module MacUnit (
	io_in_a,
	io_in_b,
	io_in_c,
	io_out_d
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_c;
	output logic [31:0] io_out_d;
	assign io_out_d =( (io_in_a * io_in_b) + io_in_c) ^ ((fiEnable && (2 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
endmodule
module PE_256 (
	clock,
	io_in_a,
	io_in_b,
	io_in_d,
	io_in_control_dataflow,
	io_in_control_propagate,
	io_in_control_shift,
	io_in_id,
	io_in_last,
	io_in_valid,
	io_out_a,
	io_out_b,
	io_out_c,
	io_out_control_dataflow,
	io_out_control_propagate,
	io_out_control_shift,
	io_out_id,
	io_out_last,
	io_out_valid
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_d;
	input io_in_control_dataflow;
	input io_in_control_propagate;
	input [4:0] io_in_control_shift;
	input [2:0] io_in_id;
	input io_in_last;
	input io_in_valid;
	output logic [31:0] io_out_a;
	output logic [31:0] io_out_b;
	output logic [31:0] io_out_c;
	output logic io_out_control_dataflow;
	output logic io_out_control_propagate;
	output logic [4:0] io_out_control_shift;
	output logic [2:0] io_out_id;
	output logic io_out_last;
	output logic io_out_valid;
	wire [31:0] _mac_unit_io_out_d;
	reg [31:0] c1;
	reg [31:0] c2;
	reg last_s;
	wire [4:0] shift_offset = (last_s != io_in_control_propagate ? io_in_control_shift : 5'h00);
	wire [31:0] _GEN = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_3 = $signed($signed(c1) >>> _GEN);
	wire [31:0] _GEN_0 = {27'h0000000, shift_offset};
	wire [31:0] _io_out_c_T = $signed($signed(c1) >>> _GEN_0);
	wire [31:0] _GEN_1 = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_8 = $signed($signed(c2) >>> _GEN_1);
	wire [31:0] _io_out_c_T_11 = $signed($signed(c2) >>> _GEN_0);
	always @(posedge clock)
		if (io_in_valid) begin
			if (io_in_control_propagate) begin
				c1 <=( io_in_d) ^ ((fiEnable && (3 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( _mac_unit_io_out_d) ^ ((fiEnable && (4 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			end
			else begin
				c1 <=( _mac_unit_io_out_d) ^ ((fiEnable && (5 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( io_in_d) ^ ((fiEnable && (6 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			end
			last_s <=( io_in_control_propagate) ^ ((fiEnable && (7 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
		end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	MacUnit mac_unit(
		.io_in_a(io_in_a),
		.io_in_b(io_in_b),
		.io_in_c((io_in_control_propagate ? c2 : c1)),
		.io_out_d(_mac_unit_io_out_d)
	,
    .fiEnable(fiEnable && ((2393 == Mesh.GlobalFiModInstNr[0]) || (2393 == Mesh.GlobalFiModInstNr[1]) || (2393 == Mesh.GlobalFiModInstNr[2]) || (2393 == Mesh.GlobalFiModInstNr[3]))));
	assign io_out_a =( io_in_a) ^ ((fiEnable && (8 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b =( io_in_b) ^ ((fiEnable && (9 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c =( (io_in_control_propagate ? _io_out_c_T + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_3[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c1 & ((32'h00000001 << _GEN) - 32'h00000001)) | _io_out_c_T[0])} : _io_out_c_T_11 + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_8[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c2 & ((32'h00000001 << _GEN_1) - 32'h00000001)) | _io_out_c_T_11[0])})) ^ ((fiEnable && (10 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_control_dataflow =( io_in_control_dataflow) ^ ((fiEnable && (11 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_propagate =( io_in_control_propagate) ^ ((fiEnable && (12 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_shift =( io_in_control_shift) ^ ((fiEnable && (13 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[4:0] : {5{1'b0}});
	assign io_out_id =( io_in_id) ^ ((fiEnable && (14 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last =( io_in_last) ^ ((fiEnable && (15 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_valid =( io_in_valid) ^ ((fiEnable && (16 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
endmodule
module Tile (
	clock,
	io_in_a_0,
	io_in_b_0,
	io_in_d_0,
	io_in_control_0_dataflow,
	io_in_control_0_propagate,
	io_in_control_0_shift,
	io_in_id_0,
	io_in_last_0,
	io_in_valid_0,
	io_out_a_0,
	io_out_c_0,
	io_out_b_0,
	io_out_control_0_dataflow,
	io_out_control_0_propagate,
	io_out_control_0_shift,
	io_out_id_0,
	io_out_last_0,
	io_out_valid_0
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a_0;
	input [31:0] io_in_b_0;
	input [31:0] io_in_d_0;
	input io_in_control_0_dataflow;
	input io_in_control_0_propagate;
	input [4:0] io_in_control_0_shift;
	input [2:0] io_in_id_0;
	input io_in_last_0;
	input io_in_valid_0;
	output logic [31:0] io_out_a_0;
	output logic [31:0] io_out_c_0;
	output logic [31:0] io_out_b_0;
	output logic io_out_control_0_dataflow;
	output logic io_out_control_0_propagate;
	output logic [4:0] io_out_control_0_shift;
	output logic [2:0] io_out_id_0;
	output logic io_out_last_0;
	output logic io_out_valid_0;
	PE_256 tile_0_0(
		.clock(clock),
		.io_in_a(io_in_a_0),
		.io_in_b(io_in_b_0),
		.io_in_d(io_in_d_0),
		.io_in_control_dataflow(io_in_control_0_dataflow),
		.io_in_control_propagate(io_in_control_0_propagate),
		.io_in_control_shift(io_in_control_0_shift),
		.io_in_id(io_in_id_0),
		.io_in_last(io_in_last_0),
		.io_in_valid(io_in_valid_0),
		.io_out_a(io_out_a_0),
		.io_out_b(io_out_b_0),
		.io_out_c(io_out_c_0),
		.io_out_control_dataflow(io_out_control_0_dataflow),
		.io_out_control_propagate(io_out_control_0_propagate),
		.io_out_control_shift(io_out_control_0_shift),
		.io_out_id(io_out_id_0),
		.io_out_last(io_out_last_0),
		.io_out_valid(io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2394 == Mesh.GlobalFiModInstNr[0]) || (2394 == Mesh.GlobalFiModInstNr[1]) || (2394 == Mesh.GlobalFiModInstNr[2]) || (2394 == Mesh.GlobalFiModInstNr[3]))));
endmodule
module Mesh (
	clock,
	io_in_a_0_0,
	io_in_a_1_0,
	io_in_a_2_0,
	io_in_a_3_0,
	io_in_a_4_0,
	io_in_a_5_0,
	io_in_a_6_0,
	io_in_a_7_0,
	io_in_a_8_0,
	io_in_a_9_0,
	io_in_a_10_0,
	io_in_a_11_0,
	io_in_a_12_0,
	io_in_a_13_0,
	io_in_a_14_0,
	io_in_a_15_0,
	io_in_b_0_0,
	io_in_b_1_0,
	io_in_b_2_0,
	io_in_b_3_0,
	io_in_b_4_0,
	io_in_b_5_0,
	io_in_b_6_0,
	io_in_b_7_0,
	io_in_b_8_0,
	io_in_b_9_0,
	io_in_b_10_0,
	io_in_b_11_0,
	io_in_b_12_0,
	io_in_b_13_0,
	io_in_b_14_0,
	io_in_b_15_0,
	io_in_d_0_0,
	io_in_d_1_0,
	io_in_d_2_0,
	io_in_d_3_0,
	io_in_d_4_0,
	io_in_d_5_0,
	io_in_d_6_0,
	io_in_d_7_0,
	io_in_d_8_0,
	io_in_d_9_0,
	io_in_d_10_0,
	io_in_d_11_0,
	io_in_d_12_0,
	io_in_d_13_0,
	io_in_d_14_0,
	io_in_d_15_0,
	io_in_control_0_0_dataflow,
	io_in_control_0_0_propagate,
	io_in_control_0_0_shift,
	io_in_control_1_0_dataflow,
	io_in_control_1_0_propagate,
	io_in_control_1_0_shift,
	io_in_control_2_0_dataflow,
	io_in_control_2_0_propagate,
	io_in_control_2_0_shift,
	io_in_control_3_0_dataflow,
	io_in_control_3_0_propagate,
	io_in_control_3_0_shift,
	io_in_control_4_0_dataflow,
	io_in_control_4_0_propagate,
	io_in_control_4_0_shift,
	io_in_control_5_0_dataflow,
	io_in_control_5_0_propagate,
	io_in_control_5_0_shift,
	io_in_control_6_0_dataflow,
	io_in_control_6_0_propagate,
	io_in_control_6_0_shift,
	io_in_control_7_0_dataflow,
	io_in_control_7_0_propagate,
	io_in_control_7_0_shift,
	io_in_control_8_0_dataflow,
	io_in_control_8_0_propagate,
	io_in_control_8_0_shift,
	io_in_control_9_0_dataflow,
	io_in_control_9_0_propagate,
	io_in_control_9_0_shift,
	io_in_control_10_0_dataflow,
	io_in_control_10_0_propagate,
	io_in_control_10_0_shift,
	io_in_control_11_0_dataflow,
	io_in_control_11_0_propagate,
	io_in_control_11_0_shift,
	io_in_control_12_0_dataflow,
	io_in_control_12_0_propagate,
	io_in_control_12_0_shift,
	io_in_control_13_0_dataflow,
	io_in_control_13_0_propagate,
	io_in_control_13_0_shift,
	io_in_control_14_0_dataflow,
	io_in_control_14_0_propagate,
	io_in_control_14_0_shift,
	io_in_control_15_0_dataflow,
	io_in_control_15_0_propagate,
	io_in_control_15_0_shift,
	io_in_id_0_0,
	io_in_id_1_0,
	io_in_id_2_0,
	io_in_id_3_0,
	io_in_id_4_0,
	io_in_id_5_0,
	io_in_id_6_0,
	io_in_id_7_0,
	io_in_id_8_0,
	io_in_id_9_0,
	io_in_id_10_0,
	io_in_id_11_0,
	io_in_id_12_0,
	io_in_id_13_0,
	io_in_id_14_0,
	io_in_id_15_0,
	io_in_last_0_0,
	io_in_last_1_0,
	io_in_last_2_0,
	io_in_last_3_0,
	io_in_last_4_0,
	io_in_last_5_0,
	io_in_last_6_0,
	io_in_last_7_0,
	io_in_last_8_0,
	io_in_last_9_0,
	io_in_last_10_0,
	io_in_last_11_0,
	io_in_last_12_0,
	io_in_last_13_0,
	io_in_last_14_0,
	io_in_last_15_0,
	io_in_valid_0_0,
	io_in_valid_1_0,
	io_in_valid_2_0,
	io_in_valid_3_0,
	io_in_valid_4_0,
	io_in_valid_5_0,
	io_in_valid_6_0,
	io_in_valid_7_0,
	io_in_valid_8_0,
	io_in_valid_9_0,
	io_in_valid_10_0,
	io_in_valid_11_0,
	io_in_valid_12_0,
	io_in_valid_13_0,
	io_in_valid_14_0,
	io_in_valid_15_0,
	io_out_b_0_0,
	io_out_b_1_0,
	io_out_b_2_0,
	io_out_b_3_0,
	io_out_b_4_0,
	io_out_b_5_0,
	io_out_b_6_0,
	io_out_b_7_0,
	io_out_b_8_0,
	io_out_b_9_0,
	io_out_b_10_0,
	io_out_b_11_0,
	io_out_b_12_0,
	io_out_b_13_0,
	io_out_b_14_0,
	io_out_b_15_0,
	io_out_c_0_0,
	io_out_c_1_0,
	io_out_c_2_0,
	io_out_c_3_0,
	io_out_c_4_0,
	io_out_c_5_0,
	io_out_c_6_0,
	io_out_c_7_0,
	io_out_c_8_0,
	io_out_c_9_0,
	io_out_c_10_0,
	io_out_c_11_0,
	io_out_c_12_0,
	io_out_c_13_0,
	io_out_c_14_0,
	io_out_c_15_0,
	io_out_valid_0_0,
	io_out_control_0_0_dataflow,
	io_out_id_0_0,
	io_out_last_0_0
, GlobalFiSignal, GlobalFiNumber, GlobalFiModInstNr);
input GlobalFiSignal;
wire [31:0] GlobalFiSignal;
input GlobalFiNumber;
wire [31:0] GlobalFiNumber;
input GlobalFiModInstNr;
wire [15:0] GlobalFiModInstNr[4];
wire fiEnable;
assign fiEnable = (1 == GlobalFiModInstNr[0]) || (1 == GlobalFiModInstNr[1]) || (1 == GlobalFiModInstNr[2]) || (1 == GlobalFiModInstNr[3]);

	input clock;
	input [31:0] io_in_a_0_0;
	input [31:0] io_in_a_1_0;
	input [31:0] io_in_a_2_0;
	input [31:0] io_in_a_3_0;
	input [31:0] io_in_a_4_0;
	input [31:0] io_in_a_5_0;
	input [31:0] io_in_a_6_0;
	input [31:0] io_in_a_7_0;
	input [31:0] io_in_a_8_0;
	input [31:0] io_in_a_9_0;
	input [31:0] io_in_a_10_0;
	input [31:0] io_in_a_11_0;
	input [31:0] io_in_a_12_0;
	input [31:0] io_in_a_13_0;
	input [31:0] io_in_a_14_0;
	input [31:0] io_in_a_15_0;
	input [31:0] io_in_b_0_0;
	input [31:0] io_in_b_1_0;
	input [31:0] io_in_b_2_0;
	input [31:0] io_in_b_3_0;
	input [31:0] io_in_b_4_0;
	input [31:0] io_in_b_5_0;
	input [31:0] io_in_b_6_0;
	input [31:0] io_in_b_7_0;
	input [31:0] io_in_b_8_0;
	input [31:0] io_in_b_9_0;
	input [31:0] io_in_b_10_0;
	input [31:0] io_in_b_11_0;
	input [31:0] io_in_b_12_0;
	input [31:0] io_in_b_13_0;
	input [31:0] io_in_b_14_0;
	input [31:0] io_in_b_15_0;
	input [31:0] io_in_d_0_0;
	input [31:0] io_in_d_1_0;
	input [31:0] io_in_d_2_0;
	input [31:0] io_in_d_3_0;
	input [31:0] io_in_d_4_0;
	input [31:0] io_in_d_5_0;
	input [31:0] io_in_d_6_0;
	input [31:0] io_in_d_7_0;
	input [31:0] io_in_d_8_0;
	input [31:0] io_in_d_9_0;
	input [31:0] io_in_d_10_0;
	input [31:0] io_in_d_11_0;
	input [31:0] io_in_d_12_0;
	input [31:0] io_in_d_13_0;
	input [31:0] io_in_d_14_0;
	input [31:0] io_in_d_15_0;
	input io_in_control_0_0_dataflow;
	input io_in_control_0_0_propagate;
	input [4:0] io_in_control_0_0_shift;
	input io_in_control_1_0_dataflow;
	input io_in_control_1_0_propagate;
	input [4:0] io_in_control_1_0_shift;
	input io_in_control_2_0_dataflow;
	input io_in_control_2_0_propagate;
	input [4:0] io_in_control_2_0_shift;
	input io_in_control_3_0_dataflow;
	input io_in_control_3_0_propagate;
	input [4:0] io_in_control_3_0_shift;
	input io_in_control_4_0_dataflow;
	input io_in_control_4_0_propagate;
	input [4:0] io_in_control_4_0_shift;
	input io_in_control_5_0_dataflow;
	input io_in_control_5_0_propagate;
	input [4:0] io_in_control_5_0_shift;
	input io_in_control_6_0_dataflow;
	input io_in_control_6_0_propagate;
	input [4:0] io_in_control_6_0_shift;
	input io_in_control_7_0_dataflow;
	input io_in_control_7_0_propagate;
	input [4:0] io_in_control_7_0_shift;
	input io_in_control_8_0_dataflow;
	input io_in_control_8_0_propagate;
	input [4:0] io_in_control_8_0_shift;
	input io_in_control_9_0_dataflow;
	input io_in_control_9_0_propagate;
	input [4:0] io_in_control_9_0_shift;
	input io_in_control_10_0_dataflow;
	input io_in_control_10_0_propagate;
	input [4:0] io_in_control_10_0_shift;
	input io_in_control_11_0_dataflow;
	input io_in_control_11_0_propagate;
	input [4:0] io_in_control_11_0_shift;
	input io_in_control_12_0_dataflow;
	input io_in_control_12_0_propagate;
	input [4:0] io_in_control_12_0_shift;
	input io_in_control_13_0_dataflow;
	input io_in_control_13_0_propagate;
	input [4:0] io_in_control_13_0_shift;
	input io_in_control_14_0_dataflow;
	input io_in_control_14_0_propagate;
	input [4:0] io_in_control_14_0_shift;
	input io_in_control_15_0_dataflow;
	input io_in_control_15_0_propagate;
	input [4:0] io_in_control_15_0_shift;
	input [2:0] io_in_id_0_0;
	input [2:0] io_in_id_1_0;
	input [2:0] io_in_id_2_0;
	input [2:0] io_in_id_3_0;
	input [2:0] io_in_id_4_0;
	input [2:0] io_in_id_5_0;
	input [2:0] io_in_id_6_0;
	input [2:0] io_in_id_7_0;
	input [2:0] io_in_id_8_0;
	input [2:0] io_in_id_9_0;
	input [2:0] io_in_id_10_0;
	input [2:0] io_in_id_11_0;
	input [2:0] io_in_id_12_0;
	input [2:0] io_in_id_13_0;
	input [2:0] io_in_id_14_0;
	input [2:0] io_in_id_15_0;
	input io_in_last_0_0;
	input io_in_last_1_0;
	input io_in_last_2_0;
	input io_in_last_3_0;
	input io_in_last_4_0;
	input io_in_last_5_0;
	input io_in_last_6_0;
	input io_in_last_7_0;
	input io_in_last_8_0;
	input io_in_last_9_0;
	input io_in_last_10_0;
	input io_in_last_11_0;
	input io_in_last_12_0;
	input io_in_last_13_0;
	input io_in_last_14_0;
	input io_in_last_15_0;
	input io_in_valid_0_0;
	input io_in_valid_1_0;
	input io_in_valid_2_0;
	input io_in_valid_3_0;
	input io_in_valid_4_0;
	input io_in_valid_5_0;
	input io_in_valid_6_0;
	input io_in_valid_7_0;
	input io_in_valid_8_0;
	input io_in_valid_9_0;
	input io_in_valid_10_0;
	input io_in_valid_11_0;
	input io_in_valid_12_0;
	input io_in_valid_13_0;
	input io_in_valid_14_0;
	input io_in_valid_15_0;
	output logic [31:0] io_out_b_0_0;
	output logic [31:0] io_out_b_1_0;
	output logic [31:0] io_out_b_2_0;
	output logic [31:0] io_out_b_3_0;
	output logic [31:0] io_out_b_4_0;
	output logic [31:0] io_out_b_5_0;
	output logic [31:0] io_out_b_6_0;
	output logic [31:0] io_out_b_7_0;
	output logic [31:0] io_out_b_8_0;
	output logic [31:0] io_out_b_9_0;
	output logic [31:0] io_out_b_10_0;
	output logic [31:0] io_out_b_11_0;
	output logic [31:0] io_out_b_12_0;
	output logic [31:0] io_out_b_13_0;
	output logic [31:0] io_out_b_14_0;
	output logic [31:0] io_out_b_15_0;
	output logic [31:0] io_out_c_0_0;
	output logic [31:0] io_out_c_1_0;
	output logic [31:0] io_out_c_2_0;
	output logic [31:0] io_out_c_3_0;
	output logic [31:0] io_out_c_4_0;
	output logic [31:0] io_out_c_5_0;
	output logic [31:0] io_out_c_6_0;
	output logic [31:0] io_out_c_7_0;
	output logic [31:0] io_out_c_8_0;
	output logic [31:0] io_out_c_9_0;
	output logic [31:0] io_out_c_10_0;
	output logic [31:0] io_out_c_11_0;
	output logic [31:0] io_out_c_12_0;
	output logic [31:0] io_out_c_13_0;
	output logic [31:0] io_out_c_14_0;
	output logic [31:0] io_out_c_15_0;
	output logic io_out_valid_0_0;
	output logic io_out_control_0_0_dataflow;
	output logic [2:0] io_out_id_0_0;
	output logic io_out_last_0_0;
	wire [31:0] _mesh_15_15_io_out_a_0;
	wire [31:0] _mesh_15_15_io_out_c_0;
	wire [31:0] _mesh_15_15_io_out_b_0;
	wire _mesh_15_15_io_out_control_0_dataflow;
	wire _mesh_15_15_io_out_control_0_propagate;
	wire [4:0] _mesh_15_15_io_out_control_0_shift;
	wire [2:0] _mesh_15_15_io_out_id_0;
	wire _mesh_15_15_io_out_last_0;
	wire _mesh_15_15_io_out_valid_0;
	wire [31:0] _mesh_15_14_io_out_a_0;
	wire [31:0] _mesh_15_14_io_out_c_0;
	wire [31:0] _mesh_15_14_io_out_b_0;
	wire _mesh_15_14_io_out_control_0_dataflow;
	wire _mesh_15_14_io_out_control_0_propagate;
	wire [4:0] _mesh_15_14_io_out_control_0_shift;
	wire [2:0] _mesh_15_14_io_out_id_0;
	wire _mesh_15_14_io_out_last_0;
	wire _mesh_15_14_io_out_valid_0;
	wire [31:0] _mesh_15_13_io_out_a_0;
	wire [31:0] _mesh_15_13_io_out_c_0;
	wire [31:0] _mesh_15_13_io_out_b_0;
	wire _mesh_15_13_io_out_control_0_dataflow;
	wire _mesh_15_13_io_out_control_0_propagate;
	wire [4:0] _mesh_15_13_io_out_control_0_shift;
	wire [2:0] _mesh_15_13_io_out_id_0;
	wire _mesh_15_13_io_out_last_0;
	wire _mesh_15_13_io_out_valid_0;
	wire [31:0] _mesh_15_12_io_out_a_0;
	wire [31:0] _mesh_15_12_io_out_c_0;
	wire [31:0] _mesh_15_12_io_out_b_0;
	wire _mesh_15_12_io_out_control_0_dataflow;
	wire _mesh_15_12_io_out_control_0_propagate;
	wire [4:0] _mesh_15_12_io_out_control_0_shift;
	wire [2:0] _mesh_15_12_io_out_id_0;
	wire _mesh_15_12_io_out_last_0;
	wire _mesh_15_12_io_out_valid_0;
	wire [31:0] _mesh_15_11_io_out_a_0;
	wire [31:0] _mesh_15_11_io_out_c_0;
	wire [31:0] _mesh_15_11_io_out_b_0;
	wire _mesh_15_11_io_out_control_0_dataflow;
	wire _mesh_15_11_io_out_control_0_propagate;
	wire [4:0] _mesh_15_11_io_out_control_0_shift;
	wire [2:0] _mesh_15_11_io_out_id_0;
	wire _mesh_15_11_io_out_last_0;
	wire _mesh_15_11_io_out_valid_0;
	wire [31:0] _mesh_15_10_io_out_a_0;
	wire [31:0] _mesh_15_10_io_out_c_0;
	wire [31:0] _mesh_15_10_io_out_b_0;
	wire _mesh_15_10_io_out_control_0_dataflow;
	wire _mesh_15_10_io_out_control_0_propagate;
	wire [4:0] _mesh_15_10_io_out_control_0_shift;
	wire [2:0] _mesh_15_10_io_out_id_0;
	wire _mesh_15_10_io_out_last_0;
	wire _mesh_15_10_io_out_valid_0;
	wire [31:0] _mesh_15_9_io_out_a_0;
	wire [31:0] _mesh_15_9_io_out_c_0;
	wire [31:0] _mesh_15_9_io_out_b_0;
	wire _mesh_15_9_io_out_control_0_dataflow;
	wire _mesh_15_9_io_out_control_0_propagate;
	wire [4:0] _mesh_15_9_io_out_control_0_shift;
	wire [2:0] _mesh_15_9_io_out_id_0;
	wire _mesh_15_9_io_out_last_0;
	wire _mesh_15_9_io_out_valid_0;
	wire [31:0] _mesh_15_8_io_out_a_0;
	wire [31:0] _mesh_15_8_io_out_c_0;
	wire [31:0] _mesh_15_8_io_out_b_0;
	wire _mesh_15_8_io_out_control_0_dataflow;
	wire _mesh_15_8_io_out_control_0_propagate;
	wire [4:0] _mesh_15_8_io_out_control_0_shift;
	wire [2:0] _mesh_15_8_io_out_id_0;
	wire _mesh_15_8_io_out_last_0;
	wire _mesh_15_8_io_out_valid_0;
	wire [31:0] _mesh_15_7_io_out_a_0;
	wire [31:0] _mesh_15_7_io_out_c_0;
	wire [31:0] _mesh_15_7_io_out_b_0;
	wire _mesh_15_7_io_out_control_0_dataflow;
	wire _mesh_15_7_io_out_control_0_propagate;
	wire [4:0] _mesh_15_7_io_out_control_0_shift;
	wire [2:0] _mesh_15_7_io_out_id_0;
	wire _mesh_15_7_io_out_last_0;
	wire _mesh_15_7_io_out_valid_0;
	wire [31:0] _mesh_15_6_io_out_a_0;
	wire [31:0] _mesh_15_6_io_out_c_0;
	wire [31:0] _mesh_15_6_io_out_b_0;
	wire _mesh_15_6_io_out_control_0_dataflow;
	wire _mesh_15_6_io_out_control_0_propagate;
	wire [4:0] _mesh_15_6_io_out_control_0_shift;
	wire [2:0] _mesh_15_6_io_out_id_0;
	wire _mesh_15_6_io_out_last_0;
	wire _mesh_15_6_io_out_valid_0;
	wire [31:0] _mesh_15_5_io_out_a_0;
	wire [31:0] _mesh_15_5_io_out_c_0;
	wire [31:0] _mesh_15_5_io_out_b_0;
	wire _mesh_15_5_io_out_control_0_dataflow;
	wire _mesh_15_5_io_out_control_0_propagate;
	wire [4:0] _mesh_15_5_io_out_control_0_shift;
	wire [2:0] _mesh_15_5_io_out_id_0;
	wire _mesh_15_5_io_out_last_0;
	wire _mesh_15_5_io_out_valid_0;
	wire [31:0] _mesh_15_4_io_out_a_0;
	wire [31:0] _mesh_15_4_io_out_c_0;
	wire [31:0] _mesh_15_4_io_out_b_0;
	wire _mesh_15_4_io_out_control_0_dataflow;
	wire _mesh_15_4_io_out_control_0_propagate;
	wire [4:0] _mesh_15_4_io_out_control_0_shift;
	wire [2:0] _mesh_15_4_io_out_id_0;
	wire _mesh_15_4_io_out_last_0;
	wire _mesh_15_4_io_out_valid_0;
	wire [31:0] _mesh_15_3_io_out_a_0;
	wire [31:0] _mesh_15_3_io_out_c_0;
	wire [31:0] _mesh_15_3_io_out_b_0;
	wire _mesh_15_3_io_out_control_0_dataflow;
	wire _mesh_15_3_io_out_control_0_propagate;
	wire [4:0] _mesh_15_3_io_out_control_0_shift;
	wire [2:0] _mesh_15_3_io_out_id_0;
	wire _mesh_15_3_io_out_last_0;
	wire _mesh_15_3_io_out_valid_0;
	wire [31:0] _mesh_15_2_io_out_a_0;
	wire [31:0] _mesh_15_2_io_out_c_0;
	wire [31:0] _mesh_15_2_io_out_b_0;
	wire _mesh_15_2_io_out_control_0_dataflow;
	wire _mesh_15_2_io_out_control_0_propagate;
	wire [4:0] _mesh_15_2_io_out_control_0_shift;
	wire [2:0] _mesh_15_2_io_out_id_0;
	wire _mesh_15_2_io_out_last_0;
	wire _mesh_15_2_io_out_valid_0;
	wire [31:0] _mesh_15_1_io_out_a_0;
	wire [31:0] _mesh_15_1_io_out_c_0;
	wire [31:0] _mesh_15_1_io_out_b_0;
	wire _mesh_15_1_io_out_control_0_dataflow;
	wire _mesh_15_1_io_out_control_0_propagate;
	wire [4:0] _mesh_15_1_io_out_control_0_shift;
	wire [2:0] _mesh_15_1_io_out_id_0;
	wire _mesh_15_1_io_out_last_0;
	wire _mesh_15_1_io_out_valid_0;
	wire [31:0] _mesh_15_0_io_out_a_0;
	wire [31:0] _mesh_15_0_io_out_c_0;
	wire [31:0] _mesh_15_0_io_out_b_0;
	wire _mesh_15_0_io_out_control_0_dataflow;
	wire _mesh_15_0_io_out_control_0_propagate;
	wire [4:0] _mesh_15_0_io_out_control_0_shift;
	wire [2:0] _mesh_15_0_io_out_id_0;
	wire _mesh_15_0_io_out_last_0;
	wire _mesh_15_0_io_out_valid_0;
	wire [31:0] _mesh_14_15_io_out_a_0;
	wire [31:0] _mesh_14_15_io_out_c_0;
	wire [31:0] _mesh_14_15_io_out_b_0;
	wire _mesh_14_15_io_out_control_0_dataflow;
	wire _mesh_14_15_io_out_control_0_propagate;
	wire [4:0] _mesh_14_15_io_out_control_0_shift;
	wire [2:0] _mesh_14_15_io_out_id_0;
	wire _mesh_14_15_io_out_last_0;
	wire _mesh_14_15_io_out_valid_0;
	wire [31:0] _mesh_14_14_io_out_a_0;
	wire [31:0] _mesh_14_14_io_out_c_0;
	wire [31:0] _mesh_14_14_io_out_b_0;
	wire _mesh_14_14_io_out_control_0_dataflow;
	wire _mesh_14_14_io_out_control_0_propagate;
	wire [4:0] _mesh_14_14_io_out_control_0_shift;
	wire [2:0] _mesh_14_14_io_out_id_0;
	wire _mesh_14_14_io_out_last_0;
	wire _mesh_14_14_io_out_valid_0;
	wire [31:0] _mesh_14_13_io_out_a_0;
	wire [31:0] _mesh_14_13_io_out_c_0;
	wire [31:0] _mesh_14_13_io_out_b_0;
	wire _mesh_14_13_io_out_control_0_dataflow;
	wire _mesh_14_13_io_out_control_0_propagate;
	wire [4:0] _mesh_14_13_io_out_control_0_shift;
	wire [2:0] _mesh_14_13_io_out_id_0;
	wire _mesh_14_13_io_out_last_0;
	wire _mesh_14_13_io_out_valid_0;
	wire [31:0] _mesh_14_12_io_out_a_0;
	wire [31:0] _mesh_14_12_io_out_c_0;
	wire [31:0] _mesh_14_12_io_out_b_0;
	wire _mesh_14_12_io_out_control_0_dataflow;
	wire _mesh_14_12_io_out_control_0_propagate;
	wire [4:0] _mesh_14_12_io_out_control_0_shift;
	wire [2:0] _mesh_14_12_io_out_id_0;
	wire _mesh_14_12_io_out_last_0;
	wire _mesh_14_12_io_out_valid_0;
	wire [31:0] _mesh_14_11_io_out_a_0;
	wire [31:0] _mesh_14_11_io_out_c_0;
	wire [31:0] _mesh_14_11_io_out_b_0;
	wire _mesh_14_11_io_out_control_0_dataflow;
	wire _mesh_14_11_io_out_control_0_propagate;
	wire [4:0] _mesh_14_11_io_out_control_0_shift;
	wire [2:0] _mesh_14_11_io_out_id_0;
	wire _mesh_14_11_io_out_last_0;
	wire _mesh_14_11_io_out_valid_0;
	wire [31:0] _mesh_14_10_io_out_a_0;
	wire [31:0] _mesh_14_10_io_out_c_0;
	wire [31:0] _mesh_14_10_io_out_b_0;
	wire _mesh_14_10_io_out_control_0_dataflow;
	wire _mesh_14_10_io_out_control_0_propagate;
	wire [4:0] _mesh_14_10_io_out_control_0_shift;
	wire [2:0] _mesh_14_10_io_out_id_0;
	wire _mesh_14_10_io_out_last_0;
	wire _mesh_14_10_io_out_valid_0;
	wire [31:0] _mesh_14_9_io_out_a_0;
	wire [31:0] _mesh_14_9_io_out_c_0;
	wire [31:0] _mesh_14_9_io_out_b_0;
	wire _mesh_14_9_io_out_control_0_dataflow;
	wire _mesh_14_9_io_out_control_0_propagate;
	wire [4:0] _mesh_14_9_io_out_control_0_shift;
	wire [2:0] _mesh_14_9_io_out_id_0;
	wire _mesh_14_9_io_out_last_0;
	wire _mesh_14_9_io_out_valid_0;
	wire [31:0] _mesh_14_8_io_out_a_0;
	wire [31:0] _mesh_14_8_io_out_c_0;
	wire [31:0] _mesh_14_8_io_out_b_0;
	wire _mesh_14_8_io_out_control_0_dataflow;
	wire _mesh_14_8_io_out_control_0_propagate;
	wire [4:0] _mesh_14_8_io_out_control_0_shift;
	wire [2:0] _mesh_14_8_io_out_id_0;
	wire _mesh_14_8_io_out_last_0;
	wire _mesh_14_8_io_out_valid_0;
	wire [31:0] _mesh_14_7_io_out_a_0;
	wire [31:0] _mesh_14_7_io_out_c_0;
	wire [31:0] _mesh_14_7_io_out_b_0;
	wire _mesh_14_7_io_out_control_0_dataflow;
	wire _mesh_14_7_io_out_control_0_propagate;
	wire [4:0] _mesh_14_7_io_out_control_0_shift;
	wire [2:0] _mesh_14_7_io_out_id_0;
	wire _mesh_14_7_io_out_last_0;
	wire _mesh_14_7_io_out_valid_0;
	wire [31:0] _mesh_14_6_io_out_a_0;
	wire [31:0] _mesh_14_6_io_out_c_0;
	wire [31:0] _mesh_14_6_io_out_b_0;
	wire _mesh_14_6_io_out_control_0_dataflow;
	wire _mesh_14_6_io_out_control_0_propagate;
	wire [4:0] _mesh_14_6_io_out_control_0_shift;
	wire [2:0] _mesh_14_6_io_out_id_0;
	wire _mesh_14_6_io_out_last_0;
	wire _mesh_14_6_io_out_valid_0;
	wire [31:0] _mesh_14_5_io_out_a_0;
	wire [31:0] _mesh_14_5_io_out_c_0;
	wire [31:0] _mesh_14_5_io_out_b_0;
	wire _mesh_14_5_io_out_control_0_dataflow;
	wire _mesh_14_5_io_out_control_0_propagate;
	wire [4:0] _mesh_14_5_io_out_control_0_shift;
	wire [2:0] _mesh_14_5_io_out_id_0;
	wire _mesh_14_5_io_out_last_0;
	wire _mesh_14_5_io_out_valid_0;
	wire [31:0] _mesh_14_4_io_out_a_0;
	wire [31:0] _mesh_14_4_io_out_c_0;
	wire [31:0] _mesh_14_4_io_out_b_0;
	wire _mesh_14_4_io_out_control_0_dataflow;
	wire _mesh_14_4_io_out_control_0_propagate;
	wire [4:0] _mesh_14_4_io_out_control_0_shift;
	wire [2:0] _mesh_14_4_io_out_id_0;
	wire _mesh_14_4_io_out_last_0;
	wire _mesh_14_4_io_out_valid_0;
	wire [31:0] _mesh_14_3_io_out_a_0;
	wire [31:0] _mesh_14_3_io_out_c_0;
	wire [31:0] _mesh_14_3_io_out_b_0;
	wire _mesh_14_3_io_out_control_0_dataflow;
	wire _mesh_14_3_io_out_control_0_propagate;
	wire [4:0] _mesh_14_3_io_out_control_0_shift;
	wire [2:0] _mesh_14_3_io_out_id_0;
	wire _mesh_14_3_io_out_last_0;
	wire _mesh_14_3_io_out_valid_0;
	wire [31:0] _mesh_14_2_io_out_a_0;
	wire [31:0] _mesh_14_2_io_out_c_0;
	wire [31:0] _mesh_14_2_io_out_b_0;
	wire _mesh_14_2_io_out_control_0_dataflow;
	wire _mesh_14_2_io_out_control_0_propagate;
	wire [4:0] _mesh_14_2_io_out_control_0_shift;
	wire [2:0] _mesh_14_2_io_out_id_0;
	wire _mesh_14_2_io_out_last_0;
	wire _mesh_14_2_io_out_valid_0;
	wire [31:0] _mesh_14_1_io_out_a_0;
	wire [31:0] _mesh_14_1_io_out_c_0;
	wire [31:0] _mesh_14_1_io_out_b_0;
	wire _mesh_14_1_io_out_control_0_dataflow;
	wire _mesh_14_1_io_out_control_0_propagate;
	wire [4:0] _mesh_14_1_io_out_control_0_shift;
	wire [2:0] _mesh_14_1_io_out_id_0;
	wire _mesh_14_1_io_out_last_0;
	wire _mesh_14_1_io_out_valid_0;
	wire [31:0] _mesh_14_0_io_out_a_0;
	wire [31:0] _mesh_14_0_io_out_c_0;
	wire [31:0] _mesh_14_0_io_out_b_0;
	wire _mesh_14_0_io_out_control_0_dataflow;
	wire _mesh_14_0_io_out_control_0_propagate;
	wire [4:0] _mesh_14_0_io_out_control_0_shift;
	wire [2:0] _mesh_14_0_io_out_id_0;
	wire _mesh_14_0_io_out_last_0;
	wire _mesh_14_0_io_out_valid_0;
	wire [31:0] _mesh_13_15_io_out_a_0;
	wire [31:0] _mesh_13_15_io_out_c_0;
	wire [31:0] _mesh_13_15_io_out_b_0;
	wire _mesh_13_15_io_out_control_0_dataflow;
	wire _mesh_13_15_io_out_control_0_propagate;
	wire [4:0] _mesh_13_15_io_out_control_0_shift;
	wire [2:0] _mesh_13_15_io_out_id_0;
	wire _mesh_13_15_io_out_last_0;
	wire _mesh_13_15_io_out_valid_0;
	wire [31:0] _mesh_13_14_io_out_a_0;
	wire [31:0] _mesh_13_14_io_out_c_0;
	wire [31:0] _mesh_13_14_io_out_b_0;
	wire _mesh_13_14_io_out_control_0_dataflow;
	wire _mesh_13_14_io_out_control_0_propagate;
	wire [4:0] _mesh_13_14_io_out_control_0_shift;
	wire [2:0] _mesh_13_14_io_out_id_0;
	wire _mesh_13_14_io_out_last_0;
	wire _mesh_13_14_io_out_valid_0;
	wire [31:0] _mesh_13_13_io_out_a_0;
	wire [31:0] _mesh_13_13_io_out_c_0;
	wire [31:0] _mesh_13_13_io_out_b_0;
	wire _mesh_13_13_io_out_control_0_dataflow;
	wire _mesh_13_13_io_out_control_0_propagate;
	wire [4:0] _mesh_13_13_io_out_control_0_shift;
	wire [2:0] _mesh_13_13_io_out_id_0;
	wire _mesh_13_13_io_out_last_0;
	wire _mesh_13_13_io_out_valid_0;
	wire [31:0] _mesh_13_12_io_out_a_0;
	wire [31:0] _mesh_13_12_io_out_c_0;
	wire [31:0] _mesh_13_12_io_out_b_0;
	wire _mesh_13_12_io_out_control_0_dataflow;
	wire _mesh_13_12_io_out_control_0_propagate;
	wire [4:0] _mesh_13_12_io_out_control_0_shift;
	wire [2:0] _mesh_13_12_io_out_id_0;
	wire _mesh_13_12_io_out_last_0;
	wire _mesh_13_12_io_out_valid_0;
	wire [31:0] _mesh_13_11_io_out_a_0;
	wire [31:0] _mesh_13_11_io_out_c_0;
	wire [31:0] _mesh_13_11_io_out_b_0;
	wire _mesh_13_11_io_out_control_0_dataflow;
	wire _mesh_13_11_io_out_control_0_propagate;
	wire [4:0] _mesh_13_11_io_out_control_0_shift;
	wire [2:0] _mesh_13_11_io_out_id_0;
	wire _mesh_13_11_io_out_last_0;
	wire _mesh_13_11_io_out_valid_0;
	wire [31:0] _mesh_13_10_io_out_a_0;
	wire [31:0] _mesh_13_10_io_out_c_0;
	wire [31:0] _mesh_13_10_io_out_b_0;
	wire _mesh_13_10_io_out_control_0_dataflow;
	wire _mesh_13_10_io_out_control_0_propagate;
	wire [4:0] _mesh_13_10_io_out_control_0_shift;
	wire [2:0] _mesh_13_10_io_out_id_0;
	wire _mesh_13_10_io_out_last_0;
	wire _mesh_13_10_io_out_valid_0;
	wire [31:0] _mesh_13_9_io_out_a_0;
	wire [31:0] _mesh_13_9_io_out_c_0;
	wire [31:0] _mesh_13_9_io_out_b_0;
	wire _mesh_13_9_io_out_control_0_dataflow;
	wire _mesh_13_9_io_out_control_0_propagate;
	wire [4:0] _mesh_13_9_io_out_control_0_shift;
	wire [2:0] _mesh_13_9_io_out_id_0;
	wire _mesh_13_9_io_out_last_0;
	wire _mesh_13_9_io_out_valid_0;
	wire [31:0] _mesh_13_8_io_out_a_0;
	wire [31:0] _mesh_13_8_io_out_c_0;
	wire [31:0] _mesh_13_8_io_out_b_0;
	wire _mesh_13_8_io_out_control_0_dataflow;
	wire _mesh_13_8_io_out_control_0_propagate;
	wire [4:0] _mesh_13_8_io_out_control_0_shift;
	wire [2:0] _mesh_13_8_io_out_id_0;
	wire _mesh_13_8_io_out_last_0;
	wire _mesh_13_8_io_out_valid_0;
	wire [31:0] _mesh_13_7_io_out_a_0;
	wire [31:0] _mesh_13_7_io_out_c_0;
	wire [31:0] _mesh_13_7_io_out_b_0;
	wire _mesh_13_7_io_out_control_0_dataflow;
	wire _mesh_13_7_io_out_control_0_propagate;
	wire [4:0] _mesh_13_7_io_out_control_0_shift;
	wire [2:0] _mesh_13_7_io_out_id_0;
	wire _mesh_13_7_io_out_last_0;
	wire _mesh_13_7_io_out_valid_0;
	wire [31:0] _mesh_13_6_io_out_a_0;
	wire [31:0] _mesh_13_6_io_out_c_0;
	wire [31:0] _mesh_13_6_io_out_b_0;
	wire _mesh_13_6_io_out_control_0_dataflow;
	wire _mesh_13_6_io_out_control_0_propagate;
	wire [4:0] _mesh_13_6_io_out_control_0_shift;
	wire [2:0] _mesh_13_6_io_out_id_0;
	wire _mesh_13_6_io_out_last_0;
	wire _mesh_13_6_io_out_valid_0;
	wire [31:0] _mesh_13_5_io_out_a_0;
	wire [31:0] _mesh_13_5_io_out_c_0;
	wire [31:0] _mesh_13_5_io_out_b_0;
	wire _mesh_13_5_io_out_control_0_dataflow;
	wire _mesh_13_5_io_out_control_0_propagate;
	wire [4:0] _mesh_13_5_io_out_control_0_shift;
	wire [2:0] _mesh_13_5_io_out_id_0;
	wire _mesh_13_5_io_out_last_0;
	wire _mesh_13_5_io_out_valid_0;
	wire [31:0] _mesh_13_4_io_out_a_0;
	wire [31:0] _mesh_13_4_io_out_c_0;
	wire [31:0] _mesh_13_4_io_out_b_0;
	wire _mesh_13_4_io_out_control_0_dataflow;
	wire _mesh_13_4_io_out_control_0_propagate;
	wire [4:0] _mesh_13_4_io_out_control_0_shift;
	wire [2:0] _mesh_13_4_io_out_id_0;
	wire _mesh_13_4_io_out_last_0;
	wire _mesh_13_4_io_out_valid_0;
	wire [31:0] _mesh_13_3_io_out_a_0;
	wire [31:0] _mesh_13_3_io_out_c_0;
	wire [31:0] _mesh_13_3_io_out_b_0;
	wire _mesh_13_3_io_out_control_0_dataflow;
	wire _mesh_13_3_io_out_control_0_propagate;
	wire [4:0] _mesh_13_3_io_out_control_0_shift;
	wire [2:0] _mesh_13_3_io_out_id_0;
	wire _mesh_13_3_io_out_last_0;
	wire _mesh_13_3_io_out_valid_0;
	wire [31:0] _mesh_13_2_io_out_a_0;
	wire [31:0] _mesh_13_2_io_out_c_0;
	wire [31:0] _mesh_13_2_io_out_b_0;
	wire _mesh_13_2_io_out_control_0_dataflow;
	wire _mesh_13_2_io_out_control_0_propagate;
	wire [4:0] _mesh_13_2_io_out_control_0_shift;
	wire [2:0] _mesh_13_2_io_out_id_0;
	wire _mesh_13_2_io_out_last_0;
	wire _mesh_13_2_io_out_valid_0;
	wire [31:0] _mesh_13_1_io_out_a_0;
	wire [31:0] _mesh_13_1_io_out_c_0;
	wire [31:0] _mesh_13_1_io_out_b_0;
	wire _mesh_13_1_io_out_control_0_dataflow;
	wire _mesh_13_1_io_out_control_0_propagate;
	wire [4:0] _mesh_13_1_io_out_control_0_shift;
	wire [2:0] _mesh_13_1_io_out_id_0;
	wire _mesh_13_1_io_out_last_0;
	wire _mesh_13_1_io_out_valid_0;
	wire [31:0] _mesh_13_0_io_out_a_0;
	wire [31:0] _mesh_13_0_io_out_c_0;
	wire [31:0] _mesh_13_0_io_out_b_0;
	wire _mesh_13_0_io_out_control_0_dataflow;
	wire _mesh_13_0_io_out_control_0_propagate;
	wire [4:0] _mesh_13_0_io_out_control_0_shift;
	wire [2:0] _mesh_13_0_io_out_id_0;
	wire _mesh_13_0_io_out_last_0;
	wire _mesh_13_0_io_out_valid_0;
	wire [31:0] _mesh_12_15_io_out_a_0;
	wire [31:0] _mesh_12_15_io_out_c_0;
	wire [31:0] _mesh_12_15_io_out_b_0;
	wire _mesh_12_15_io_out_control_0_dataflow;
	wire _mesh_12_15_io_out_control_0_propagate;
	wire [4:0] _mesh_12_15_io_out_control_0_shift;
	wire [2:0] _mesh_12_15_io_out_id_0;
	wire _mesh_12_15_io_out_last_0;
	wire _mesh_12_15_io_out_valid_0;
	wire [31:0] _mesh_12_14_io_out_a_0;
	wire [31:0] _mesh_12_14_io_out_c_0;
	wire [31:0] _mesh_12_14_io_out_b_0;
	wire _mesh_12_14_io_out_control_0_dataflow;
	wire _mesh_12_14_io_out_control_0_propagate;
	wire [4:0] _mesh_12_14_io_out_control_0_shift;
	wire [2:0] _mesh_12_14_io_out_id_0;
	wire _mesh_12_14_io_out_last_0;
	wire _mesh_12_14_io_out_valid_0;
	wire [31:0] _mesh_12_13_io_out_a_0;
	wire [31:0] _mesh_12_13_io_out_c_0;
	wire [31:0] _mesh_12_13_io_out_b_0;
	wire _mesh_12_13_io_out_control_0_dataflow;
	wire _mesh_12_13_io_out_control_0_propagate;
	wire [4:0] _mesh_12_13_io_out_control_0_shift;
	wire [2:0] _mesh_12_13_io_out_id_0;
	wire _mesh_12_13_io_out_last_0;
	wire _mesh_12_13_io_out_valid_0;
	wire [31:0] _mesh_12_12_io_out_a_0;
	wire [31:0] _mesh_12_12_io_out_c_0;
	wire [31:0] _mesh_12_12_io_out_b_0;
	wire _mesh_12_12_io_out_control_0_dataflow;
	wire _mesh_12_12_io_out_control_0_propagate;
	wire [4:0] _mesh_12_12_io_out_control_0_shift;
	wire [2:0] _mesh_12_12_io_out_id_0;
	wire _mesh_12_12_io_out_last_0;
	wire _mesh_12_12_io_out_valid_0;
	wire [31:0] _mesh_12_11_io_out_a_0;
	wire [31:0] _mesh_12_11_io_out_c_0;
	wire [31:0] _mesh_12_11_io_out_b_0;
	wire _mesh_12_11_io_out_control_0_dataflow;
	wire _mesh_12_11_io_out_control_0_propagate;
	wire [4:0] _mesh_12_11_io_out_control_0_shift;
	wire [2:0] _mesh_12_11_io_out_id_0;
	wire _mesh_12_11_io_out_last_0;
	wire _mesh_12_11_io_out_valid_0;
	wire [31:0] _mesh_12_10_io_out_a_0;
	wire [31:0] _mesh_12_10_io_out_c_0;
	wire [31:0] _mesh_12_10_io_out_b_0;
	wire _mesh_12_10_io_out_control_0_dataflow;
	wire _mesh_12_10_io_out_control_0_propagate;
	wire [4:0] _mesh_12_10_io_out_control_0_shift;
	wire [2:0] _mesh_12_10_io_out_id_0;
	wire _mesh_12_10_io_out_last_0;
	wire _mesh_12_10_io_out_valid_0;
	wire [31:0] _mesh_12_9_io_out_a_0;
	wire [31:0] _mesh_12_9_io_out_c_0;
	wire [31:0] _mesh_12_9_io_out_b_0;
	wire _mesh_12_9_io_out_control_0_dataflow;
	wire _mesh_12_9_io_out_control_0_propagate;
	wire [4:0] _mesh_12_9_io_out_control_0_shift;
	wire [2:0] _mesh_12_9_io_out_id_0;
	wire _mesh_12_9_io_out_last_0;
	wire _mesh_12_9_io_out_valid_0;
	wire [31:0] _mesh_12_8_io_out_a_0;
	wire [31:0] _mesh_12_8_io_out_c_0;
	wire [31:0] _mesh_12_8_io_out_b_0;
	wire _mesh_12_8_io_out_control_0_dataflow;
	wire _mesh_12_8_io_out_control_0_propagate;
	wire [4:0] _mesh_12_8_io_out_control_0_shift;
	wire [2:0] _mesh_12_8_io_out_id_0;
	wire _mesh_12_8_io_out_last_0;
	wire _mesh_12_8_io_out_valid_0;
	wire [31:0] _mesh_12_7_io_out_a_0;
	wire [31:0] _mesh_12_7_io_out_c_0;
	wire [31:0] _mesh_12_7_io_out_b_0;
	wire _mesh_12_7_io_out_control_0_dataflow;
	wire _mesh_12_7_io_out_control_0_propagate;
	wire [4:0] _mesh_12_7_io_out_control_0_shift;
	wire [2:0] _mesh_12_7_io_out_id_0;
	wire _mesh_12_7_io_out_last_0;
	wire _mesh_12_7_io_out_valid_0;
	wire [31:0] _mesh_12_6_io_out_a_0;
	wire [31:0] _mesh_12_6_io_out_c_0;
	wire [31:0] _mesh_12_6_io_out_b_0;
	wire _mesh_12_6_io_out_control_0_dataflow;
	wire _mesh_12_6_io_out_control_0_propagate;
	wire [4:0] _mesh_12_6_io_out_control_0_shift;
	wire [2:0] _mesh_12_6_io_out_id_0;
	wire _mesh_12_6_io_out_last_0;
	wire _mesh_12_6_io_out_valid_0;
	wire [31:0] _mesh_12_5_io_out_a_0;
	wire [31:0] _mesh_12_5_io_out_c_0;
	wire [31:0] _mesh_12_5_io_out_b_0;
	wire _mesh_12_5_io_out_control_0_dataflow;
	wire _mesh_12_5_io_out_control_0_propagate;
	wire [4:0] _mesh_12_5_io_out_control_0_shift;
	wire [2:0] _mesh_12_5_io_out_id_0;
	wire _mesh_12_5_io_out_last_0;
	wire _mesh_12_5_io_out_valid_0;
	wire [31:0] _mesh_12_4_io_out_a_0;
	wire [31:0] _mesh_12_4_io_out_c_0;
	wire [31:0] _mesh_12_4_io_out_b_0;
	wire _mesh_12_4_io_out_control_0_dataflow;
	wire _mesh_12_4_io_out_control_0_propagate;
	wire [4:0] _mesh_12_4_io_out_control_0_shift;
	wire [2:0] _mesh_12_4_io_out_id_0;
	wire _mesh_12_4_io_out_last_0;
	wire _mesh_12_4_io_out_valid_0;
	wire [31:0] _mesh_12_3_io_out_a_0;
	wire [31:0] _mesh_12_3_io_out_c_0;
	wire [31:0] _mesh_12_3_io_out_b_0;
	wire _mesh_12_3_io_out_control_0_dataflow;
	wire _mesh_12_3_io_out_control_0_propagate;
	wire [4:0] _mesh_12_3_io_out_control_0_shift;
	wire [2:0] _mesh_12_3_io_out_id_0;
	wire _mesh_12_3_io_out_last_0;
	wire _mesh_12_3_io_out_valid_0;
	wire [31:0] _mesh_12_2_io_out_a_0;
	wire [31:0] _mesh_12_2_io_out_c_0;
	wire [31:0] _mesh_12_2_io_out_b_0;
	wire _mesh_12_2_io_out_control_0_dataflow;
	wire _mesh_12_2_io_out_control_0_propagate;
	wire [4:0] _mesh_12_2_io_out_control_0_shift;
	wire [2:0] _mesh_12_2_io_out_id_0;
	wire _mesh_12_2_io_out_last_0;
	wire _mesh_12_2_io_out_valid_0;
	wire [31:0] _mesh_12_1_io_out_a_0;
	wire [31:0] _mesh_12_1_io_out_c_0;
	wire [31:0] _mesh_12_1_io_out_b_0;
	wire _mesh_12_1_io_out_control_0_dataflow;
	wire _mesh_12_1_io_out_control_0_propagate;
	wire [4:0] _mesh_12_1_io_out_control_0_shift;
	wire [2:0] _mesh_12_1_io_out_id_0;
	wire _mesh_12_1_io_out_last_0;
	wire _mesh_12_1_io_out_valid_0;
	wire [31:0] _mesh_12_0_io_out_a_0;
	wire [31:0] _mesh_12_0_io_out_c_0;
	wire [31:0] _mesh_12_0_io_out_b_0;
	wire _mesh_12_0_io_out_control_0_dataflow;
	wire _mesh_12_0_io_out_control_0_propagate;
	wire [4:0] _mesh_12_0_io_out_control_0_shift;
	wire [2:0] _mesh_12_0_io_out_id_0;
	wire _mesh_12_0_io_out_last_0;
	wire _mesh_12_0_io_out_valid_0;
	wire [31:0] _mesh_11_15_io_out_a_0;
	wire [31:0] _mesh_11_15_io_out_c_0;
	wire [31:0] _mesh_11_15_io_out_b_0;
	wire _mesh_11_15_io_out_control_0_dataflow;
	wire _mesh_11_15_io_out_control_0_propagate;
	wire [4:0] _mesh_11_15_io_out_control_0_shift;
	wire [2:0] _mesh_11_15_io_out_id_0;
	wire _mesh_11_15_io_out_last_0;
	wire _mesh_11_15_io_out_valid_0;
	wire [31:0] _mesh_11_14_io_out_a_0;
	wire [31:0] _mesh_11_14_io_out_c_0;
	wire [31:0] _mesh_11_14_io_out_b_0;
	wire _mesh_11_14_io_out_control_0_dataflow;
	wire _mesh_11_14_io_out_control_0_propagate;
	wire [4:0] _mesh_11_14_io_out_control_0_shift;
	wire [2:0] _mesh_11_14_io_out_id_0;
	wire _mesh_11_14_io_out_last_0;
	wire _mesh_11_14_io_out_valid_0;
	wire [31:0] _mesh_11_13_io_out_a_0;
	wire [31:0] _mesh_11_13_io_out_c_0;
	wire [31:0] _mesh_11_13_io_out_b_0;
	wire _mesh_11_13_io_out_control_0_dataflow;
	wire _mesh_11_13_io_out_control_0_propagate;
	wire [4:0] _mesh_11_13_io_out_control_0_shift;
	wire [2:0] _mesh_11_13_io_out_id_0;
	wire _mesh_11_13_io_out_last_0;
	wire _mesh_11_13_io_out_valid_0;
	wire [31:0] _mesh_11_12_io_out_a_0;
	wire [31:0] _mesh_11_12_io_out_c_0;
	wire [31:0] _mesh_11_12_io_out_b_0;
	wire _mesh_11_12_io_out_control_0_dataflow;
	wire _mesh_11_12_io_out_control_0_propagate;
	wire [4:0] _mesh_11_12_io_out_control_0_shift;
	wire [2:0] _mesh_11_12_io_out_id_0;
	wire _mesh_11_12_io_out_last_0;
	wire _mesh_11_12_io_out_valid_0;
	wire [31:0] _mesh_11_11_io_out_a_0;
	wire [31:0] _mesh_11_11_io_out_c_0;
	wire [31:0] _mesh_11_11_io_out_b_0;
	wire _mesh_11_11_io_out_control_0_dataflow;
	wire _mesh_11_11_io_out_control_0_propagate;
	wire [4:0] _mesh_11_11_io_out_control_0_shift;
	wire [2:0] _mesh_11_11_io_out_id_0;
	wire _mesh_11_11_io_out_last_0;
	wire _mesh_11_11_io_out_valid_0;
	wire [31:0] _mesh_11_10_io_out_a_0;
	wire [31:0] _mesh_11_10_io_out_c_0;
	wire [31:0] _mesh_11_10_io_out_b_0;
	wire _mesh_11_10_io_out_control_0_dataflow;
	wire _mesh_11_10_io_out_control_0_propagate;
	wire [4:0] _mesh_11_10_io_out_control_0_shift;
	wire [2:0] _mesh_11_10_io_out_id_0;
	wire _mesh_11_10_io_out_last_0;
	wire _mesh_11_10_io_out_valid_0;
	wire [31:0] _mesh_11_9_io_out_a_0;
	wire [31:0] _mesh_11_9_io_out_c_0;
	wire [31:0] _mesh_11_9_io_out_b_0;
	wire _mesh_11_9_io_out_control_0_dataflow;
	wire _mesh_11_9_io_out_control_0_propagate;
	wire [4:0] _mesh_11_9_io_out_control_0_shift;
	wire [2:0] _mesh_11_9_io_out_id_0;
	wire _mesh_11_9_io_out_last_0;
	wire _mesh_11_9_io_out_valid_0;
	wire [31:0] _mesh_11_8_io_out_a_0;
	wire [31:0] _mesh_11_8_io_out_c_0;
	wire [31:0] _mesh_11_8_io_out_b_0;
	wire _mesh_11_8_io_out_control_0_dataflow;
	wire _mesh_11_8_io_out_control_0_propagate;
	wire [4:0] _mesh_11_8_io_out_control_0_shift;
	wire [2:0] _mesh_11_8_io_out_id_0;
	wire _mesh_11_8_io_out_last_0;
	wire _mesh_11_8_io_out_valid_0;
	wire [31:0] _mesh_11_7_io_out_a_0;
	wire [31:0] _mesh_11_7_io_out_c_0;
	wire [31:0] _mesh_11_7_io_out_b_0;
	wire _mesh_11_7_io_out_control_0_dataflow;
	wire _mesh_11_7_io_out_control_0_propagate;
	wire [4:0] _mesh_11_7_io_out_control_0_shift;
	wire [2:0] _mesh_11_7_io_out_id_0;
	wire _mesh_11_7_io_out_last_0;
	wire _mesh_11_7_io_out_valid_0;
	wire [31:0] _mesh_11_6_io_out_a_0;
	wire [31:0] _mesh_11_6_io_out_c_0;
	wire [31:0] _mesh_11_6_io_out_b_0;
	wire _mesh_11_6_io_out_control_0_dataflow;
	wire _mesh_11_6_io_out_control_0_propagate;
	wire [4:0] _mesh_11_6_io_out_control_0_shift;
	wire [2:0] _mesh_11_6_io_out_id_0;
	wire _mesh_11_6_io_out_last_0;
	wire _mesh_11_6_io_out_valid_0;
	wire [31:0] _mesh_11_5_io_out_a_0;
	wire [31:0] _mesh_11_5_io_out_c_0;
	wire [31:0] _mesh_11_5_io_out_b_0;
	wire _mesh_11_5_io_out_control_0_dataflow;
	wire _mesh_11_5_io_out_control_0_propagate;
	wire [4:0] _mesh_11_5_io_out_control_0_shift;
	wire [2:0] _mesh_11_5_io_out_id_0;
	wire _mesh_11_5_io_out_last_0;
	wire _mesh_11_5_io_out_valid_0;
	wire [31:0] _mesh_11_4_io_out_a_0;
	wire [31:0] _mesh_11_4_io_out_c_0;
	wire [31:0] _mesh_11_4_io_out_b_0;
	wire _mesh_11_4_io_out_control_0_dataflow;
	wire _mesh_11_4_io_out_control_0_propagate;
	wire [4:0] _mesh_11_4_io_out_control_0_shift;
	wire [2:0] _mesh_11_4_io_out_id_0;
	wire _mesh_11_4_io_out_last_0;
	wire _mesh_11_4_io_out_valid_0;
	wire [31:0] _mesh_11_3_io_out_a_0;
	wire [31:0] _mesh_11_3_io_out_c_0;
	wire [31:0] _mesh_11_3_io_out_b_0;
	wire _mesh_11_3_io_out_control_0_dataflow;
	wire _mesh_11_3_io_out_control_0_propagate;
	wire [4:0] _mesh_11_3_io_out_control_0_shift;
	wire [2:0] _mesh_11_3_io_out_id_0;
	wire _mesh_11_3_io_out_last_0;
	wire _mesh_11_3_io_out_valid_0;
	wire [31:0] _mesh_11_2_io_out_a_0;
	wire [31:0] _mesh_11_2_io_out_c_0;
	wire [31:0] _mesh_11_2_io_out_b_0;
	wire _mesh_11_2_io_out_control_0_dataflow;
	wire _mesh_11_2_io_out_control_0_propagate;
	wire [4:0] _mesh_11_2_io_out_control_0_shift;
	wire [2:0] _mesh_11_2_io_out_id_0;
	wire _mesh_11_2_io_out_last_0;
	wire _mesh_11_2_io_out_valid_0;
	wire [31:0] _mesh_11_1_io_out_a_0;
	wire [31:0] _mesh_11_1_io_out_c_0;
	wire [31:0] _mesh_11_1_io_out_b_0;
	wire _mesh_11_1_io_out_control_0_dataflow;
	wire _mesh_11_1_io_out_control_0_propagate;
	wire [4:0] _mesh_11_1_io_out_control_0_shift;
	wire [2:0] _mesh_11_1_io_out_id_0;
	wire _mesh_11_1_io_out_last_0;
	wire _mesh_11_1_io_out_valid_0;
	wire [31:0] _mesh_11_0_io_out_a_0;
	wire [31:0] _mesh_11_0_io_out_c_0;
	wire [31:0] _mesh_11_0_io_out_b_0;
	wire _mesh_11_0_io_out_control_0_dataflow;
	wire _mesh_11_0_io_out_control_0_propagate;
	wire [4:0] _mesh_11_0_io_out_control_0_shift;
	wire [2:0] _mesh_11_0_io_out_id_0;
	wire _mesh_11_0_io_out_last_0;
	wire _mesh_11_0_io_out_valid_0;
	wire [31:0] _mesh_10_15_io_out_a_0;
	wire [31:0] _mesh_10_15_io_out_c_0;
	wire [31:0] _mesh_10_15_io_out_b_0;
	wire _mesh_10_15_io_out_control_0_dataflow;
	wire _mesh_10_15_io_out_control_0_propagate;
	wire [4:0] _mesh_10_15_io_out_control_0_shift;
	wire [2:0] _mesh_10_15_io_out_id_0;
	wire _mesh_10_15_io_out_last_0;
	wire _mesh_10_15_io_out_valid_0;
	wire [31:0] _mesh_10_14_io_out_a_0;
	wire [31:0] _mesh_10_14_io_out_c_0;
	wire [31:0] _mesh_10_14_io_out_b_0;
	wire _mesh_10_14_io_out_control_0_dataflow;
	wire _mesh_10_14_io_out_control_0_propagate;
	wire [4:0] _mesh_10_14_io_out_control_0_shift;
	wire [2:0] _mesh_10_14_io_out_id_0;
	wire _mesh_10_14_io_out_last_0;
	wire _mesh_10_14_io_out_valid_0;
	wire [31:0] _mesh_10_13_io_out_a_0;
	wire [31:0] _mesh_10_13_io_out_c_0;
	wire [31:0] _mesh_10_13_io_out_b_0;
	wire _mesh_10_13_io_out_control_0_dataflow;
	wire _mesh_10_13_io_out_control_0_propagate;
	wire [4:0] _mesh_10_13_io_out_control_0_shift;
	wire [2:0] _mesh_10_13_io_out_id_0;
	wire _mesh_10_13_io_out_last_0;
	wire _mesh_10_13_io_out_valid_0;
	wire [31:0] _mesh_10_12_io_out_a_0;
	wire [31:0] _mesh_10_12_io_out_c_0;
	wire [31:0] _mesh_10_12_io_out_b_0;
	wire _mesh_10_12_io_out_control_0_dataflow;
	wire _mesh_10_12_io_out_control_0_propagate;
	wire [4:0] _mesh_10_12_io_out_control_0_shift;
	wire [2:0] _mesh_10_12_io_out_id_0;
	wire _mesh_10_12_io_out_last_0;
	wire _mesh_10_12_io_out_valid_0;
	wire [31:0] _mesh_10_11_io_out_a_0;
	wire [31:0] _mesh_10_11_io_out_c_0;
	wire [31:0] _mesh_10_11_io_out_b_0;
	wire _mesh_10_11_io_out_control_0_dataflow;
	wire _mesh_10_11_io_out_control_0_propagate;
	wire [4:0] _mesh_10_11_io_out_control_0_shift;
	wire [2:0] _mesh_10_11_io_out_id_0;
	wire _mesh_10_11_io_out_last_0;
	wire _mesh_10_11_io_out_valid_0;
	wire [31:0] _mesh_10_10_io_out_a_0;
	wire [31:0] _mesh_10_10_io_out_c_0;
	wire [31:0] _mesh_10_10_io_out_b_0;
	wire _mesh_10_10_io_out_control_0_dataflow;
	wire _mesh_10_10_io_out_control_0_propagate;
	wire [4:0] _mesh_10_10_io_out_control_0_shift;
	wire [2:0] _mesh_10_10_io_out_id_0;
	wire _mesh_10_10_io_out_last_0;
	wire _mesh_10_10_io_out_valid_0;
	wire [31:0] _mesh_10_9_io_out_a_0;
	wire [31:0] _mesh_10_9_io_out_c_0;
	wire [31:0] _mesh_10_9_io_out_b_0;
	wire _mesh_10_9_io_out_control_0_dataflow;
	wire _mesh_10_9_io_out_control_0_propagate;
	wire [4:0] _mesh_10_9_io_out_control_0_shift;
	wire [2:0] _mesh_10_9_io_out_id_0;
	wire _mesh_10_9_io_out_last_0;
	wire _mesh_10_9_io_out_valid_0;
	wire [31:0] _mesh_10_8_io_out_a_0;
	wire [31:0] _mesh_10_8_io_out_c_0;
	wire [31:0] _mesh_10_8_io_out_b_0;
	wire _mesh_10_8_io_out_control_0_dataflow;
	wire _mesh_10_8_io_out_control_0_propagate;
	wire [4:0] _mesh_10_8_io_out_control_0_shift;
	wire [2:0] _mesh_10_8_io_out_id_0;
	wire _mesh_10_8_io_out_last_0;
	wire _mesh_10_8_io_out_valid_0;
	wire [31:0] _mesh_10_7_io_out_a_0;
	wire [31:0] _mesh_10_7_io_out_c_0;
	wire [31:0] _mesh_10_7_io_out_b_0;
	wire _mesh_10_7_io_out_control_0_dataflow;
	wire _mesh_10_7_io_out_control_0_propagate;
	wire [4:0] _mesh_10_7_io_out_control_0_shift;
	wire [2:0] _mesh_10_7_io_out_id_0;
	wire _mesh_10_7_io_out_last_0;
	wire _mesh_10_7_io_out_valid_0;
	wire [31:0] _mesh_10_6_io_out_a_0;
	wire [31:0] _mesh_10_6_io_out_c_0;
	wire [31:0] _mesh_10_6_io_out_b_0;
	wire _mesh_10_6_io_out_control_0_dataflow;
	wire _mesh_10_6_io_out_control_0_propagate;
	wire [4:0] _mesh_10_6_io_out_control_0_shift;
	wire [2:0] _mesh_10_6_io_out_id_0;
	wire _mesh_10_6_io_out_last_0;
	wire _mesh_10_6_io_out_valid_0;
	wire [31:0] _mesh_10_5_io_out_a_0;
	wire [31:0] _mesh_10_5_io_out_c_0;
	wire [31:0] _mesh_10_5_io_out_b_0;
	wire _mesh_10_5_io_out_control_0_dataflow;
	wire _mesh_10_5_io_out_control_0_propagate;
	wire [4:0] _mesh_10_5_io_out_control_0_shift;
	wire [2:0] _mesh_10_5_io_out_id_0;
	wire _mesh_10_5_io_out_last_0;
	wire _mesh_10_5_io_out_valid_0;
	wire [31:0] _mesh_10_4_io_out_a_0;
	wire [31:0] _mesh_10_4_io_out_c_0;
	wire [31:0] _mesh_10_4_io_out_b_0;
	wire _mesh_10_4_io_out_control_0_dataflow;
	wire _mesh_10_4_io_out_control_0_propagate;
	wire [4:0] _mesh_10_4_io_out_control_0_shift;
	wire [2:0] _mesh_10_4_io_out_id_0;
	wire _mesh_10_4_io_out_last_0;
	wire _mesh_10_4_io_out_valid_0;
	wire [31:0] _mesh_10_3_io_out_a_0;
	wire [31:0] _mesh_10_3_io_out_c_0;
	wire [31:0] _mesh_10_3_io_out_b_0;
	wire _mesh_10_3_io_out_control_0_dataflow;
	wire _mesh_10_3_io_out_control_0_propagate;
	wire [4:0] _mesh_10_3_io_out_control_0_shift;
	wire [2:0] _mesh_10_3_io_out_id_0;
	wire _mesh_10_3_io_out_last_0;
	wire _mesh_10_3_io_out_valid_0;
	wire [31:0] _mesh_10_2_io_out_a_0;
	wire [31:0] _mesh_10_2_io_out_c_0;
	wire [31:0] _mesh_10_2_io_out_b_0;
	wire _mesh_10_2_io_out_control_0_dataflow;
	wire _mesh_10_2_io_out_control_0_propagate;
	wire [4:0] _mesh_10_2_io_out_control_0_shift;
	wire [2:0] _mesh_10_2_io_out_id_0;
	wire _mesh_10_2_io_out_last_0;
	wire _mesh_10_2_io_out_valid_0;
	wire [31:0] _mesh_10_1_io_out_a_0;
	wire [31:0] _mesh_10_1_io_out_c_0;
	wire [31:0] _mesh_10_1_io_out_b_0;
	wire _mesh_10_1_io_out_control_0_dataflow;
	wire _mesh_10_1_io_out_control_0_propagate;
	wire [4:0] _mesh_10_1_io_out_control_0_shift;
	wire [2:0] _mesh_10_1_io_out_id_0;
	wire _mesh_10_1_io_out_last_0;
	wire _mesh_10_1_io_out_valid_0;
	wire [31:0] _mesh_10_0_io_out_a_0;
	wire [31:0] _mesh_10_0_io_out_c_0;
	wire [31:0] _mesh_10_0_io_out_b_0;
	wire _mesh_10_0_io_out_control_0_dataflow;
	wire _mesh_10_0_io_out_control_0_propagate;
	wire [4:0] _mesh_10_0_io_out_control_0_shift;
	wire [2:0] _mesh_10_0_io_out_id_0;
	wire _mesh_10_0_io_out_last_0;
	wire _mesh_10_0_io_out_valid_0;
	wire [31:0] _mesh_9_15_io_out_a_0;
	wire [31:0] _mesh_9_15_io_out_c_0;
	wire [31:0] _mesh_9_15_io_out_b_0;
	wire _mesh_9_15_io_out_control_0_dataflow;
	wire _mesh_9_15_io_out_control_0_propagate;
	wire [4:0] _mesh_9_15_io_out_control_0_shift;
	wire [2:0] _mesh_9_15_io_out_id_0;
	wire _mesh_9_15_io_out_last_0;
	wire _mesh_9_15_io_out_valid_0;
	wire [31:0] _mesh_9_14_io_out_a_0;
	wire [31:0] _mesh_9_14_io_out_c_0;
	wire [31:0] _mesh_9_14_io_out_b_0;
	wire _mesh_9_14_io_out_control_0_dataflow;
	wire _mesh_9_14_io_out_control_0_propagate;
	wire [4:0] _mesh_9_14_io_out_control_0_shift;
	wire [2:0] _mesh_9_14_io_out_id_0;
	wire _mesh_9_14_io_out_last_0;
	wire _mesh_9_14_io_out_valid_0;
	wire [31:0] _mesh_9_13_io_out_a_0;
	wire [31:0] _mesh_9_13_io_out_c_0;
	wire [31:0] _mesh_9_13_io_out_b_0;
	wire _mesh_9_13_io_out_control_0_dataflow;
	wire _mesh_9_13_io_out_control_0_propagate;
	wire [4:0] _mesh_9_13_io_out_control_0_shift;
	wire [2:0] _mesh_9_13_io_out_id_0;
	wire _mesh_9_13_io_out_last_0;
	wire _mesh_9_13_io_out_valid_0;
	wire [31:0] _mesh_9_12_io_out_a_0;
	wire [31:0] _mesh_9_12_io_out_c_0;
	wire [31:0] _mesh_9_12_io_out_b_0;
	wire _mesh_9_12_io_out_control_0_dataflow;
	wire _mesh_9_12_io_out_control_0_propagate;
	wire [4:0] _mesh_9_12_io_out_control_0_shift;
	wire [2:0] _mesh_9_12_io_out_id_0;
	wire _mesh_9_12_io_out_last_0;
	wire _mesh_9_12_io_out_valid_0;
	wire [31:0] _mesh_9_11_io_out_a_0;
	wire [31:0] _mesh_9_11_io_out_c_0;
	wire [31:0] _mesh_9_11_io_out_b_0;
	wire _mesh_9_11_io_out_control_0_dataflow;
	wire _mesh_9_11_io_out_control_0_propagate;
	wire [4:0] _mesh_9_11_io_out_control_0_shift;
	wire [2:0] _mesh_9_11_io_out_id_0;
	wire _mesh_9_11_io_out_last_0;
	wire _mesh_9_11_io_out_valid_0;
	wire [31:0] _mesh_9_10_io_out_a_0;
	wire [31:0] _mesh_9_10_io_out_c_0;
	wire [31:0] _mesh_9_10_io_out_b_0;
	wire _mesh_9_10_io_out_control_0_dataflow;
	wire _mesh_9_10_io_out_control_0_propagate;
	wire [4:0] _mesh_9_10_io_out_control_0_shift;
	wire [2:0] _mesh_9_10_io_out_id_0;
	wire _mesh_9_10_io_out_last_0;
	wire _mesh_9_10_io_out_valid_0;
	wire [31:0] _mesh_9_9_io_out_a_0;
	wire [31:0] _mesh_9_9_io_out_c_0;
	wire [31:0] _mesh_9_9_io_out_b_0;
	wire _mesh_9_9_io_out_control_0_dataflow;
	wire _mesh_9_9_io_out_control_0_propagate;
	wire [4:0] _mesh_9_9_io_out_control_0_shift;
	wire [2:0] _mesh_9_9_io_out_id_0;
	wire _mesh_9_9_io_out_last_0;
	wire _mesh_9_9_io_out_valid_0;
	wire [31:0] _mesh_9_8_io_out_a_0;
	wire [31:0] _mesh_9_8_io_out_c_0;
	wire [31:0] _mesh_9_8_io_out_b_0;
	wire _mesh_9_8_io_out_control_0_dataflow;
	wire _mesh_9_8_io_out_control_0_propagate;
	wire [4:0] _mesh_9_8_io_out_control_0_shift;
	wire [2:0] _mesh_9_8_io_out_id_0;
	wire _mesh_9_8_io_out_last_0;
	wire _mesh_9_8_io_out_valid_0;
	wire [31:0] _mesh_9_7_io_out_a_0;
	wire [31:0] _mesh_9_7_io_out_c_0;
	wire [31:0] _mesh_9_7_io_out_b_0;
	wire _mesh_9_7_io_out_control_0_dataflow;
	wire _mesh_9_7_io_out_control_0_propagate;
	wire [4:0] _mesh_9_7_io_out_control_0_shift;
	wire [2:0] _mesh_9_7_io_out_id_0;
	wire _mesh_9_7_io_out_last_0;
	wire _mesh_9_7_io_out_valid_0;
	wire [31:0] _mesh_9_6_io_out_a_0;
	wire [31:0] _mesh_9_6_io_out_c_0;
	wire [31:0] _mesh_9_6_io_out_b_0;
	wire _mesh_9_6_io_out_control_0_dataflow;
	wire _mesh_9_6_io_out_control_0_propagate;
	wire [4:0] _mesh_9_6_io_out_control_0_shift;
	wire [2:0] _mesh_9_6_io_out_id_0;
	wire _mesh_9_6_io_out_last_0;
	wire _mesh_9_6_io_out_valid_0;
	wire [31:0] _mesh_9_5_io_out_a_0;
	wire [31:0] _mesh_9_5_io_out_c_0;
	wire [31:0] _mesh_9_5_io_out_b_0;
	wire _mesh_9_5_io_out_control_0_dataflow;
	wire _mesh_9_5_io_out_control_0_propagate;
	wire [4:0] _mesh_9_5_io_out_control_0_shift;
	wire [2:0] _mesh_9_5_io_out_id_0;
	wire _mesh_9_5_io_out_last_0;
	wire _mesh_9_5_io_out_valid_0;
	wire [31:0] _mesh_9_4_io_out_a_0;
	wire [31:0] _mesh_9_4_io_out_c_0;
	wire [31:0] _mesh_9_4_io_out_b_0;
	wire _mesh_9_4_io_out_control_0_dataflow;
	wire _mesh_9_4_io_out_control_0_propagate;
	wire [4:0] _mesh_9_4_io_out_control_0_shift;
	wire [2:0] _mesh_9_4_io_out_id_0;
	wire _mesh_9_4_io_out_last_0;
	wire _mesh_9_4_io_out_valid_0;
	wire [31:0] _mesh_9_3_io_out_a_0;
	wire [31:0] _mesh_9_3_io_out_c_0;
	wire [31:0] _mesh_9_3_io_out_b_0;
	wire _mesh_9_3_io_out_control_0_dataflow;
	wire _mesh_9_3_io_out_control_0_propagate;
	wire [4:0] _mesh_9_3_io_out_control_0_shift;
	wire [2:0] _mesh_9_3_io_out_id_0;
	wire _mesh_9_3_io_out_last_0;
	wire _mesh_9_3_io_out_valid_0;
	wire [31:0] _mesh_9_2_io_out_a_0;
	wire [31:0] _mesh_9_2_io_out_c_0;
	wire [31:0] _mesh_9_2_io_out_b_0;
	wire _mesh_9_2_io_out_control_0_dataflow;
	wire _mesh_9_2_io_out_control_0_propagate;
	wire [4:0] _mesh_9_2_io_out_control_0_shift;
	wire [2:0] _mesh_9_2_io_out_id_0;
	wire _mesh_9_2_io_out_last_0;
	wire _mesh_9_2_io_out_valid_0;
	wire [31:0] _mesh_9_1_io_out_a_0;
	wire [31:0] _mesh_9_1_io_out_c_0;
	wire [31:0] _mesh_9_1_io_out_b_0;
	wire _mesh_9_1_io_out_control_0_dataflow;
	wire _mesh_9_1_io_out_control_0_propagate;
	wire [4:0] _mesh_9_1_io_out_control_0_shift;
	wire [2:0] _mesh_9_1_io_out_id_0;
	wire _mesh_9_1_io_out_last_0;
	wire _mesh_9_1_io_out_valid_0;
	wire [31:0] _mesh_9_0_io_out_a_0;
	wire [31:0] _mesh_9_0_io_out_c_0;
	wire [31:0] _mesh_9_0_io_out_b_0;
	wire _mesh_9_0_io_out_control_0_dataflow;
	wire _mesh_9_0_io_out_control_0_propagate;
	wire [4:0] _mesh_9_0_io_out_control_0_shift;
	wire [2:0] _mesh_9_0_io_out_id_0;
	wire _mesh_9_0_io_out_last_0;
	wire _mesh_9_0_io_out_valid_0;
	wire [31:0] _mesh_8_15_io_out_a_0;
	wire [31:0] _mesh_8_15_io_out_c_0;
	wire [31:0] _mesh_8_15_io_out_b_0;
	wire _mesh_8_15_io_out_control_0_dataflow;
	wire _mesh_8_15_io_out_control_0_propagate;
	wire [4:0] _mesh_8_15_io_out_control_0_shift;
	wire [2:0] _mesh_8_15_io_out_id_0;
	wire _mesh_8_15_io_out_last_0;
	wire _mesh_8_15_io_out_valid_0;
	wire [31:0] _mesh_8_14_io_out_a_0;
	wire [31:0] _mesh_8_14_io_out_c_0;
	wire [31:0] _mesh_8_14_io_out_b_0;
	wire _mesh_8_14_io_out_control_0_dataflow;
	wire _mesh_8_14_io_out_control_0_propagate;
	wire [4:0] _mesh_8_14_io_out_control_0_shift;
	wire [2:0] _mesh_8_14_io_out_id_0;
	wire _mesh_8_14_io_out_last_0;
	wire _mesh_8_14_io_out_valid_0;
	wire [31:0] _mesh_8_13_io_out_a_0;
	wire [31:0] _mesh_8_13_io_out_c_0;
	wire [31:0] _mesh_8_13_io_out_b_0;
	wire _mesh_8_13_io_out_control_0_dataflow;
	wire _mesh_8_13_io_out_control_0_propagate;
	wire [4:0] _mesh_8_13_io_out_control_0_shift;
	wire [2:0] _mesh_8_13_io_out_id_0;
	wire _mesh_8_13_io_out_last_0;
	wire _mesh_8_13_io_out_valid_0;
	wire [31:0] _mesh_8_12_io_out_a_0;
	wire [31:0] _mesh_8_12_io_out_c_0;
	wire [31:0] _mesh_8_12_io_out_b_0;
	wire _mesh_8_12_io_out_control_0_dataflow;
	wire _mesh_8_12_io_out_control_0_propagate;
	wire [4:0] _mesh_8_12_io_out_control_0_shift;
	wire [2:0] _mesh_8_12_io_out_id_0;
	wire _mesh_8_12_io_out_last_0;
	wire _mesh_8_12_io_out_valid_0;
	wire [31:0] _mesh_8_11_io_out_a_0;
	wire [31:0] _mesh_8_11_io_out_c_0;
	wire [31:0] _mesh_8_11_io_out_b_0;
	wire _mesh_8_11_io_out_control_0_dataflow;
	wire _mesh_8_11_io_out_control_0_propagate;
	wire [4:0] _mesh_8_11_io_out_control_0_shift;
	wire [2:0] _mesh_8_11_io_out_id_0;
	wire _mesh_8_11_io_out_last_0;
	wire _mesh_8_11_io_out_valid_0;
	wire [31:0] _mesh_8_10_io_out_a_0;
	wire [31:0] _mesh_8_10_io_out_c_0;
	wire [31:0] _mesh_8_10_io_out_b_0;
	wire _mesh_8_10_io_out_control_0_dataflow;
	wire _mesh_8_10_io_out_control_0_propagate;
	wire [4:0] _mesh_8_10_io_out_control_0_shift;
	wire [2:0] _mesh_8_10_io_out_id_0;
	wire _mesh_8_10_io_out_last_0;
	wire _mesh_8_10_io_out_valid_0;
	wire [31:0] _mesh_8_9_io_out_a_0;
	wire [31:0] _mesh_8_9_io_out_c_0;
	wire [31:0] _mesh_8_9_io_out_b_0;
	wire _mesh_8_9_io_out_control_0_dataflow;
	wire _mesh_8_9_io_out_control_0_propagate;
	wire [4:0] _mesh_8_9_io_out_control_0_shift;
	wire [2:0] _mesh_8_9_io_out_id_0;
	wire _mesh_8_9_io_out_last_0;
	wire _mesh_8_9_io_out_valid_0;
	wire [31:0] _mesh_8_8_io_out_a_0;
	wire [31:0] _mesh_8_8_io_out_c_0;
	wire [31:0] _mesh_8_8_io_out_b_0;
	wire _mesh_8_8_io_out_control_0_dataflow;
	wire _mesh_8_8_io_out_control_0_propagate;
	wire [4:0] _mesh_8_8_io_out_control_0_shift;
	wire [2:0] _mesh_8_8_io_out_id_0;
	wire _mesh_8_8_io_out_last_0;
	wire _mesh_8_8_io_out_valid_0;
	wire [31:0] _mesh_8_7_io_out_a_0;
	wire [31:0] _mesh_8_7_io_out_c_0;
	wire [31:0] _mesh_8_7_io_out_b_0;
	wire _mesh_8_7_io_out_control_0_dataflow;
	wire _mesh_8_7_io_out_control_0_propagate;
	wire [4:0] _mesh_8_7_io_out_control_0_shift;
	wire [2:0] _mesh_8_7_io_out_id_0;
	wire _mesh_8_7_io_out_last_0;
	wire _mesh_8_7_io_out_valid_0;
	wire [31:0] _mesh_8_6_io_out_a_0;
	wire [31:0] _mesh_8_6_io_out_c_0;
	wire [31:0] _mesh_8_6_io_out_b_0;
	wire _mesh_8_6_io_out_control_0_dataflow;
	wire _mesh_8_6_io_out_control_0_propagate;
	wire [4:0] _mesh_8_6_io_out_control_0_shift;
	wire [2:0] _mesh_8_6_io_out_id_0;
	wire _mesh_8_6_io_out_last_0;
	wire _mesh_8_6_io_out_valid_0;
	wire [31:0] _mesh_8_5_io_out_a_0;
	wire [31:0] _mesh_8_5_io_out_c_0;
	wire [31:0] _mesh_8_5_io_out_b_0;
	wire _mesh_8_5_io_out_control_0_dataflow;
	wire _mesh_8_5_io_out_control_0_propagate;
	wire [4:0] _mesh_8_5_io_out_control_0_shift;
	wire [2:0] _mesh_8_5_io_out_id_0;
	wire _mesh_8_5_io_out_last_0;
	wire _mesh_8_5_io_out_valid_0;
	wire [31:0] _mesh_8_4_io_out_a_0;
	wire [31:0] _mesh_8_4_io_out_c_0;
	wire [31:0] _mesh_8_4_io_out_b_0;
	wire _mesh_8_4_io_out_control_0_dataflow;
	wire _mesh_8_4_io_out_control_0_propagate;
	wire [4:0] _mesh_8_4_io_out_control_0_shift;
	wire [2:0] _mesh_8_4_io_out_id_0;
	wire _mesh_8_4_io_out_last_0;
	wire _mesh_8_4_io_out_valid_0;
	wire [31:0] _mesh_8_3_io_out_a_0;
	wire [31:0] _mesh_8_3_io_out_c_0;
	wire [31:0] _mesh_8_3_io_out_b_0;
	wire _mesh_8_3_io_out_control_0_dataflow;
	wire _mesh_8_3_io_out_control_0_propagate;
	wire [4:0] _mesh_8_3_io_out_control_0_shift;
	wire [2:0] _mesh_8_3_io_out_id_0;
	wire _mesh_8_3_io_out_last_0;
	wire _mesh_8_3_io_out_valid_0;
	wire [31:0] _mesh_8_2_io_out_a_0;
	wire [31:0] _mesh_8_2_io_out_c_0;
	wire [31:0] _mesh_8_2_io_out_b_0;
	wire _mesh_8_2_io_out_control_0_dataflow;
	wire _mesh_8_2_io_out_control_0_propagate;
	wire [4:0] _mesh_8_2_io_out_control_0_shift;
	wire [2:0] _mesh_8_2_io_out_id_0;
	wire _mesh_8_2_io_out_last_0;
	wire _mesh_8_2_io_out_valid_0;
	wire [31:0] _mesh_8_1_io_out_a_0;
	wire [31:0] _mesh_8_1_io_out_c_0;
	wire [31:0] _mesh_8_1_io_out_b_0;
	wire _mesh_8_1_io_out_control_0_dataflow;
	wire _mesh_8_1_io_out_control_0_propagate;
	wire [4:0] _mesh_8_1_io_out_control_0_shift;
	wire [2:0] _mesh_8_1_io_out_id_0;
	wire _mesh_8_1_io_out_last_0;
	wire _mesh_8_1_io_out_valid_0;
	wire [31:0] _mesh_8_0_io_out_a_0;
	wire [31:0] _mesh_8_0_io_out_c_0;
	wire [31:0] _mesh_8_0_io_out_b_0;
	wire _mesh_8_0_io_out_control_0_dataflow;
	wire _mesh_8_0_io_out_control_0_propagate;
	wire [4:0] _mesh_8_0_io_out_control_0_shift;
	wire [2:0] _mesh_8_0_io_out_id_0;
	wire _mesh_8_0_io_out_last_0;
	wire _mesh_8_0_io_out_valid_0;
	wire [31:0] _mesh_7_15_io_out_a_0;
	wire [31:0] _mesh_7_15_io_out_c_0;
	wire [31:0] _mesh_7_15_io_out_b_0;
	wire _mesh_7_15_io_out_control_0_dataflow;
	wire _mesh_7_15_io_out_control_0_propagate;
	wire [4:0] _mesh_7_15_io_out_control_0_shift;
	wire [2:0] _mesh_7_15_io_out_id_0;
	wire _mesh_7_15_io_out_last_0;
	wire _mesh_7_15_io_out_valid_0;
	wire [31:0] _mesh_7_14_io_out_a_0;
	wire [31:0] _mesh_7_14_io_out_c_0;
	wire [31:0] _mesh_7_14_io_out_b_0;
	wire _mesh_7_14_io_out_control_0_dataflow;
	wire _mesh_7_14_io_out_control_0_propagate;
	wire [4:0] _mesh_7_14_io_out_control_0_shift;
	wire [2:0] _mesh_7_14_io_out_id_0;
	wire _mesh_7_14_io_out_last_0;
	wire _mesh_7_14_io_out_valid_0;
	wire [31:0] _mesh_7_13_io_out_a_0;
	wire [31:0] _mesh_7_13_io_out_c_0;
	wire [31:0] _mesh_7_13_io_out_b_0;
	wire _mesh_7_13_io_out_control_0_dataflow;
	wire _mesh_7_13_io_out_control_0_propagate;
	wire [4:0] _mesh_7_13_io_out_control_0_shift;
	wire [2:0] _mesh_7_13_io_out_id_0;
	wire _mesh_7_13_io_out_last_0;
	wire _mesh_7_13_io_out_valid_0;
	wire [31:0] _mesh_7_12_io_out_a_0;
	wire [31:0] _mesh_7_12_io_out_c_0;
	wire [31:0] _mesh_7_12_io_out_b_0;
	wire _mesh_7_12_io_out_control_0_dataflow;
	wire _mesh_7_12_io_out_control_0_propagate;
	wire [4:0] _mesh_7_12_io_out_control_0_shift;
	wire [2:0] _mesh_7_12_io_out_id_0;
	wire _mesh_7_12_io_out_last_0;
	wire _mesh_7_12_io_out_valid_0;
	wire [31:0] _mesh_7_11_io_out_a_0;
	wire [31:0] _mesh_7_11_io_out_c_0;
	wire [31:0] _mesh_7_11_io_out_b_0;
	wire _mesh_7_11_io_out_control_0_dataflow;
	wire _mesh_7_11_io_out_control_0_propagate;
	wire [4:0] _mesh_7_11_io_out_control_0_shift;
	wire [2:0] _mesh_7_11_io_out_id_0;
	wire _mesh_7_11_io_out_last_0;
	wire _mesh_7_11_io_out_valid_0;
	wire [31:0] _mesh_7_10_io_out_a_0;
	wire [31:0] _mesh_7_10_io_out_c_0;
	wire [31:0] _mesh_7_10_io_out_b_0;
	wire _mesh_7_10_io_out_control_0_dataflow;
	wire _mesh_7_10_io_out_control_0_propagate;
	wire [4:0] _mesh_7_10_io_out_control_0_shift;
	wire [2:0] _mesh_7_10_io_out_id_0;
	wire _mesh_7_10_io_out_last_0;
	wire _mesh_7_10_io_out_valid_0;
	wire [31:0] _mesh_7_9_io_out_a_0;
	wire [31:0] _mesh_7_9_io_out_c_0;
	wire [31:0] _mesh_7_9_io_out_b_0;
	wire _mesh_7_9_io_out_control_0_dataflow;
	wire _mesh_7_9_io_out_control_0_propagate;
	wire [4:0] _mesh_7_9_io_out_control_0_shift;
	wire [2:0] _mesh_7_9_io_out_id_0;
	wire _mesh_7_9_io_out_last_0;
	wire _mesh_7_9_io_out_valid_0;
	wire [31:0] _mesh_7_8_io_out_a_0;
	wire [31:0] _mesh_7_8_io_out_c_0;
	wire [31:0] _mesh_7_8_io_out_b_0;
	wire _mesh_7_8_io_out_control_0_dataflow;
	wire _mesh_7_8_io_out_control_0_propagate;
	wire [4:0] _mesh_7_8_io_out_control_0_shift;
	wire [2:0] _mesh_7_8_io_out_id_0;
	wire _mesh_7_8_io_out_last_0;
	wire _mesh_7_8_io_out_valid_0;
	wire [31:0] _mesh_7_7_io_out_a_0;
	wire [31:0] _mesh_7_7_io_out_c_0;
	wire [31:0] _mesh_7_7_io_out_b_0;
	wire _mesh_7_7_io_out_control_0_dataflow;
	wire _mesh_7_7_io_out_control_0_propagate;
	wire [4:0] _mesh_7_7_io_out_control_0_shift;
	wire [2:0] _mesh_7_7_io_out_id_0;
	wire _mesh_7_7_io_out_last_0;
	wire _mesh_7_7_io_out_valid_0;
	wire [31:0] _mesh_7_6_io_out_a_0;
	wire [31:0] _mesh_7_6_io_out_c_0;
	wire [31:0] _mesh_7_6_io_out_b_0;
	wire _mesh_7_6_io_out_control_0_dataflow;
	wire _mesh_7_6_io_out_control_0_propagate;
	wire [4:0] _mesh_7_6_io_out_control_0_shift;
	wire [2:0] _mesh_7_6_io_out_id_0;
	wire _mesh_7_6_io_out_last_0;
	wire _mesh_7_6_io_out_valid_0;
	wire [31:0] _mesh_7_5_io_out_a_0;
	wire [31:0] _mesh_7_5_io_out_c_0;
	wire [31:0] _mesh_7_5_io_out_b_0;
	wire _mesh_7_5_io_out_control_0_dataflow;
	wire _mesh_7_5_io_out_control_0_propagate;
	wire [4:0] _mesh_7_5_io_out_control_0_shift;
	wire [2:0] _mesh_7_5_io_out_id_0;
	wire _mesh_7_5_io_out_last_0;
	wire _mesh_7_5_io_out_valid_0;
	wire [31:0] _mesh_7_4_io_out_a_0;
	wire [31:0] _mesh_7_4_io_out_c_0;
	wire [31:0] _mesh_7_4_io_out_b_0;
	wire _mesh_7_4_io_out_control_0_dataflow;
	wire _mesh_7_4_io_out_control_0_propagate;
	wire [4:0] _mesh_7_4_io_out_control_0_shift;
	wire [2:0] _mesh_7_4_io_out_id_0;
	wire _mesh_7_4_io_out_last_0;
	wire _mesh_7_4_io_out_valid_0;
	wire [31:0] _mesh_7_3_io_out_a_0;
	wire [31:0] _mesh_7_3_io_out_c_0;
	wire [31:0] _mesh_7_3_io_out_b_0;
	wire _mesh_7_3_io_out_control_0_dataflow;
	wire _mesh_7_3_io_out_control_0_propagate;
	wire [4:0] _mesh_7_3_io_out_control_0_shift;
	wire [2:0] _mesh_7_3_io_out_id_0;
	wire _mesh_7_3_io_out_last_0;
	wire _mesh_7_3_io_out_valid_0;
	wire [31:0] _mesh_7_2_io_out_a_0;
	wire [31:0] _mesh_7_2_io_out_c_0;
	wire [31:0] _mesh_7_2_io_out_b_0;
	wire _mesh_7_2_io_out_control_0_dataflow;
	wire _mesh_7_2_io_out_control_0_propagate;
	wire [4:0] _mesh_7_2_io_out_control_0_shift;
	wire [2:0] _mesh_7_2_io_out_id_0;
	wire _mesh_7_2_io_out_last_0;
	wire _mesh_7_2_io_out_valid_0;
	wire [31:0] _mesh_7_1_io_out_a_0;
	wire [31:0] _mesh_7_1_io_out_c_0;
	wire [31:0] _mesh_7_1_io_out_b_0;
	wire _mesh_7_1_io_out_control_0_dataflow;
	wire _mesh_7_1_io_out_control_0_propagate;
	wire [4:0] _mesh_7_1_io_out_control_0_shift;
	wire [2:0] _mesh_7_1_io_out_id_0;
	wire _mesh_7_1_io_out_last_0;
	wire _mesh_7_1_io_out_valid_0;
	wire [31:0] _mesh_7_0_io_out_a_0;
	wire [31:0] _mesh_7_0_io_out_c_0;
	wire [31:0] _mesh_7_0_io_out_b_0;
	wire _mesh_7_0_io_out_control_0_dataflow;
	wire _mesh_7_0_io_out_control_0_propagate;
	wire [4:0] _mesh_7_0_io_out_control_0_shift;
	wire [2:0] _mesh_7_0_io_out_id_0;
	wire _mesh_7_0_io_out_last_0;
	wire _mesh_7_0_io_out_valid_0;
	wire [31:0] _mesh_6_15_io_out_a_0;
	wire [31:0] _mesh_6_15_io_out_c_0;
	wire [31:0] _mesh_6_15_io_out_b_0;
	wire _mesh_6_15_io_out_control_0_dataflow;
	wire _mesh_6_15_io_out_control_0_propagate;
	wire [4:0] _mesh_6_15_io_out_control_0_shift;
	wire [2:0] _mesh_6_15_io_out_id_0;
	wire _mesh_6_15_io_out_last_0;
	wire _mesh_6_15_io_out_valid_0;
	wire [31:0] _mesh_6_14_io_out_a_0;
	wire [31:0] _mesh_6_14_io_out_c_0;
	wire [31:0] _mesh_6_14_io_out_b_0;
	wire _mesh_6_14_io_out_control_0_dataflow;
	wire _mesh_6_14_io_out_control_0_propagate;
	wire [4:0] _mesh_6_14_io_out_control_0_shift;
	wire [2:0] _mesh_6_14_io_out_id_0;
	wire _mesh_6_14_io_out_last_0;
	wire _mesh_6_14_io_out_valid_0;
	wire [31:0] _mesh_6_13_io_out_a_0;
	wire [31:0] _mesh_6_13_io_out_c_0;
	wire [31:0] _mesh_6_13_io_out_b_0;
	wire _mesh_6_13_io_out_control_0_dataflow;
	wire _mesh_6_13_io_out_control_0_propagate;
	wire [4:0] _mesh_6_13_io_out_control_0_shift;
	wire [2:0] _mesh_6_13_io_out_id_0;
	wire _mesh_6_13_io_out_last_0;
	wire _mesh_6_13_io_out_valid_0;
	wire [31:0] _mesh_6_12_io_out_a_0;
	wire [31:0] _mesh_6_12_io_out_c_0;
	wire [31:0] _mesh_6_12_io_out_b_0;
	wire _mesh_6_12_io_out_control_0_dataflow;
	wire _mesh_6_12_io_out_control_0_propagate;
	wire [4:0] _mesh_6_12_io_out_control_0_shift;
	wire [2:0] _mesh_6_12_io_out_id_0;
	wire _mesh_6_12_io_out_last_0;
	wire _mesh_6_12_io_out_valid_0;
	wire [31:0] _mesh_6_11_io_out_a_0;
	wire [31:0] _mesh_6_11_io_out_c_0;
	wire [31:0] _mesh_6_11_io_out_b_0;
	wire _mesh_6_11_io_out_control_0_dataflow;
	wire _mesh_6_11_io_out_control_0_propagate;
	wire [4:0] _mesh_6_11_io_out_control_0_shift;
	wire [2:0] _mesh_6_11_io_out_id_0;
	wire _mesh_6_11_io_out_last_0;
	wire _mesh_6_11_io_out_valid_0;
	wire [31:0] _mesh_6_10_io_out_a_0;
	wire [31:0] _mesh_6_10_io_out_c_0;
	wire [31:0] _mesh_6_10_io_out_b_0;
	wire _mesh_6_10_io_out_control_0_dataflow;
	wire _mesh_6_10_io_out_control_0_propagate;
	wire [4:0] _mesh_6_10_io_out_control_0_shift;
	wire [2:0] _mesh_6_10_io_out_id_0;
	wire _mesh_6_10_io_out_last_0;
	wire _mesh_6_10_io_out_valid_0;
	wire [31:0] _mesh_6_9_io_out_a_0;
	wire [31:0] _mesh_6_9_io_out_c_0;
	wire [31:0] _mesh_6_9_io_out_b_0;
	wire _mesh_6_9_io_out_control_0_dataflow;
	wire _mesh_6_9_io_out_control_0_propagate;
	wire [4:0] _mesh_6_9_io_out_control_0_shift;
	wire [2:0] _mesh_6_9_io_out_id_0;
	wire _mesh_6_9_io_out_last_0;
	wire _mesh_6_9_io_out_valid_0;
	wire [31:0] _mesh_6_8_io_out_a_0;
	wire [31:0] _mesh_6_8_io_out_c_0;
	wire [31:0] _mesh_6_8_io_out_b_0;
	wire _mesh_6_8_io_out_control_0_dataflow;
	wire _mesh_6_8_io_out_control_0_propagate;
	wire [4:0] _mesh_6_8_io_out_control_0_shift;
	wire [2:0] _mesh_6_8_io_out_id_0;
	wire _mesh_6_8_io_out_last_0;
	wire _mesh_6_8_io_out_valid_0;
	wire [31:0] _mesh_6_7_io_out_a_0;
	wire [31:0] _mesh_6_7_io_out_c_0;
	wire [31:0] _mesh_6_7_io_out_b_0;
	wire _mesh_6_7_io_out_control_0_dataflow;
	wire _mesh_6_7_io_out_control_0_propagate;
	wire [4:0] _mesh_6_7_io_out_control_0_shift;
	wire [2:0] _mesh_6_7_io_out_id_0;
	wire _mesh_6_7_io_out_last_0;
	wire _mesh_6_7_io_out_valid_0;
	wire [31:0] _mesh_6_6_io_out_a_0;
	wire [31:0] _mesh_6_6_io_out_c_0;
	wire [31:0] _mesh_6_6_io_out_b_0;
	wire _mesh_6_6_io_out_control_0_dataflow;
	wire _mesh_6_6_io_out_control_0_propagate;
	wire [4:0] _mesh_6_6_io_out_control_0_shift;
	wire [2:0] _mesh_6_6_io_out_id_0;
	wire _mesh_6_6_io_out_last_0;
	wire _mesh_6_6_io_out_valid_0;
	wire [31:0] _mesh_6_5_io_out_a_0;
	wire [31:0] _mesh_6_5_io_out_c_0;
	wire [31:0] _mesh_6_5_io_out_b_0;
	wire _mesh_6_5_io_out_control_0_dataflow;
	wire _mesh_6_5_io_out_control_0_propagate;
	wire [4:0] _mesh_6_5_io_out_control_0_shift;
	wire [2:0] _mesh_6_5_io_out_id_0;
	wire _mesh_6_5_io_out_last_0;
	wire _mesh_6_5_io_out_valid_0;
	wire [31:0] _mesh_6_4_io_out_a_0;
	wire [31:0] _mesh_6_4_io_out_c_0;
	wire [31:0] _mesh_6_4_io_out_b_0;
	wire _mesh_6_4_io_out_control_0_dataflow;
	wire _mesh_6_4_io_out_control_0_propagate;
	wire [4:0] _mesh_6_4_io_out_control_0_shift;
	wire [2:0] _mesh_6_4_io_out_id_0;
	wire _mesh_6_4_io_out_last_0;
	wire _mesh_6_4_io_out_valid_0;
	wire [31:0] _mesh_6_3_io_out_a_0;
	wire [31:0] _mesh_6_3_io_out_c_0;
	wire [31:0] _mesh_6_3_io_out_b_0;
	wire _mesh_6_3_io_out_control_0_dataflow;
	wire _mesh_6_3_io_out_control_0_propagate;
	wire [4:0] _mesh_6_3_io_out_control_0_shift;
	wire [2:0] _mesh_6_3_io_out_id_0;
	wire _mesh_6_3_io_out_last_0;
	wire _mesh_6_3_io_out_valid_0;
	wire [31:0] _mesh_6_2_io_out_a_0;
	wire [31:0] _mesh_6_2_io_out_c_0;
	wire [31:0] _mesh_6_2_io_out_b_0;
	wire _mesh_6_2_io_out_control_0_dataflow;
	wire _mesh_6_2_io_out_control_0_propagate;
	wire [4:0] _mesh_6_2_io_out_control_0_shift;
	wire [2:0] _mesh_6_2_io_out_id_0;
	wire _mesh_6_2_io_out_last_0;
	wire _mesh_6_2_io_out_valid_0;
	wire [31:0] _mesh_6_1_io_out_a_0;
	wire [31:0] _mesh_6_1_io_out_c_0;
	wire [31:0] _mesh_6_1_io_out_b_0;
	wire _mesh_6_1_io_out_control_0_dataflow;
	wire _mesh_6_1_io_out_control_0_propagate;
	wire [4:0] _mesh_6_1_io_out_control_0_shift;
	wire [2:0] _mesh_6_1_io_out_id_0;
	wire _mesh_6_1_io_out_last_0;
	wire _mesh_6_1_io_out_valid_0;
	wire [31:0] _mesh_6_0_io_out_a_0;
	wire [31:0] _mesh_6_0_io_out_c_0;
	wire [31:0] _mesh_6_0_io_out_b_0;
	wire _mesh_6_0_io_out_control_0_dataflow;
	wire _mesh_6_0_io_out_control_0_propagate;
	wire [4:0] _mesh_6_0_io_out_control_0_shift;
	wire [2:0] _mesh_6_0_io_out_id_0;
	wire _mesh_6_0_io_out_last_0;
	wire _mesh_6_0_io_out_valid_0;
	wire [31:0] _mesh_5_15_io_out_a_0;
	wire [31:0] _mesh_5_15_io_out_c_0;
	wire [31:0] _mesh_5_15_io_out_b_0;
	wire _mesh_5_15_io_out_control_0_dataflow;
	wire _mesh_5_15_io_out_control_0_propagate;
	wire [4:0] _mesh_5_15_io_out_control_0_shift;
	wire [2:0] _mesh_5_15_io_out_id_0;
	wire _mesh_5_15_io_out_last_0;
	wire _mesh_5_15_io_out_valid_0;
	wire [31:0] _mesh_5_14_io_out_a_0;
	wire [31:0] _mesh_5_14_io_out_c_0;
	wire [31:0] _mesh_5_14_io_out_b_0;
	wire _mesh_5_14_io_out_control_0_dataflow;
	wire _mesh_5_14_io_out_control_0_propagate;
	wire [4:0] _mesh_5_14_io_out_control_0_shift;
	wire [2:0] _mesh_5_14_io_out_id_0;
	wire _mesh_5_14_io_out_last_0;
	wire _mesh_5_14_io_out_valid_0;
	wire [31:0] _mesh_5_13_io_out_a_0;
	wire [31:0] _mesh_5_13_io_out_c_0;
	wire [31:0] _mesh_5_13_io_out_b_0;
	wire _mesh_5_13_io_out_control_0_dataflow;
	wire _mesh_5_13_io_out_control_0_propagate;
	wire [4:0] _mesh_5_13_io_out_control_0_shift;
	wire [2:0] _mesh_5_13_io_out_id_0;
	wire _mesh_5_13_io_out_last_0;
	wire _mesh_5_13_io_out_valid_0;
	wire [31:0] _mesh_5_12_io_out_a_0;
	wire [31:0] _mesh_5_12_io_out_c_0;
	wire [31:0] _mesh_5_12_io_out_b_0;
	wire _mesh_5_12_io_out_control_0_dataflow;
	wire _mesh_5_12_io_out_control_0_propagate;
	wire [4:0] _mesh_5_12_io_out_control_0_shift;
	wire [2:0] _mesh_5_12_io_out_id_0;
	wire _mesh_5_12_io_out_last_0;
	wire _mesh_5_12_io_out_valid_0;
	wire [31:0] _mesh_5_11_io_out_a_0;
	wire [31:0] _mesh_5_11_io_out_c_0;
	wire [31:0] _mesh_5_11_io_out_b_0;
	wire _mesh_5_11_io_out_control_0_dataflow;
	wire _mesh_5_11_io_out_control_0_propagate;
	wire [4:0] _mesh_5_11_io_out_control_0_shift;
	wire [2:0] _mesh_5_11_io_out_id_0;
	wire _mesh_5_11_io_out_last_0;
	wire _mesh_5_11_io_out_valid_0;
	wire [31:0] _mesh_5_10_io_out_a_0;
	wire [31:0] _mesh_5_10_io_out_c_0;
	wire [31:0] _mesh_5_10_io_out_b_0;
	wire _mesh_5_10_io_out_control_0_dataflow;
	wire _mesh_5_10_io_out_control_0_propagate;
	wire [4:0] _mesh_5_10_io_out_control_0_shift;
	wire [2:0] _mesh_5_10_io_out_id_0;
	wire _mesh_5_10_io_out_last_0;
	wire _mesh_5_10_io_out_valid_0;
	wire [31:0] _mesh_5_9_io_out_a_0;
	wire [31:0] _mesh_5_9_io_out_c_0;
	wire [31:0] _mesh_5_9_io_out_b_0;
	wire _mesh_5_9_io_out_control_0_dataflow;
	wire _mesh_5_9_io_out_control_0_propagate;
	wire [4:0] _mesh_5_9_io_out_control_0_shift;
	wire [2:0] _mesh_5_9_io_out_id_0;
	wire _mesh_5_9_io_out_last_0;
	wire _mesh_5_9_io_out_valid_0;
	wire [31:0] _mesh_5_8_io_out_a_0;
	wire [31:0] _mesh_5_8_io_out_c_0;
	wire [31:0] _mesh_5_8_io_out_b_0;
	wire _mesh_5_8_io_out_control_0_dataflow;
	wire _mesh_5_8_io_out_control_0_propagate;
	wire [4:0] _mesh_5_8_io_out_control_0_shift;
	wire [2:0] _mesh_5_8_io_out_id_0;
	wire _mesh_5_8_io_out_last_0;
	wire _mesh_5_8_io_out_valid_0;
	wire [31:0] _mesh_5_7_io_out_a_0;
	wire [31:0] _mesh_5_7_io_out_c_0;
	wire [31:0] _mesh_5_7_io_out_b_0;
	wire _mesh_5_7_io_out_control_0_dataflow;
	wire _mesh_5_7_io_out_control_0_propagate;
	wire [4:0] _mesh_5_7_io_out_control_0_shift;
	wire [2:0] _mesh_5_7_io_out_id_0;
	wire _mesh_5_7_io_out_last_0;
	wire _mesh_5_7_io_out_valid_0;
	wire [31:0] _mesh_5_6_io_out_a_0;
	wire [31:0] _mesh_5_6_io_out_c_0;
	wire [31:0] _mesh_5_6_io_out_b_0;
	wire _mesh_5_6_io_out_control_0_dataflow;
	wire _mesh_5_6_io_out_control_0_propagate;
	wire [4:0] _mesh_5_6_io_out_control_0_shift;
	wire [2:0] _mesh_5_6_io_out_id_0;
	wire _mesh_5_6_io_out_last_0;
	wire _mesh_5_6_io_out_valid_0;
	wire [31:0] _mesh_5_5_io_out_a_0;
	wire [31:0] _mesh_5_5_io_out_c_0;
	wire [31:0] _mesh_5_5_io_out_b_0;
	wire _mesh_5_5_io_out_control_0_dataflow;
	wire _mesh_5_5_io_out_control_0_propagate;
	wire [4:0] _mesh_5_5_io_out_control_0_shift;
	wire [2:0] _mesh_5_5_io_out_id_0;
	wire _mesh_5_5_io_out_last_0;
	wire _mesh_5_5_io_out_valid_0;
	wire [31:0] _mesh_5_4_io_out_a_0;
	wire [31:0] _mesh_5_4_io_out_c_0;
	wire [31:0] _mesh_5_4_io_out_b_0;
	wire _mesh_5_4_io_out_control_0_dataflow;
	wire _mesh_5_4_io_out_control_0_propagate;
	wire [4:0] _mesh_5_4_io_out_control_0_shift;
	wire [2:0] _mesh_5_4_io_out_id_0;
	wire _mesh_5_4_io_out_last_0;
	wire _mesh_5_4_io_out_valid_0;
	wire [31:0] _mesh_5_3_io_out_a_0;
	wire [31:0] _mesh_5_3_io_out_c_0;
	wire [31:0] _mesh_5_3_io_out_b_0;
	wire _mesh_5_3_io_out_control_0_dataflow;
	wire _mesh_5_3_io_out_control_0_propagate;
	wire [4:0] _mesh_5_3_io_out_control_0_shift;
	wire [2:0] _mesh_5_3_io_out_id_0;
	wire _mesh_5_3_io_out_last_0;
	wire _mesh_5_3_io_out_valid_0;
	wire [31:0] _mesh_5_2_io_out_a_0;
	wire [31:0] _mesh_5_2_io_out_c_0;
	wire [31:0] _mesh_5_2_io_out_b_0;
	wire _mesh_5_2_io_out_control_0_dataflow;
	wire _mesh_5_2_io_out_control_0_propagate;
	wire [4:0] _mesh_5_2_io_out_control_0_shift;
	wire [2:0] _mesh_5_2_io_out_id_0;
	wire _mesh_5_2_io_out_last_0;
	wire _mesh_5_2_io_out_valid_0;
	wire [31:0] _mesh_5_1_io_out_a_0;
	wire [31:0] _mesh_5_1_io_out_c_0;
	wire [31:0] _mesh_5_1_io_out_b_0;
	wire _mesh_5_1_io_out_control_0_dataflow;
	wire _mesh_5_1_io_out_control_0_propagate;
	wire [4:0] _mesh_5_1_io_out_control_0_shift;
	wire [2:0] _mesh_5_1_io_out_id_0;
	wire _mesh_5_1_io_out_last_0;
	wire _mesh_5_1_io_out_valid_0;
	wire [31:0] _mesh_5_0_io_out_a_0;
	wire [31:0] _mesh_5_0_io_out_c_0;
	wire [31:0] _mesh_5_0_io_out_b_0;
	wire _mesh_5_0_io_out_control_0_dataflow;
	wire _mesh_5_0_io_out_control_0_propagate;
	wire [4:0] _mesh_5_0_io_out_control_0_shift;
	wire [2:0] _mesh_5_0_io_out_id_0;
	wire _mesh_5_0_io_out_last_0;
	wire _mesh_5_0_io_out_valid_0;
	wire [31:0] _mesh_4_15_io_out_a_0;
	wire [31:0] _mesh_4_15_io_out_c_0;
	wire [31:0] _mesh_4_15_io_out_b_0;
	wire _mesh_4_15_io_out_control_0_dataflow;
	wire _mesh_4_15_io_out_control_0_propagate;
	wire [4:0] _mesh_4_15_io_out_control_0_shift;
	wire [2:0] _mesh_4_15_io_out_id_0;
	wire _mesh_4_15_io_out_last_0;
	wire _mesh_4_15_io_out_valid_0;
	wire [31:0] _mesh_4_14_io_out_a_0;
	wire [31:0] _mesh_4_14_io_out_c_0;
	wire [31:0] _mesh_4_14_io_out_b_0;
	wire _mesh_4_14_io_out_control_0_dataflow;
	wire _mesh_4_14_io_out_control_0_propagate;
	wire [4:0] _mesh_4_14_io_out_control_0_shift;
	wire [2:0] _mesh_4_14_io_out_id_0;
	wire _mesh_4_14_io_out_last_0;
	wire _mesh_4_14_io_out_valid_0;
	wire [31:0] _mesh_4_13_io_out_a_0;
	wire [31:0] _mesh_4_13_io_out_c_0;
	wire [31:0] _mesh_4_13_io_out_b_0;
	wire _mesh_4_13_io_out_control_0_dataflow;
	wire _mesh_4_13_io_out_control_0_propagate;
	wire [4:0] _mesh_4_13_io_out_control_0_shift;
	wire [2:0] _mesh_4_13_io_out_id_0;
	wire _mesh_4_13_io_out_last_0;
	wire _mesh_4_13_io_out_valid_0;
	wire [31:0] _mesh_4_12_io_out_a_0;
	wire [31:0] _mesh_4_12_io_out_c_0;
	wire [31:0] _mesh_4_12_io_out_b_0;
	wire _mesh_4_12_io_out_control_0_dataflow;
	wire _mesh_4_12_io_out_control_0_propagate;
	wire [4:0] _mesh_4_12_io_out_control_0_shift;
	wire [2:0] _mesh_4_12_io_out_id_0;
	wire _mesh_4_12_io_out_last_0;
	wire _mesh_4_12_io_out_valid_0;
	wire [31:0] _mesh_4_11_io_out_a_0;
	wire [31:0] _mesh_4_11_io_out_c_0;
	wire [31:0] _mesh_4_11_io_out_b_0;
	wire _mesh_4_11_io_out_control_0_dataflow;
	wire _mesh_4_11_io_out_control_0_propagate;
	wire [4:0] _mesh_4_11_io_out_control_0_shift;
	wire [2:0] _mesh_4_11_io_out_id_0;
	wire _mesh_4_11_io_out_last_0;
	wire _mesh_4_11_io_out_valid_0;
	wire [31:0] _mesh_4_10_io_out_a_0;
	wire [31:0] _mesh_4_10_io_out_c_0;
	wire [31:0] _mesh_4_10_io_out_b_0;
	wire _mesh_4_10_io_out_control_0_dataflow;
	wire _mesh_4_10_io_out_control_0_propagate;
	wire [4:0] _mesh_4_10_io_out_control_0_shift;
	wire [2:0] _mesh_4_10_io_out_id_0;
	wire _mesh_4_10_io_out_last_0;
	wire _mesh_4_10_io_out_valid_0;
	wire [31:0] _mesh_4_9_io_out_a_0;
	wire [31:0] _mesh_4_9_io_out_c_0;
	wire [31:0] _mesh_4_9_io_out_b_0;
	wire _mesh_4_9_io_out_control_0_dataflow;
	wire _mesh_4_9_io_out_control_0_propagate;
	wire [4:0] _mesh_4_9_io_out_control_0_shift;
	wire [2:0] _mesh_4_9_io_out_id_0;
	wire _mesh_4_9_io_out_last_0;
	wire _mesh_4_9_io_out_valid_0;
	wire [31:0] _mesh_4_8_io_out_a_0;
	wire [31:0] _mesh_4_8_io_out_c_0;
	wire [31:0] _mesh_4_8_io_out_b_0;
	wire _mesh_4_8_io_out_control_0_dataflow;
	wire _mesh_4_8_io_out_control_0_propagate;
	wire [4:0] _mesh_4_8_io_out_control_0_shift;
	wire [2:0] _mesh_4_8_io_out_id_0;
	wire _mesh_4_8_io_out_last_0;
	wire _mesh_4_8_io_out_valid_0;
	wire [31:0] _mesh_4_7_io_out_a_0;
	wire [31:0] _mesh_4_7_io_out_c_0;
	wire [31:0] _mesh_4_7_io_out_b_0;
	wire _mesh_4_7_io_out_control_0_dataflow;
	wire _mesh_4_7_io_out_control_0_propagate;
	wire [4:0] _mesh_4_7_io_out_control_0_shift;
	wire [2:0] _mesh_4_7_io_out_id_0;
	wire _mesh_4_7_io_out_last_0;
	wire _mesh_4_7_io_out_valid_0;
	wire [31:0] _mesh_4_6_io_out_a_0;
	wire [31:0] _mesh_4_6_io_out_c_0;
	wire [31:0] _mesh_4_6_io_out_b_0;
	wire _mesh_4_6_io_out_control_0_dataflow;
	wire _mesh_4_6_io_out_control_0_propagate;
	wire [4:0] _mesh_4_6_io_out_control_0_shift;
	wire [2:0] _mesh_4_6_io_out_id_0;
	wire _mesh_4_6_io_out_last_0;
	wire _mesh_4_6_io_out_valid_0;
	wire [31:0] _mesh_4_5_io_out_a_0;
	wire [31:0] _mesh_4_5_io_out_c_0;
	wire [31:0] _mesh_4_5_io_out_b_0;
	wire _mesh_4_5_io_out_control_0_dataflow;
	wire _mesh_4_5_io_out_control_0_propagate;
	wire [4:0] _mesh_4_5_io_out_control_0_shift;
	wire [2:0] _mesh_4_5_io_out_id_0;
	wire _mesh_4_5_io_out_last_0;
	wire _mesh_4_5_io_out_valid_0;
	wire [31:0] _mesh_4_4_io_out_a_0;
	wire [31:0] _mesh_4_4_io_out_c_0;
	wire [31:0] _mesh_4_4_io_out_b_0;
	wire _mesh_4_4_io_out_control_0_dataflow;
	wire _mesh_4_4_io_out_control_0_propagate;
	wire [4:0] _mesh_4_4_io_out_control_0_shift;
	wire [2:0] _mesh_4_4_io_out_id_0;
	wire _mesh_4_4_io_out_last_0;
	wire _mesh_4_4_io_out_valid_0;
	wire [31:0] _mesh_4_3_io_out_a_0;
	wire [31:0] _mesh_4_3_io_out_c_0;
	wire [31:0] _mesh_4_3_io_out_b_0;
	wire _mesh_4_3_io_out_control_0_dataflow;
	wire _mesh_4_3_io_out_control_0_propagate;
	wire [4:0] _mesh_4_3_io_out_control_0_shift;
	wire [2:0] _mesh_4_3_io_out_id_0;
	wire _mesh_4_3_io_out_last_0;
	wire _mesh_4_3_io_out_valid_0;
	wire [31:0] _mesh_4_2_io_out_a_0;
	wire [31:0] _mesh_4_2_io_out_c_0;
	wire [31:0] _mesh_4_2_io_out_b_0;
	wire _mesh_4_2_io_out_control_0_dataflow;
	wire _mesh_4_2_io_out_control_0_propagate;
	wire [4:0] _mesh_4_2_io_out_control_0_shift;
	wire [2:0] _mesh_4_2_io_out_id_0;
	wire _mesh_4_2_io_out_last_0;
	wire _mesh_4_2_io_out_valid_0;
	wire [31:0] _mesh_4_1_io_out_a_0;
	wire [31:0] _mesh_4_1_io_out_c_0;
	wire [31:0] _mesh_4_1_io_out_b_0;
	wire _mesh_4_1_io_out_control_0_dataflow;
	wire _mesh_4_1_io_out_control_0_propagate;
	wire [4:0] _mesh_4_1_io_out_control_0_shift;
	wire [2:0] _mesh_4_1_io_out_id_0;
	wire _mesh_4_1_io_out_last_0;
	wire _mesh_4_1_io_out_valid_0;
	wire [31:0] _mesh_4_0_io_out_a_0;
	wire [31:0] _mesh_4_0_io_out_c_0;
	wire [31:0] _mesh_4_0_io_out_b_0;
	wire _mesh_4_0_io_out_control_0_dataflow;
	wire _mesh_4_0_io_out_control_0_propagate;
	wire [4:0] _mesh_4_0_io_out_control_0_shift;
	wire [2:0] _mesh_4_0_io_out_id_0;
	wire _mesh_4_0_io_out_last_0;
	wire _mesh_4_0_io_out_valid_0;
	wire [31:0] _mesh_3_15_io_out_a_0;
	wire [31:0] _mesh_3_15_io_out_c_0;
	wire [31:0] _mesh_3_15_io_out_b_0;
	wire _mesh_3_15_io_out_control_0_dataflow;
	wire _mesh_3_15_io_out_control_0_propagate;
	wire [4:0] _mesh_3_15_io_out_control_0_shift;
	wire [2:0] _mesh_3_15_io_out_id_0;
	wire _mesh_3_15_io_out_last_0;
	wire _mesh_3_15_io_out_valid_0;
	wire [31:0] _mesh_3_14_io_out_a_0;
	wire [31:0] _mesh_3_14_io_out_c_0;
	wire [31:0] _mesh_3_14_io_out_b_0;
	wire _mesh_3_14_io_out_control_0_dataflow;
	wire _mesh_3_14_io_out_control_0_propagate;
	wire [4:0] _mesh_3_14_io_out_control_0_shift;
	wire [2:0] _mesh_3_14_io_out_id_0;
	wire _mesh_3_14_io_out_last_0;
	wire _mesh_3_14_io_out_valid_0;
	wire [31:0] _mesh_3_13_io_out_a_0;
	wire [31:0] _mesh_3_13_io_out_c_0;
	wire [31:0] _mesh_3_13_io_out_b_0;
	wire _mesh_3_13_io_out_control_0_dataflow;
	wire _mesh_3_13_io_out_control_0_propagate;
	wire [4:0] _mesh_3_13_io_out_control_0_shift;
	wire [2:0] _mesh_3_13_io_out_id_0;
	wire _mesh_3_13_io_out_last_0;
	wire _mesh_3_13_io_out_valid_0;
	wire [31:0] _mesh_3_12_io_out_a_0;
	wire [31:0] _mesh_3_12_io_out_c_0;
	wire [31:0] _mesh_3_12_io_out_b_0;
	wire _mesh_3_12_io_out_control_0_dataflow;
	wire _mesh_3_12_io_out_control_0_propagate;
	wire [4:0] _mesh_3_12_io_out_control_0_shift;
	wire [2:0] _mesh_3_12_io_out_id_0;
	wire _mesh_3_12_io_out_last_0;
	wire _mesh_3_12_io_out_valid_0;
	wire [31:0] _mesh_3_11_io_out_a_0;
	wire [31:0] _mesh_3_11_io_out_c_0;
	wire [31:0] _mesh_3_11_io_out_b_0;
	wire _mesh_3_11_io_out_control_0_dataflow;
	wire _mesh_3_11_io_out_control_0_propagate;
	wire [4:0] _mesh_3_11_io_out_control_0_shift;
	wire [2:0] _mesh_3_11_io_out_id_0;
	wire _mesh_3_11_io_out_last_0;
	wire _mesh_3_11_io_out_valid_0;
	wire [31:0] _mesh_3_10_io_out_a_0;
	wire [31:0] _mesh_3_10_io_out_c_0;
	wire [31:0] _mesh_3_10_io_out_b_0;
	wire _mesh_3_10_io_out_control_0_dataflow;
	wire _mesh_3_10_io_out_control_0_propagate;
	wire [4:0] _mesh_3_10_io_out_control_0_shift;
	wire [2:0] _mesh_3_10_io_out_id_0;
	wire _mesh_3_10_io_out_last_0;
	wire _mesh_3_10_io_out_valid_0;
	wire [31:0] _mesh_3_9_io_out_a_0;
	wire [31:0] _mesh_3_9_io_out_c_0;
	wire [31:0] _mesh_3_9_io_out_b_0;
	wire _mesh_3_9_io_out_control_0_dataflow;
	wire _mesh_3_9_io_out_control_0_propagate;
	wire [4:0] _mesh_3_9_io_out_control_0_shift;
	wire [2:0] _mesh_3_9_io_out_id_0;
	wire _mesh_3_9_io_out_last_0;
	wire _mesh_3_9_io_out_valid_0;
	wire [31:0] _mesh_3_8_io_out_a_0;
	wire [31:0] _mesh_3_8_io_out_c_0;
	wire [31:0] _mesh_3_8_io_out_b_0;
	wire _mesh_3_8_io_out_control_0_dataflow;
	wire _mesh_3_8_io_out_control_0_propagate;
	wire [4:0] _mesh_3_8_io_out_control_0_shift;
	wire [2:0] _mesh_3_8_io_out_id_0;
	wire _mesh_3_8_io_out_last_0;
	wire _mesh_3_8_io_out_valid_0;
	wire [31:0] _mesh_3_7_io_out_a_0;
	wire [31:0] _mesh_3_7_io_out_c_0;
	wire [31:0] _mesh_3_7_io_out_b_0;
	wire _mesh_3_7_io_out_control_0_dataflow;
	wire _mesh_3_7_io_out_control_0_propagate;
	wire [4:0] _mesh_3_7_io_out_control_0_shift;
	wire [2:0] _mesh_3_7_io_out_id_0;
	wire _mesh_3_7_io_out_last_0;
	wire _mesh_3_7_io_out_valid_0;
	wire [31:0] _mesh_3_6_io_out_a_0;
	wire [31:0] _mesh_3_6_io_out_c_0;
	wire [31:0] _mesh_3_6_io_out_b_0;
	wire _mesh_3_6_io_out_control_0_dataflow;
	wire _mesh_3_6_io_out_control_0_propagate;
	wire [4:0] _mesh_3_6_io_out_control_0_shift;
	wire [2:0] _mesh_3_6_io_out_id_0;
	wire _mesh_3_6_io_out_last_0;
	wire _mesh_3_6_io_out_valid_0;
	wire [31:0] _mesh_3_5_io_out_a_0;
	wire [31:0] _mesh_3_5_io_out_c_0;
	wire [31:0] _mesh_3_5_io_out_b_0;
	wire _mesh_3_5_io_out_control_0_dataflow;
	wire _mesh_3_5_io_out_control_0_propagate;
	wire [4:0] _mesh_3_5_io_out_control_0_shift;
	wire [2:0] _mesh_3_5_io_out_id_0;
	wire _mesh_3_5_io_out_last_0;
	wire _mesh_3_5_io_out_valid_0;
	wire [31:0] _mesh_3_4_io_out_a_0;
	wire [31:0] _mesh_3_4_io_out_c_0;
	wire [31:0] _mesh_3_4_io_out_b_0;
	wire _mesh_3_4_io_out_control_0_dataflow;
	wire _mesh_3_4_io_out_control_0_propagate;
	wire [4:0] _mesh_3_4_io_out_control_0_shift;
	wire [2:0] _mesh_3_4_io_out_id_0;
	wire _mesh_3_4_io_out_last_0;
	wire _mesh_3_4_io_out_valid_0;
	wire [31:0] _mesh_3_3_io_out_a_0;
	wire [31:0] _mesh_3_3_io_out_c_0;
	wire [31:0] _mesh_3_3_io_out_b_0;
	wire _mesh_3_3_io_out_control_0_dataflow;
	wire _mesh_3_3_io_out_control_0_propagate;
	wire [4:0] _mesh_3_3_io_out_control_0_shift;
	wire [2:0] _mesh_3_3_io_out_id_0;
	wire _mesh_3_3_io_out_last_0;
	wire _mesh_3_3_io_out_valid_0;
	wire [31:0] _mesh_3_2_io_out_a_0;
	wire [31:0] _mesh_3_2_io_out_c_0;
	wire [31:0] _mesh_3_2_io_out_b_0;
	wire _mesh_3_2_io_out_control_0_dataflow;
	wire _mesh_3_2_io_out_control_0_propagate;
	wire [4:0] _mesh_3_2_io_out_control_0_shift;
	wire [2:0] _mesh_3_2_io_out_id_0;
	wire _mesh_3_2_io_out_last_0;
	wire _mesh_3_2_io_out_valid_0;
	wire [31:0] _mesh_3_1_io_out_a_0;
	wire [31:0] _mesh_3_1_io_out_c_0;
	wire [31:0] _mesh_3_1_io_out_b_0;
	wire _mesh_3_1_io_out_control_0_dataflow;
	wire _mesh_3_1_io_out_control_0_propagate;
	wire [4:0] _mesh_3_1_io_out_control_0_shift;
	wire [2:0] _mesh_3_1_io_out_id_0;
	wire _mesh_3_1_io_out_last_0;
	wire _mesh_3_1_io_out_valid_0;
	wire [31:0] _mesh_3_0_io_out_a_0;
	wire [31:0] _mesh_3_0_io_out_c_0;
	wire [31:0] _mesh_3_0_io_out_b_0;
	wire _mesh_3_0_io_out_control_0_dataflow;
	wire _mesh_3_0_io_out_control_0_propagate;
	wire [4:0] _mesh_3_0_io_out_control_0_shift;
	wire [2:0] _mesh_3_0_io_out_id_0;
	wire _mesh_3_0_io_out_last_0;
	wire _mesh_3_0_io_out_valid_0;
	wire [31:0] _mesh_2_15_io_out_a_0;
	wire [31:0] _mesh_2_15_io_out_c_0;
	wire [31:0] _mesh_2_15_io_out_b_0;
	wire _mesh_2_15_io_out_control_0_dataflow;
	wire _mesh_2_15_io_out_control_0_propagate;
	wire [4:0] _mesh_2_15_io_out_control_0_shift;
	wire [2:0] _mesh_2_15_io_out_id_0;
	wire _mesh_2_15_io_out_last_0;
	wire _mesh_2_15_io_out_valid_0;
	wire [31:0] _mesh_2_14_io_out_a_0;
	wire [31:0] _mesh_2_14_io_out_c_0;
	wire [31:0] _mesh_2_14_io_out_b_0;
	wire _mesh_2_14_io_out_control_0_dataflow;
	wire _mesh_2_14_io_out_control_0_propagate;
	wire [4:0] _mesh_2_14_io_out_control_0_shift;
	wire [2:0] _mesh_2_14_io_out_id_0;
	wire _mesh_2_14_io_out_last_0;
	wire _mesh_2_14_io_out_valid_0;
	wire [31:0] _mesh_2_13_io_out_a_0;
	wire [31:0] _mesh_2_13_io_out_c_0;
	wire [31:0] _mesh_2_13_io_out_b_0;
	wire _mesh_2_13_io_out_control_0_dataflow;
	wire _mesh_2_13_io_out_control_0_propagate;
	wire [4:0] _mesh_2_13_io_out_control_0_shift;
	wire [2:0] _mesh_2_13_io_out_id_0;
	wire _mesh_2_13_io_out_last_0;
	wire _mesh_2_13_io_out_valid_0;
	wire [31:0] _mesh_2_12_io_out_a_0;
	wire [31:0] _mesh_2_12_io_out_c_0;
	wire [31:0] _mesh_2_12_io_out_b_0;
	wire _mesh_2_12_io_out_control_0_dataflow;
	wire _mesh_2_12_io_out_control_0_propagate;
	wire [4:0] _mesh_2_12_io_out_control_0_shift;
	wire [2:0] _mesh_2_12_io_out_id_0;
	wire _mesh_2_12_io_out_last_0;
	wire _mesh_2_12_io_out_valid_0;
	wire [31:0] _mesh_2_11_io_out_a_0;
	wire [31:0] _mesh_2_11_io_out_c_0;
	wire [31:0] _mesh_2_11_io_out_b_0;
	wire _mesh_2_11_io_out_control_0_dataflow;
	wire _mesh_2_11_io_out_control_0_propagate;
	wire [4:0] _mesh_2_11_io_out_control_0_shift;
	wire [2:0] _mesh_2_11_io_out_id_0;
	wire _mesh_2_11_io_out_last_0;
	wire _mesh_2_11_io_out_valid_0;
	wire [31:0] _mesh_2_10_io_out_a_0;
	wire [31:0] _mesh_2_10_io_out_c_0;
	wire [31:0] _mesh_2_10_io_out_b_0;
	wire _mesh_2_10_io_out_control_0_dataflow;
	wire _mesh_2_10_io_out_control_0_propagate;
	wire [4:0] _mesh_2_10_io_out_control_0_shift;
	wire [2:0] _mesh_2_10_io_out_id_0;
	wire _mesh_2_10_io_out_last_0;
	wire _mesh_2_10_io_out_valid_0;
	wire [31:0] _mesh_2_9_io_out_a_0;
	wire [31:0] _mesh_2_9_io_out_c_0;
	wire [31:0] _mesh_2_9_io_out_b_0;
	wire _mesh_2_9_io_out_control_0_dataflow;
	wire _mesh_2_9_io_out_control_0_propagate;
	wire [4:0] _mesh_2_9_io_out_control_0_shift;
	wire [2:0] _mesh_2_9_io_out_id_0;
	wire _mesh_2_9_io_out_last_0;
	wire _mesh_2_9_io_out_valid_0;
	wire [31:0] _mesh_2_8_io_out_a_0;
	wire [31:0] _mesh_2_8_io_out_c_0;
	wire [31:0] _mesh_2_8_io_out_b_0;
	wire _mesh_2_8_io_out_control_0_dataflow;
	wire _mesh_2_8_io_out_control_0_propagate;
	wire [4:0] _mesh_2_8_io_out_control_0_shift;
	wire [2:0] _mesh_2_8_io_out_id_0;
	wire _mesh_2_8_io_out_last_0;
	wire _mesh_2_8_io_out_valid_0;
	wire [31:0] _mesh_2_7_io_out_a_0;
	wire [31:0] _mesh_2_7_io_out_c_0;
	wire [31:0] _mesh_2_7_io_out_b_0;
	wire _mesh_2_7_io_out_control_0_dataflow;
	wire _mesh_2_7_io_out_control_0_propagate;
	wire [4:0] _mesh_2_7_io_out_control_0_shift;
	wire [2:0] _mesh_2_7_io_out_id_0;
	wire _mesh_2_7_io_out_last_0;
	wire _mesh_2_7_io_out_valid_0;
	wire [31:0] _mesh_2_6_io_out_a_0;
	wire [31:0] _mesh_2_6_io_out_c_0;
	wire [31:0] _mesh_2_6_io_out_b_0;
	wire _mesh_2_6_io_out_control_0_dataflow;
	wire _mesh_2_6_io_out_control_0_propagate;
	wire [4:0] _mesh_2_6_io_out_control_0_shift;
	wire [2:0] _mesh_2_6_io_out_id_0;
	wire _mesh_2_6_io_out_last_0;
	wire _mesh_2_6_io_out_valid_0;
	wire [31:0] _mesh_2_5_io_out_a_0;
	wire [31:0] _mesh_2_5_io_out_c_0;
	wire [31:0] _mesh_2_5_io_out_b_0;
	wire _mesh_2_5_io_out_control_0_dataflow;
	wire _mesh_2_5_io_out_control_0_propagate;
	wire [4:0] _mesh_2_5_io_out_control_0_shift;
	wire [2:0] _mesh_2_5_io_out_id_0;
	wire _mesh_2_5_io_out_last_0;
	wire _mesh_2_5_io_out_valid_0;
	wire [31:0] _mesh_2_4_io_out_a_0;
	wire [31:0] _mesh_2_4_io_out_c_0;
	wire [31:0] _mesh_2_4_io_out_b_0;
	wire _mesh_2_4_io_out_control_0_dataflow;
	wire _mesh_2_4_io_out_control_0_propagate;
	wire [4:0] _mesh_2_4_io_out_control_0_shift;
	wire [2:0] _mesh_2_4_io_out_id_0;
	wire _mesh_2_4_io_out_last_0;
	wire _mesh_2_4_io_out_valid_0;
	wire [31:0] _mesh_2_3_io_out_a_0;
	wire [31:0] _mesh_2_3_io_out_c_0;
	wire [31:0] _mesh_2_3_io_out_b_0;
	wire _mesh_2_3_io_out_control_0_dataflow;
	wire _mesh_2_3_io_out_control_0_propagate;
	wire [4:0] _mesh_2_3_io_out_control_0_shift;
	wire [2:0] _mesh_2_3_io_out_id_0;
	wire _mesh_2_3_io_out_last_0;
	wire _mesh_2_3_io_out_valid_0;
	wire [31:0] _mesh_2_2_io_out_a_0;
	wire [31:0] _mesh_2_2_io_out_c_0;
	wire [31:0] _mesh_2_2_io_out_b_0;
	wire _mesh_2_2_io_out_control_0_dataflow;
	wire _mesh_2_2_io_out_control_0_propagate;
	wire [4:0] _mesh_2_2_io_out_control_0_shift;
	wire [2:0] _mesh_2_2_io_out_id_0;
	wire _mesh_2_2_io_out_last_0;
	wire _mesh_2_2_io_out_valid_0;
	wire [31:0] _mesh_2_1_io_out_a_0;
	wire [31:0] _mesh_2_1_io_out_c_0;
	wire [31:0] _mesh_2_1_io_out_b_0;
	wire _mesh_2_1_io_out_control_0_dataflow;
	wire _mesh_2_1_io_out_control_0_propagate;
	wire [4:0] _mesh_2_1_io_out_control_0_shift;
	wire [2:0] _mesh_2_1_io_out_id_0;
	wire _mesh_2_1_io_out_last_0;
	wire _mesh_2_1_io_out_valid_0;
	wire [31:0] _mesh_2_0_io_out_a_0;
	wire [31:0] _mesh_2_0_io_out_c_0;
	wire [31:0] _mesh_2_0_io_out_b_0;
	wire _mesh_2_0_io_out_control_0_dataflow;
	wire _mesh_2_0_io_out_control_0_propagate;
	wire [4:0] _mesh_2_0_io_out_control_0_shift;
	wire [2:0] _mesh_2_0_io_out_id_0;
	wire _mesh_2_0_io_out_last_0;
	wire _mesh_2_0_io_out_valid_0;
	wire [31:0] _mesh_1_15_io_out_a_0;
	wire [31:0] _mesh_1_15_io_out_c_0;
	wire [31:0] _mesh_1_15_io_out_b_0;
	wire _mesh_1_15_io_out_control_0_dataflow;
	wire _mesh_1_15_io_out_control_0_propagate;
	wire [4:0] _mesh_1_15_io_out_control_0_shift;
	wire [2:0] _mesh_1_15_io_out_id_0;
	wire _mesh_1_15_io_out_last_0;
	wire _mesh_1_15_io_out_valid_0;
	wire [31:0] _mesh_1_14_io_out_a_0;
	wire [31:0] _mesh_1_14_io_out_c_0;
	wire [31:0] _mesh_1_14_io_out_b_0;
	wire _mesh_1_14_io_out_control_0_dataflow;
	wire _mesh_1_14_io_out_control_0_propagate;
	wire [4:0] _mesh_1_14_io_out_control_0_shift;
	wire [2:0] _mesh_1_14_io_out_id_0;
	wire _mesh_1_14_io_out_last_0;
	wire _mesh_1_14_io_out_valid_0;
	wire [31:0] _mesh_1_13_io_out_a_0;
	wire [31:0] _mesh_1_13_io_out_c_0;
	wire [31:0] _mesh_1_13_io_out_b_0;
	wire _mesh_1_13_io_out_control_0_dataflow;
	wire _mesh_1_13_io_out_control_0_propagate;
	wire [4:0] _mesh_1_13_io_out_control_0_shift;
	wire [2:0] _mesh_1_13_io_out_id_0;
	wire _mesh_1_13_io_out_last_0;
	wire _mesh_1_13_io_out_valid_0;
	wire [31:0] _mesh_1_12_io_out_a_0;
	wire [31:0] _mesh_1_12_io_out_c_0;
	wire [31:0] _mesh_1_12_io_out_b_0;
	wire _mesh_1_12_io_out_control_0_dataflow;
	wire _mesh_1_12_io_out_control_0_propagate;
	wire [4:0] _mesh_1_12_io_out_control_0_shift;
	wire [2:0] _mesh_1_12_io_out_id_0;
	wire _mesh_1_12_io_out_last_0;
	wire _mesh_1_12_io_out_valid_0;
	wire [31:0] _mesh_1_11_io_out_a_0;
	wire [31:0] _mesh_1_11_io_out_c_0;
	wire [31:0] _mesh_1_11_io_out_b_0;
	wire _mesh_1_11_io_out_control_0_dataflow;
	wire _mesh_1_11_io_out_control_0_propagate;
	wire [4:0] _mesh_1_11_io_out_control_0_shift;
	wire [2:0] _mesh_1_11_io_out_id_0;
	wire _mesh_1_11_io_out_last_0;
	wire _mesh_1_11_io_out_valid_0;
	wire [31:0] _mesh_1_10_io_out_a_0;
	wire [31:0] _mesh_1_10_io_out_c_0;
	wire [31:0] _mesh_1_10_io_out_b_0;
	wire _mesh_1_10_io_out_control_0_dataflow;
	wire _mesh_1_10_io_out_control_0_propagate;
	wire [4:0] _mesh_1_10_io_out_control_0_shift;
	wire [2:0] _mesh_1_10_io_out_id_0;
	wire _mesh_1_10_io_out_last_0;
	wire _mesh_1_10_io_out_valid_0;
	wire [31:0] _mesh_1_9_io_out_a_0;
	wire [31:0] _mesh_1_9_io_out_c_0;
	wire [31:0] _mesh_1_9_io_out_b_0;
	wire _mesh_1_9_io_out_control_0_dataflow;
	wire _mesh_1_9_io_out_control_0_propagate;
	wire [4:0] _mesh_1_9_io_out_control_0_shift;
	wire [2:0] _mesh_1_9_io_out_id_0;
	wire _mesh_1_9_io_out_last_0;
	wire _mesh_1_9_io_out_valid_0;
	wire [31:0] _mesh_1_8_io_out_a_0;
	wire [31:0] _mesh_1_8_io_out_c_0;
	wire [31:0] _mesh_1_8_io_out_b_0;
	wire _mesh_1_8_io_out_control_0_dataflow;
	wire _mesh_1_8_io_out_control_0_propagate;
	wire [4:0] _mesh_1_8_io_out_control_0_shift;
	wire [2:0] _mesh_1_8_io_out_id_0;
	wire _mesh_1_8_io_out_last_0;
	wire _mesh_1_8_io_out_valid_0;
	wire [31:0] _mesh_1_7_io_out_a_0;
	wire [31:0] _mesh_1_7_io_out_c_0;
	wire [31:0] _mesh_1_7_io_out_b_0;
	wire _mesh_1_7_io_out_control_0_dataflow;
	wire _mesh_1_7_io_out_control_0_propagate;
	wire [4:0] _mesh_1_7_io_out_control_0_shift;
	wire [2:0] _mesh_1_7_io_out_id_0;
	wire _mesh_1_7_io_out_last_0;
	wire _mesh_1_7_io_out_valid_0;
	wire [31:0] _mesh_1_6_io_out_a_0;
	wire [31:0] _mesh_1_6_io_out_c_0;
	wire [31:0] _mesh_1_6_io_out_b_0;
	wire _mesh_1_6_io_out_control_0_dataflow;
	wire _mesh_1_6_io_out_control_0_propagate;
	wire [4:0] _mesh_1_6_io_out_control_0_shift;
	wire [2:0] _mesh_1_6_io_out_id_0;
	wire _mesh_1_6_io_out_last_0;
	wire _mesh_1_6_io_out_valid_0;
	wire [31:0] _mesh_1_5_io_out_a_0;
	wire [31:0] _mesh_1_5_io_out_c_0;
	wire [31:0] _mesh_1_5_io_out_b_0;
	wire _mesh_1_5_io_out_control_0_dataflow;
	wire _mesh_1_5_io_out_control_0_propagate;
	wire [4:0] _mesh_1_5_io_out_control_0_shift;
	wire [2:0] _mesh_1_5_io_out_id_0;
	wire _mesh_1_5_io_out_last_0;
	wire _mesh_1_5_io_out_valid_0;
	wire [31:0] _mesh_1_4_io_out_a_0;
	wire [31:0] _mesh_1_4_io_out_c_0;
	wire [31:0] _mesh_1_4_io_out_b_0;
	wire _mesh_1_4_io_out_control_0_dataflow;
	wire _mesh_1_4_io_out_control_0_propagate;
	wire [4:0] _mesh_1_4_io_out_control_0_shift;
	wire [2:0] _mesh_1_4_io_out_id_0;
	wire _mesh_1_4_io_out_last_0;
	wire _mesh_1_4_io_out_valid_0;
	wire [31:0] _mesh_1_3_io_out_a_0;
	wire [31:0] _mesh_1_3_io_out_c_0;
	wire [31:0] _mesh_1_3_io_out_b_0;
	wire _mesh_1_3_io_out_control_0_dataflow;
	wire _mesh_1_3_io_out_control_0_propagate;
	wire [4:0] _mesh_1_3_io_out_control_0_shift;
	wire [2:0] _mesh_1_3_io_out_id_0;
	wire _mesh_1_3_io_out_last_0;
	wire _mesh_1_3_io_out_valid_0;
	wire [31:0] _mesh_1_2_io_out_a_0;
	wire [31:0] _mesh_1_2_io_out_c_0;
	wire [31:0] _mesh_1_2_io_out_b_0;
	wire _mesh_1_2_io_out_control_0_dataflow;
	wire _mesh_1_2_io_out_control_0_propagate;
	wire [4:0] _mesh_1_2_io_out_control_0_shift;
	wire [2:0] _mesh_1_2_io_out_id_0;
	wire _mesh_1_2_io_out_last_0;
	wire _mesh_1_2_io_out_valid_0;
	wire [31:0] _mesh_1_1_io_out_a_0;
	wire [31:0] _mesh_1_1_io_out_c_0;
	wire [31:0] _mesh_1_1_io_out_b_0;
	wire _mesh_1_1_io_out_control_0_dataflow;
	wire _mesh_1_1_io_out_control_0_propagate;
	wire [4:0] _mesh_1_1_io_out_control_0_shift;
	wire [2:0] _mesh_1_1_io_out_id_0;
	wire _mesh_1_1_io_out_last_0;
	wire _mesh_1_1_io_out_valid_0;
	wire [31:0] _mesh_1_0_io_out_a_0;
	wire [31:0] _mesh_1_0_io_out_c_0;
	wire [31:0] _mesh_1_0_io_out_b_0;
	wire _mesh_1_0_io_out_control_0_dataflow;
	wire _mesh_1_0_io_out_control_0_propagate;
	wire [4:0] _mesh_1_0_io_out_control_0_shift;
	wire [2:0] _mesh_1_0_io_out_id_0;
	wire _mesh_1_0_io_out_last_0;
	wire _mesh_1_0_io_out_valid_0;
	wire [31:0] _mesh_0_15_io_out_a_0;
	wire [31:0] _mesh_0_15_io_out_c_0;
	wire [31:0] _mesh_0_15_io_out_b_0;
	wire _mesh_0_15_io_out_control_0_dataflow;
	wire _mesh_0_15_io_out_control_0_propagate;
	wire [4:0] _mesh_0_15_io_out_control_0_shift;
	wire [2:0] _mesh_0_15_io_out_id_0;
	wire _mesh_0_15_io_out_last_0;
	wire _mesh_0_15_io_out_valid_0;
	wire [31:0] _mesh_0_14_io_out_a_0;
	wire [31:0] _mesh_0_14_io_out_c_0;
	wire [31:0] _mesh_0_14_io_out_b_0;
	wire _mesh_0_14_io_out_control_0_dataflow;
	wire _mesh_0_14_io_out_control_0_propagate;
	wire [4:0] _mesh_0_14_io_out_control_0_shift;
	wire [2:0] _mesh_0_14_io_out_id_0;
	wire _mesh_0_14_io_out_last_0;
	wire _mesh_0_14_io_out_valid_0;
	wire [31:0] _mesh_0_13_io_out_a_0;
	wire [31:0] _mesh_0_13_io_out_c_0;
	wire [31:0] _mesh_0_13_io_out_b_0;
	wire _mesh_0_13_io_out_control_0_dataflow;
	wire _mesh_0_13_io_out_control_0_propagate;
	wire [4:0] _mesh_0_13_io_out_control_0_shift;
	wire [2:0] _mesh_0_13_io_out_id_0;
	wire _mesh_0_13_io_out_last_0;
	wire _mesh_0_13_io_out_valid_0;
	wire [31:0] _mesh_0_12_io_out_a_0;
	wire [31:0] _mesh_0_12_io_out_c_0;
	wire [31:0] _mesh_0_12_io_out_b_0;
	wire _mesh_0_12_io_out_control_0_dataflow;
	wire _mesh_0_12_io_out_control_0_propagate;
	wire [4:0] _mesh_0_12_io_out_control_0_shift;
	wire [2:0] _mesh_0_12_io_out_id_0;
	wire _mesh_0_12_io_out_last_0;
	wire _mesh_0_12_io_out_valid_0;
	wire [31:0] _mesh_0_11_io_out_a_0;
	wire [31:0] _mesh_0_11_io_out_c_0;
	wire [31:0] _mesh_0_11_io_out_b_0;
	wire _mesh_0_11_io_out_control_0_dataflow;
	wire _mesh_0_11_io_out_control_0_propagate;
	wire [4:0] _mesh_0_11_io_out_control_0_shift;
	wire [2:0] _mesh_0_11_io_out_id_0;
	wire _mesh_0_11_io_out_last_0;
	wire _mesh_0_11_io_out_valid_0;
	wire [31:0] _mesh_0_10_io_out_a_0;
	wire [31:0] _mesh_0_10_io_out_c_0;
	wire [31:0] _mesh_0_10_io_out_b_0;
	wire _mesh_0_10_io_out_control_0_dataflow;
	wire _mesh_0_10_io_out_control_0_propagate;
	wire [4:0] _mesh_0_10_io_out_control_0_shift;
	wire [2:0] _mesh_0_10_io_out_id_0;
	wire _mesh_0_10_io_out_last_0;
	wire _mesh_0_10_io_out_valid_0;
	wire [31:0] _mesh_0_9_io_out_a_0;
	wire [31:0] _mesh_0_9_io_out_c_0;
	wire [31:0] _mesh_0_9_io_out_b_0;
	wire _mesh_0_9_io_out_control_0_dataflow;
	wire _mesh_0_9_io_out_control_0_propagate;
	wire [4:0] _mesh_0_9_io_out_control_0_shift;
	wire [2:0] _mesh_0_9_io_out_id_0;
	wire _mesh_0_9_io_out_last_0;
	wire _mesh_0_9_io_out_valid_0;
	wire [31:0] _mesh_0_8_io_out_a_0;
	wire [31:0] _mesh_0_8_io_out_c_0;
	wire [31:0] _mesh_0_8_io_out_b_0;
	wire _mesh_0_8_io_out_control_0_dataflow;
	wire _mesh_0_8_io_out_control_0_propagate;
	wire [4:0] _mesh_0_8_io_out_control_0_shift;
	wire [2:0] _mesh_0_8_io_out_id_0;
	wire _mesh_0_8_io_out_last_0;
	wire _mesh_0_8_io_out_valid_0;
	wire [31:0] _mesh_0_7_io_out_a_0;
	wire [31:0] _mesh_0_7_io_out_c_0;
	wire [31:0] _mesh_0_7_io_out_b_0;
	wire _mesh_0_7_io_out_control_0_dataflow;
	wire _mesh_0_7_io_out_control_0_propagate;
	wire [4:0] _mesh_0_7_io_out_control_0_shift;
	wire [2:0] _mesh_0_7_io_out_id_0;
	wire _mesh_0_7_io_out_last_0;
	wire _mesh_0_7_io_out_valid_0;
	wire [31:0] _mesh_0_6_io_out_a_0;
	wire [31:0] _mesh_0_6_io_out_c_0;
	wire [31:0] _mesh_0_6_io_out_b_0;
	wire _mesh_0_6_io_out_control_0_dataflow;
	wire _mesh_0_6_io_out_control_0_propagate;
	wire [4:0] _mesh_0_6_io_out_control_0_shift;
	wire [2:0] _mesh_0_6_io_out_id_0;
	wire _mesh_0_6_io_out_last_0;
	wire _mesh_0_6_io_out_valid_0;
	wire [31:0] _mesh_0_5_io_out_a_0;
	wire [31:0] _mesh_0_5_io_out_c_0;
	wire [31:0] _mesh_0_5_io_out_b_0;
	wire _mesh_0_5_io_out_control_0_dataflow;
	wire _mesh_0_5_io_out_control_0_propagate;
	wire [4:0] _mesh_0_5_io_out_control_0_shift;
	wire [2:0] _mesh_0_5_io_out_id_0;
	wire _mesh_0_5_io_out_last_0;
	wire _mesh_0_5_io_out_valid_0;
	wire [31:0] _mesh_0_4_io_out_a_0;
	wire [31:0] _mesh_0_4_io_out_c_0;
	wire [31:0] _mesh_0_4_io_out_b_0;
	wire _mesh_0_4_io_out_control_0_dataflow;
	wire _mesh_0_4_io_out_control_0_propagate;
	wire [4:0] _mesh_0_4_io_out_control_0_shift;
	wire [2:0] _mesh_0_4_io_out_id_0;
	wire _mesh_0_4_io_out_last_0;
	wire _mesh_0_4_io_out_valid_0;
	wire [31:0] _mesh_0_3_io_out_a_0;
	wire [31:0] _mesh_0_3_io_out_c_0;
	wire [31:0] _mesh_0_3_io_out_b_0;
	wire _mesh_0_3_io_out_control_0_dataflow;
	wire _mesh_0_3_io_out_control_0_propagate;
	wire [4:0] _mesh_0_3_io_out_control_0_shift;
	wire [2:0] _mesh_0_3_io_out_id_0;
	wire _mesh_0_3_io_out_last_0;
	wire _mesh_0_3_io_out_valid_0;
	wire [31:0] _mesh_0_2_io_out_a_0;
	wire [31:0] _mesh_0_2_io_out_c_0;
	wire [31:0] _mesh_0_2_io_out_b_0;
	wire _mesh_0_2_io_out_control_0_dataflow;
	wire _mesh_0_2_io_out_control_0_propagate;
	wire [4:0] _mesh_0_2_io_out_control_0_shift;
	wire [2:0] _mesh_0_2_io_out_id_0;
	wire _mesh_0_2_io_out_last_0;
	wire _mesh_0_2_io_out_valid_0;
	wire [31:0] _mesh_0_1_io_out_a_0;
	wire [31:0] _mesh_0_1_io_out_c_0;
	wire [31:0] _mesh_0_1_io_out_b_0;
	wire _mesh_0_1_io_out_control_0_dataflow;
	wire _mesh_0_1_io_out_control_0_propagate;
	wire [4:0] _mesh_0_1_io_out_control_0_shift;
	wire [2:0] _mesh_0_1_io_out_id_0;
	wire _mesh_0_1_io_out_last_0;
	wire _mesh_0_1_io_out_valid_0;
	wire [31:0] _mesh_0_0_io_out_a_0;
	wire [31:0] _mesh_0_0_io_out_c_0;
	wire [31:0] _mesh_0_0_io_out_b_0;
	wire _mesh_0_0_io_out_control_0_dataflow;
	wire _mesh_0_0_io_out_control_0_propagate;
	wire [4:0] _mesh_0_0_io_out_control_0_shift;
	wire [2:0] _mesh_0_0_io_out_id_0;
	wire _mesh_0_0_io_out_last_0;
	wire _mesh_0_0_io_out_valid_0;
	reg [31:0] r_0;
	reg [31:0] r_1_0;
	reg [31:0] r_2_0;
	reg [31:0] r_3_0;
	reg [31:0] r_4_0;
	reg [31:0] r_5_0;
	reg [31:0] r_6_0;
	reg [31:0] r_7_0;
	reg [31:0] r_8_0;
	reg [31:0] r_9_0;
	reg [31:0] r_10_0;
	reg [31:0] r_11_0;
	reg [31:0] r_12_0;
	reg [31:0] r_13_0;
	reg [31:0] r_14_0;
	reg [31:0] r_15_0;
	reg [31:0] r_16_0;
	reg [31:0] r_17_0;
	reg [31:0] r_18_0;
	reg [31:0] r_19_0;
	reg [31:0] r_20_0;
	reg [31:0] r_21_0;
	reg [31:0] r_22_0;
	reg [31:0] r_23_0;
	reg [31:0] r_24_0;
	reg [31:0] r_25_0;
	reg [31:0] r_26_0;
	reg [31:0] r_27_0;
	reg [31:0] r_28_0;
	reg [31:0] r_29_0;
	reg [31:0] r_30_0;
	reg [31:0] r_31_0;
	reg [31:0] r_32_0;
	reg [31:0] r_33_0;
	reg [31:0] r_34_0;
	reg [31:0] r_35_0;
	reg [31:0] r_36_0;
	reg [31:0] r_37_0;
	reg [31:0] r_38_0;
	reg [31:0] r_39_0;
	reg [31:0] r_40_0;
	reg [31:0] r_41_0;
	reg [31:0] r_42_0;
	reg [31:0] r_43_0;
	reg [31:0] r_44_0;
	reg [31:0] r_45_0;
	reg [31:0] r_46_0;
	reg [31:0] r_47_0;
	reg [31:0] r_48_0;
	reg [31:0] r_49_0;
	reg [31:0] r_50_0;
	reg [31:0] r_51_0;
	reg [31:0] r_52_0;
	reg [31:0] r_53_0;
	reg [31:0] r_54_0;
	reg [31:0] r_55_0;
	reg [31:0] r_56_0;
	reg [31:0] r_57_0;
	reg [31:0] r_58_0;
	reg [31:0] r_59_0;
	reg [31:0] r_60_0;
	reg [31:0] r_61_0;
	reg [31:0] r_62_0;
	reg [31:0] r_63_0;
	reg [31:0] r_64_0;
	reg [31:0] r_65_0;
	reg [31:0] r_66_0;
	reg [31:0] r_67_0;
	reg [31:0] r_68_0;
	reg [31:0] r_69_0;
	reg [31:0] r_70_0;
	reg [31:0] r_71_0;
	reg [31:0] r_72_0;
	reg [31:0] r_73_0;
	reg [31:0] r_74_0;
	reg [31:0] r_75_0;
	reg [31:0] r_76_0;
	reg [31:0] r_77_0;
	reg [31:0] r_78_0;
	reg [31:0] r_79_0;
	reg [31:0] r_80_0;
	reg [31:0] r_81_0;
	reg [31:0] r_82_0;
	reg [31:0] r_83_0;
	reg [31:0] r_84_0;
	reg [31:0] r_85_0;
	reg [31:0] r_86_0;
	reg [31:0] r_87_0;
	reg [31:0] r_88_0;
	reg [31:0] r_89_0;
	reg [31:0] r_90_0;
	reg [31:0] r_91_0;
	reg [31:0] r_92_0;
	reg [31:0] r_93_0;
	reg [31:0] r_94_0;
	reg [31:0] r_95_0;
	reg [31:0] r_96_0;
	reg [31:0] r_97_0;
	reg [31:0] r_98_0;
	reg [31:0] r_99_0;
	reg [31:0] r_100_0;
	reg [31:0] r_101_0;
	reg [31:0] r_102_0;
	reg [31:0] r_103_0;
	reg [31:0] r_104_0;
	reg [31:0] r_105_0;
	reg [31:0] r_106_0;
	reg [31:0] r_107_0;
	reg [31:0] r_108_0;
	reg [31:0] r_109_0;
	reg [31:0] r_110_0;
	reg [31:0] r_111_0;
	reg [31:0] r_112_0;
	reg [31:0] r_113_0;
	reg [31:0] r_114_0;
	reg [31:0] r_115_0;
	reg [31:0] r_116_0;
	reg [31:0] r_117_0;
	reg [31:0] r_118_0;
	reg [31:0] r_119_0;
	reg [31:0] r_120_0;
	reg [31:0] r_121_0;
	reg [31:0] r_122_0;
	reg [31:0] r_123_0;
	reg [31:0] r_124_0;
	reg [31:0] r_125_0;
	reg [31:0] r_126_0;
	reg [31:0] r_127_0;
	reg [31:0] r_128_0;
	reg [31:0] r_129_0;
	reg [31:0] r_130_0;
	reg [31:0] r_131_0;
	reg [31:0] r_132_0;
	reg [31:0] r_133_0;
	reg [31:0] r_134_0;
	reg [31:0] r_135_0;
	reg [31:0] r_136_0;
	reg [31:0] r_137_0;
	reg [31:0] r_138_0;
	reg [31:0] r_139_0;
	reg [31:0] r_140_0;
	reg [31:0] r_141_0;
	reg [31:0] r_142_0;
	reg [31:0] r_143_0;
	reg [31:0] r_144_0;
	reg [31:0] r_145_0;
	reg [31:0] r_146_0;
	reg [31:0] r_147_0;
	reg [31:0] r_148_0;
	reg [31:0] r_149_0;
	reg [31:0] r_150_0;
	reg [31:0] r_151_0;
	reg [31:0] r_152_0;
	reg [31:0] r_153_0;
	reg [31:0] r_154_0;
	reg [31:0] r_155_0;
	reg [31:0] r_156_0;
	reg [31:0] r_157_0;
	reg [31:0] r_158_0;
	reg [31:0] r_159_0;
	reg [31:0] r_160_0;
	reg [31:0] r_161_0;
	reg [31:0] r_162_0;
	reg [31:0] r_163_0;
	reg [31:0] r_164_0;
	reg [31:0] r_165_0;
	reg [31:0] r_166_0;
	reg [31:0] r_167_0;
	reg [31:0] r_168_0;
	reg [31:0] r_169_0;
	reg [31:0] r_170_0;
	reg [31:0] r_171_0;
	reg [31:0] r_172_0;
	reg [31:0] r_173_0;
	reg [31:0] r_174_0;
	reg [31:0] r_175_0;
	reg [31:0] r_176_0;
	reg [31:0] r_177_0;
	reg [31:0] r_178_0;
	reg [31:0] r_179_0;
	reg [31:0] r_180_0;
	reg [31:0] r_181_0;
	reg [31:0] r_182_0;
	reg [31:0] r_183_0;
	reg [31:0] r_184_0;
	reg [31:0] r_185_0;
	reg [31:0] r_186_0;
	reg [31:0] r_187_0;
	reg [31:0] r_188_0;
	reg [31:0] r_189_0;
	reg [31:0] r_190_0;
	reg [31:0] r_191_0;
	reg [31:0] r_192_0;
	reg [31:0] r_193_0;
	reg [31:0] r_194_0;
	reg [31:0] r_195_0;
	reg [31:0] r_196_0;
	reg [31:0] r_197_0;
	reg [31:0] r_198_0;
	reg [31:0] r_199_0;
	reg [31:0] r_200_0;
	reg [31:0] r_201_0;
	reg [31:0] r_202_0;
	reg [31:0] r_203_0;
	reg [31:0] r_204_0;
	reg [31:0] r_205_0;
	reg [31:0] r_206_0;
	reg [31:0] r_207_0;
	reg [31:0] r_208_0;
	reg [31:0] r_209_0;
	reg [31:0] r_210_0;
	reg [31:0] r_211_0;
	reg [31:0] r_212_0;
	reg [31:0] r_213_0;
	reg [31:0] r_214_0;
	reg [31:0] r_215_0;
	reg [31:0] r_216_0;
	reg [31:0] r_217_0;
	reg [31:0] r_218_0;
	reg [31:0] r_219_0;
	reg [31:0] r_220_0;
	reg [31:0] r_221_0;
	reg [31:0] r_222_0;
	reg [31:0] r_223_0;
	reg [31:0] r_224_0;
	reg [31:0] r_225_0;
	reg [31:0] r_226_0;
	reg [31:0] r_227_0;
	reg [31:0] r_228_0;
	reg [31:0] r_229_0;
	reg [31:0] r_230_0;
	reg [31:0] r_231_0;
	reg [31:0] r_232_0;
	reg [31:0] r_233_0;
	reg [31:0] r_234_0;
	reg [31:0] r_235_0;
	reg [31:0] r_236_0;
	reg [31:0] r_237_0;
	reg [31:0] r_238_0;
	reg [31:0] r_239_0;
	reg [31:0] r_240_0;
	reg [31:0] r_241_0;
	reg [31:0] r_242_0;
	reg [31:0] r_243_0;
	reg [31:0] r_244_0;
	reg [31:0] r_245_0;
	reg [31:0] r_246_0;
	reg [31:0] r_247_0;
	reg [31:0] r_248_0;
	reg [31:0] r_249_0;
	reg [31:0] r_250_0;
	reg [31:0] r_251_0;
	reg [31:0] r_252_0;
	reg [31:0] r_253_0;
	reg [31:0] r_254_0;
	reg [31:0] r_255_0;
	reg [31:0] b_0;
	reg [31:0] b_1_0;
	reg [31:0] b_2_0;
	reg [31:0] b_3_0;
	reg [31:0] b_4_0;
	reg [31:0] b_5_0;
	reg [31:0] b_6_0;
	reg [31:0] b_7_0;
	reg [31:0] b_8_0;
	reg [31:0] b_9_0;
	reg [31:0] b_10_0;
	reg [31:0] b_11_0;
	reg [31:0] b_12_0;
	reg [31:0] b_13_0;
	reg [31:0] b_14_0;
	reg [31:0] b_15_0;
	reg [31:0] b_16_0;
	reg [31:0] b_17_0;
	reg [31:0] b_18_0;
	reg [31:0] b_19_0;
	reg [31:0] b_20_0;
	reg [31:0] b_21_0;
	reg [31:0] b_22_0;
	reg [31:0] b_23_0;
	reg [31:0] b_24_0;
	reg [31:0] b_25_0;
	reg [31:0] b_26_0;
	reg [31:0] b_27_0;
	reg [31:0] b_28_0;
	reg [31:0] b_29_0;
	reg [31:0] b_30_0;
	reg [31:0] b_31_0;
	reg [31:0] b_32_0;
	reg [31:0] b_33_0;
	reg [31:0] b_34_0;
	reg [31:0] b_35_0;
	reg [31:0] b_36_0;
	reg [31:0] b_37_0;
	reg [31:0] b_38_0;
	reg [31:0] b_39_0;
	reg [31:0] b_40_0;
	reg [31:0] b_41_0;
	reg [31:0] b_42_0;
	reg [31:0] b_43_0;
	reg [31:0] b_44_0;
	reg [31:0] b_45_0;
	reg [31:0] b_46_0;
	reg [31:0] b_47_0;
	reg [31:0] b_48_0;
	reg [31:0] b_49_0;
	reg [31:0] b_50_0;
	reg [31:0] b_51_0;
	reg [31:0] b_52_0;
	reg [31:0] b_53_0;
	reg [31:0] b_54_0;
	reg [31:0] b_55_0;
	reg [31:0] b_56_0;
	reg [31:0] b_57_0;
	reg [31:0] b_58_0;
	reg [31:0] b_59_0;
	reg [31:0] b_60_0;
	reg [31:0] b_61_0;
	reg [31:0] b_62_0;
	reg [31:0] b_63_0;
	reg [31:0] b_64_0;
	reg [31:0] b_65_0;
	reg [31:0] b_66_0;
	reg [31:0] b_67_0;
	reg [31:0] b_68_0;
	reg [31:0] b_69_0;
	reg [31:0] b_70_0;
	reg [31:0] b_71_0;
	reg [31:0] b_72_0;
	reg [31:0] b_73_0;
	reg [31:0] b_74_0;
	reg [31:0] b_75_0;
	reg [31:0] b_76_0;
	reg [31:0] b_77_0;
	reg [31:0] b_78_0;
	reg [31:0] b_79_0;
	reg [31:0] b_80_0;
	reg [31:0] b_81_0;
	reg [31:0] b_82_0;
	reg [31:0] b_83_0;
	reg [31:0] b_84_0;
	reg [31:0] b_85_0;
	reg [31:0] b_86_0;
	reg [31:0] b_87_0;
	reg [31:0] b_88_0;
	reg [31:0] b_89_0;
	reg [31:0] b_90_0;
	reg [31:0] b_91_0;
	reg [31:0] b_92_0;
	reg [31:0] b_93_0;
	reg [31:0] b_94_0;
	reg [31:0] b_95_0;
	reg [31:0] b_96_0;
	reg [31:0] b_97_0;
	reg [31:0] b_98_0;
	reg [31:0] b_99_0;
	reg [31:0] b_100_0;
	reg [31:0] b_101_0;
	reg [31:0] b_102_0;
	reg [31:0] b_103_0;
	reg [31:0] b_104_0;
	reg [31:0] b_105_0;
	reg [31:0] b_106_0;
	reg [31:0] b_107_0;
	reg [31:0] b_108_0;
	reg [31:0] b_109_0;
	reg [31:0] b_110_0;
	reg [31:0] b_111_0;
	reg [31:0] b_112_0;
	reg [31:0] b_113_0;
	reg [31:0] b_114_0;
	reg [31:0] b_115_0;
	reg [31:0] b_116_0;
	reg [31:0] b_117_0;
	reg [31:0] b_118_0;
	reg [31:0] b_119_0;
	reg [31:0] b_120_0;
	reg [31:0] b_121_0;
	reg [31:0] b_122_0;
	reg [31:0] b_123_0;
	reg [31:0] b_124_0;
	reg [31:0] b_125_0;
	reg [31:0] b_126_0;
	reg [31:0] b_127_0;
	reg [31:0] b_128_0;
	reg [31:0] b_129_0;
	reg [31:0] b_130_0;
	reg [31:0] b_131_0;
	reg [31:0] b_132_0;
	reg [31:0] b_133_0;
	reg [31:0] b_134_0;
	reg [31:0] b_135_0;
	reg [31:0] b_136_0;
	reg [31:0] b_137_0;
	reg [31:0] b_138_0;
	reg [31:0] b_139_0;
	reg [31:0] b_140_0;
	reg [31:0] b_141_0;
	reg [31:0] b_142_0;
	reg [31:0] b_143_0;
	reg [31:0] b_144_0;
	reg [31:0] b_145_0;
	reg [31:0] b_146_0;
	reg [31:0] b_147_0;
	reg [31:0] b_148_0;
	reg [31:0] b_149_0;
	reg [31:0] b_150_0;
	reg [31:0] b_151_0;
	reg [31:0] b_152_0;
	reg [31:0] b_153_0;
	reg [31:0] b_154_0;
	reg [31:0] b_155_0;
	reg [31:0] b_156_0;
	reg [31:0] b_157_0;
	reg [31:0] b_158_0;
	reg [31:0] b_159_0;
	reg [31:0] b_160_0;
	reg [31:0] b_161_0;
	reg [31:0] b_162_0;
	reg [31:0] b_163_0;
	reg [31:0] b_164_0;
	reg [31:0] b_165_0;
	reg [31:0] b_166_0;
	reg [31:0] b_167_0;
	reg [31:0] b_168_0;
	reg [31:0] b_169_0;
	reg [31:0] b_170_0;
	reg [31:0] b_171_0;
	reg [31:0] b_172_0;
	reg [31:0] b_173_0;
	reg [31:0] b_174_0;
	reg [31:0] b_175_0;
	reg [31:0] b_176_0;
	reg [31:0] b_177_0;
	reg [31:0] b_178_0;
	reg [31:0] b_179_0;
	reg [31:0] b_180_0;
	reg [31:0] b_181_0;
	reg [31:0] b_182_0;
	reg [31:0] b_183_0;
	reg [31:0] b_184_0;
	reg [31:0] b_185_0;
	reg [31:0] b_186_0;
	reg [31:0] b_187_0;
	reg [31:0] b_188_0;
	reg [31:0] b_189_0;
	reg [31:0] b_190_0;
	reg [31:0] b_191_0;
	reg [31:0] b_192_0;
	reg [31:0] b_193_0;
	reg [31:0] b_194_0;
	reg [31:0] b_195_0;
	reg [31:0] b_196_0;
	reg [31:0] b_197_0;
	reg [31:0] b_198_0;
	reg [31:0] b_199_0;
	reg [31:0] b_200_0;
	reg [31:0] b_201_0;
	reg [31:0] b_202_0;
	reg [31:0] b_203_0;
	reg [31:0] b_204_0;
	reg [31:0] b_205_0;
	reg [31:0] b_206_0;
	reg [31:0] b_207_0;
	reg [31:0] b_208_0;
	reg [31:0] b_209_0;
	reg [31:0] b_210_0;
	reg [31:0] b_211_0;
	reg [31:0] b_212_0;
	reg [31:0] b_213_0;
	reg [31:0] b_214_0;
	reg [31:0] b_215_0;
	reg [31:0] b_216_0;
	reg [31:0] b_217_0;
	reg [31:0] b_218_0;
	reg [31:0] b_219_0;
	reg [31:0] b_220_0;
	reg [31:0] b_221_0;
	reg [31:0] b_222_0;
	reg [31:0] b_223_0;
	reg [31:0] b_224_0;
	reg [31:0] b_225_0;
	reg [31:0] b_226_0;
	reg [31:0] b_227_0;
	reg [31:0] b_228_0;
	reg [31:0] b_229_0;
	reg [31:0] b_230_0;
	reg [31:0] b_231_0;
	reg [31:0] b_232_0;
	reg [31:0] b_233_0;
	reg [31:0] b_234_0;
	reg [31:0] b_235_0;
	reg [31:0] b_236_0;
	reg [31:0] b_237_0;
	reg [31:0] b_238_0;
	reg [31:0] b_239_0;
	reg [31:0] b_240_0;
	reg [31:0] b_241_0;
	reg [31:0] b_242_0;
	reg [31:0] b_243_0;
	reg [31:0] b_244_0;
	reg [31:0] b_245_0;
	reg [31:0] b_246_0;
	reg [31:0] b_247_0;
	reg [31:0] b_248_0;
	reg [31:0] b_249_0;
	reg [31:0] b_250_0;
	reg [31:0] b_251_0;
	reg [31:0] b_252_0;
	reg [31:0] b_253_0;
	reg [31:0] b_254_0;
	reg [31:0] b_255_0;
	reg [31:0] b_256_0;
	reg [31:0] b_257_0;
	reg [31:0] b_258_0;
	reg [31:0] b_259_0;
	reg [31:0] b_260_0;
	reg [31:0] b_261_0;
	reg [31:0] b_262_0;
	reg [31:0] b_263_0;
	reg [31:0] b_264_0;
	reg [31:0] b_265_0;
	reg [31:0] b_266_0;
	reg [31:0] b_267_0;
	reg [31:0] b_268_0;
	reg [31:0] b_269_0;
	reg [31:0] b_270_0;
	reg [31:0] b_271_0;
	reg [31:0] b_272_0;
	reg [31:0] b_273_0;
	reg [31:0] b_274_0;
	reg [31:0] b_275_0;
	reg [31:0] b_276_0;
	reg [31:0] b_277_0;
	reg [31:0] b_278_0;
	reg [31:0] b_279_0;
	reg [31:0] b_280_0;
	reg [31:0] b_281_0;
	reg [31:0] b_282_0;
	reg [31:0] b_283_0;
	reg [31:0] b_284_0;
	reg [31:0] b_285_0;
	reg [31:0] b_286_0;
	reg [31:0] b_287_0;
	reg [31:0] b_288_0;
	reg [31:0] b_289_0;
	reg [31:0] b_290_0;
	reg [31:0] b_291_0;
	reg [31:0] b_292_0;
	reg [31:0] b_293_0;
	reg [31:0] b_294_0;
	reg [31:0] b_295_0;
	reg [31:0] b_296_0;
	reg [31:0] b_297_0;
	reg [31:0] b_298_0;
	reg [31:0] b_299_0;
	reg [31:0] b_300_0;
	reg [31:0] b_301_0;
	reg [31:0] b_302_0;
	reg [31:0] b_303_0;
	reg [31:0] b_304_0;
	reg [31:0] b_305_0;
	reg [31:0] b_306_0;
	reg [31:0] b_307_0;
	reg [31:0] b_308_0;
	reg [31:0] b_309_0;
	reg [31:0] b_310_0;
	reg [31:0] b_311_0;
	reg [31:0] b_312_0;
	reg [31:0] b_313_0;
	reg [31:0] b_314_0;
	reg [31:0] b_315_0;
	reg [31:0] b_316_0;
	reg [31:0] b_317_0;
	reg [31:0] b_318_0;
	reg [31:0] b_319_0;
	reg [31:0] b_320_0;
	reg [31:0] b_321_0;
	reg [31:0] b_322_0;
	reg [31:0] b_323_0;
	reg [31:0] b_324_0;
	reg [31:0] b_325_0;
	reg [31:0] b_326_0;
	reg [31:0] b_327_0;
	reg [31:0] b_328_0;
	reg [31:0] b_329_0;
	reg [31:0] b_330_0;
	reg [31:0] b_331_0;
	reg [31:0] b_332_0;
	reg [31:0] b_333_0;
	reg [31:0] b_334_0;
	reg [31:0] b_335_0;
	reg [31:0] b_336_0;
	reg [31:0] b_337_0;
	reg [31:0] b_338_0;
	reg [31:0] b_339_0;
	reg [31:0] b_340_0;
	reg [31:0] b_341_0;
	reg [31:0] b_342_0;
	reg [31:0] b_343_0;
	reg [31:0] b_344_0;
	reg [31:0] b_345_0;
	reg [31:0] b_346_0;
	reg [31:0] b_347_0;
	reg [31:0] b_348_0;
	reg [31:0] b_349_0;
	reg [31:0] b_350_0;
	reg [31:0] b_351_0;
	reg [31:0] b_352_0;
	reg [31:0] b_353_0;
	reg [31:0] b_354_0;
	reg [31:0] b_355_0;
	reg [31:0] b_356_0;
	reg [31:0] b_357_0;
	reg [31:0] b_358_0;
	reg [31:0] b_359_0;
	reg [31:0] b_360_0;
	reg [31:0] b_361_0;
	reg [31:0] b_362_0;
	reg [31:0] b_363_0;
	reg [31:0] b_364_0;
	reg [31:0] b_365_0;
	reg [31:0] b_366_0;
	reg [31:0] b_367_0;
	reg [31:0] b_368_0;
	reg [31:0] b_369_0;
	reg [31:0] b_370_0;
	reg [31:0] b_371_0;
	reg [31:0] b_372_0;
	reg [31:0] b_373_0;
	reg [31:0] b_374_0;
	reg [31:0] b_375_0;
	reg [31:0] b_376_0;
	reg [31:0] b_377_0;
	reg [31:0] b_378_0;
	reg [31:0] b_379_0;
	reg [31:0] b_380_0;
	reg [31:0] b_381_0;
	reg [31:0] b_382_0;
	reg [31:0] b_383_0;
	reg [31:0] b_384_0;
	reg [31:0] b_385_0;
	reg [31:0] b_386_0;
	reg [31:0] b_387_0;
	reg [31:0] b_388_0;
	reg [31:0] b_389_0;
	reg [31:0] b_390_0;
	reg [31:0] b_391_0;
	reg [31:0] b_392_0;
	reg [31:0] b_393_0;
	reg [31:0] b_394_0;
	reg [31:0] b_395_0;
	reg [31:0] b_396_0;
	reg [31:0] b_397_0;
	reg [31:0] b_398_0;
	reg [31:0] b_399_0;
	reg [31:0] b_400_0;
	reg [31:0] b_401_0;
	reg [31:0] b_402_0;
	reg [31:0] b_403_0;
	reg [31:0] b_404_0;
	reg [31:0] b_405_0;
	reg [31:0] b_406_0;
	reg [31:0] b_407_0;
	reg [31:0] b_408_0;
	reg [31:0] b_409_0;
	reg [31:0] b_410_0;
	reg [31:0] b_411_0;
	reg [31:0] b_412_0;
	reg [31:0] b_413_0;
	reg [31:0] b_414_0;
	reg [31:0] b_415_0;
	reg [31:0] b_416_0;
	reg [31:0] b_417_0;
	reg [31:0] b_418_0;
	reg [31:0] b_419_0;
	reg [31:0] b_420_0;
	reg [31:0] b_421_0;
	reg [31:0] b_422_0;
	reg [31:0] b_423_0;
	reg [31:0] b_424_0;
	reg [31:0] b_425_0;
	reg [31:0] b_426_0;
	reg [31:0] b_427_0;
	reg [31:0] b_428_0;
	reg [31:0] b_429_0;
	reg [31:0] b_430_0;
	reg [31:0] b_431_0;
	reg [31:0] b_432_0;
	reg [31:0] b_433_0;
	reg [31:0] b_434_0;
	reg [31:0] b_435_0;
	reg [31:0] b_436_0;
	reg [31:0] b_437_0;
	reg [31:0] b_438_0;
	reg [31:0] b_439_0;
	reg [31:0] b_440_0;
	reg [31:0] b_441_0;
	reg [31:0] b_442_0;
	reg [31:0] b_443_0;
	reg [31:0] b_444_0;
	reg [31:0] b_445_0;
	reg [31:0] b_446_0;
	reg [31:0] b_447_0;
	reg [31:0] b_448_0;
	reg [31:0] b_449_0;
	reg [31:0] b_450_0;
	reg [31:0] b_451_0;
	reg [31:0] b_452_0;
	reg [31:0] b_453_0;
	reg [31:0] b_454_0;
	reg [31:0] b_455_0;
	reg [31:0] b_456_0;
	reg [31:0] b_457_0;
	reg [31:0] b_458_0;
	reg [31:0] b_459_0;
	reg [31:0] b_460_0;
	reg [31:0] b_461_0;
	reg [31:0] b_462_0;
	reg [31:0] b_463_0;
	reg [31:0] b_464_0;
	reg [31:0] b_465_0;
	reg [31:0] b_466_0;
	reg [31:0] b_467_0;
	reg [31:0] b_468_0;
	reg [31:0] b_469_0;
	reg [31:0] b_470_0;
	reg [31:0] b_471_0;
	reg [31:0] b_472_0;
	reg [31:0] b_473_0;
	reg [31:0] b_474_0;
	reg [31:0] b_475_0;
	reg [31:0] b_476_0;
	reg [31:0] b_477_0;
	reg [31:0] b_478_0;
	reg [31:0] b_479_0;
	reg [31:0] b_480_0;
	reg [31:0] b_481_0;
	reg [31:0] b_482_0;
	reg [31:0] b_483_0;
	reg [31:0] b_484_0;
	reg [31:0] b_485_0;
	reg [31:0] b_486_0;
	reg [31:0] b_487_0;
	reg [31:0] b_488_0;
	reg [31:0] b_489_0;
	reg [31:0] b_490_0;
	reg [31:0] b_491_0;
	reg [31:0] b_492_0;
	reg [31:0] b_493_0;
	reg [31:0] b_494_0;
	reg [31:0] b_495_0;
	reg [31:0] b_496_0;
	reg [31:0] b_497_0;
	reg [31:0] b_498_0;
	reg [31:0] b_499_0;
	reg [31:0] b_500_0;
	reg [31:0] b_501_0;
	reg [31:0] b_502_0;
	reg [31:0] b_503_0;
	reg [31:0] b_504_0;
	reg [31:0] b_505_0;
	reg [31:0] b_506_0;
	reg [31:0] b_507_0;
	reg [31:0] b_508_0;
	reg [31:0] b_509_0;
	reg [31:0] b_510_0;
	reg [31:0] b_511_0;
	reg [4:0] mesh_0_0_io_in_control_0_shift_b;
	reg mesh_0_0_io_in_control_0_dataflow_b;
	reg mesh_0_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_0_io_in_control_0_shift_b;
	reg mesh_1_0_io_in_control_0_dataflow_b;
	reg mesh_1_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_0_io_in_control_0_shift_b;
	reg mesh_2_0_io_in_control_0_dataflow_b;
	reg mesh_2_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_0_io_in_control_0_shift_b;
	reg mesh_3_0_io_in_control_0_dataflow_b;
	reg mesh_3_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_0_io_in_control_0_shift_b;
	reg mesh_4_0_io_in_control_0_dataflow_b;
	reg mesh_4_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_0_io_in_control_0_shift_b;
	reg mesh_5_0_io_in_control_0_dataflow_b;
	reg mesh_5_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_0_io_in_control_0_shift_b;
	reg mesh_6_0_io_in_control_0_dataflow_b;
	reg mesh_6_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_0_io_in_control_0_shift_b;
	reg mesh_7_0_io_in_control_0_dataflow_b;
	reg mesh_7_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_0_io_in_control_0_shift_b;
	reg mesh_8_0_io_in_control_0_dataflow_b;
	reg mesh_8_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_0_io_in_control_0_shift_b;
	reg mesh_9_0_io_in_control_0_dataflow_b;
	reg mesh_9_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_0_io_in_control_0_shift_b;
	reg mesh_10_0_io_in_control_0_dataflow_b;
	reg mesh_10_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_0_io_in_control_0_shift_b;
	reg mesh_11_0_io_in_control_0_dataflow_b;
	reg mesh_11_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_0_io_in_control_0_shift_b;
	reg mesh_12_0_io_in_control_0_dataflow_b;
	reg mesh_12_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_0_io_in_control_0_shift_b;
	reg mesh_13_0_io_in_control_0_dataflow_b;
	reg mesh_13_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_0_io_in_control_0_shift_b;
	reg mesh_14_0_io_in_control_0_dataflow_b;
	reg mesh_14_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_0_io_in_control_0_shift_b;
	reg mesh_15_0_io_in_control_0_dataflow_b;
	reg mesh_15_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_1_io_in_control_0_shift_b;
	reg mesh_0_1_io_in_control_0_dataflow_b;
	reg mesh_0_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_1_io_in_control_0_shift_b;
	reg mesh_1_1_io_in_control_0_dataflow_b;
	reg mesh_1_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_1_io_in_control_0_shift_b;
	reg mesh_2_1_io_in_control_0_dataflow_b;
	reg mesh_2_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_1_io_in_control_0_shift_b;
	reg mesh_3_1_io_in_control_0_dataflow_b;
	reg mesh_3_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_1_io_in_control_0_shift_b;
	reg mesh_4_1_io_in_control_0_dataflow_b;
	reg mesh_4_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_1_io_in_control_0_shift_b;
	reg mesh_5_1_io_in_control_0_dataflow_b;
	reg mesh_5_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_1_io_in_control_0_shift_b;
	reg mesh_6_1_io_in_control_0_dataflow_b;
	reg mesh_6_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_1_io_in_control_0_shift_b;
	reg mesh_7_1_io_in_control_0_dataflow_b;
	reg mesh_7_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_1_io_in_control_0_shift_b;
	reg mesh_8_1_io_in_control_0_dataflow_b;
	reg mesh_8_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_1_io_in_control_0_shift_b;
	reg mesh_9_1_io_in_control_0_dataflow_b;
	reg mesh_9_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_1_io_in_control_0_shift_b;
	reg mesh_10_1_io_in_control_0_dataflow_b;
	reg mesh_10_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_1_io_in_control_0_shift_b;
	reg mesh_11_1_io_in_control_0_dataflow_b;
	reg mesh_11_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_1_io_in_control_0_shift_b;
	reg mesh_12_1_io_in_control_0_dataflow_b;
	reg mesh_12_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_1_io_in_control_0_shift_b;
	reg mesh_13_1_io_in_control_0_dataflow_b;
	reg mesh_13_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_1_io_in_control_0_shift_b;
	reg mesh_14_1_io_in_control_0_dataflow_b;
	reg mesh_14_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_1_io_in_control_0_shift_b;
	reg mesh_15_1_io_in_control_0_dataflow_b;
	reg mesh_15_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_2_io_in_control_0_shift_b;
	reg mesh_0_2_io_in_control_0_dataflow_b;
	reg mesh_0_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_2_io_in_control_0_shift_b;
	reg mesh_1_2_io_in_control_0_dataflow_b;
	reg mesh_1_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_2_io_in_control_0_shift_b;
	reg mesh_2_2_io_in_control_0_dataflow_b;
	reg mesh_2_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_2_io_in_control_0_shift_b;
	reg mesh_3_2_io_in_control_0_dataflow_b;
	reg mesh_3_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_2_io_in_control_0_shift_b;
	reg mesh_4_2_io_in_control_0_dataflow_b;
	reg mesh_4_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_2_io_in_control_0_shift_b;
	reg mesh_5_2_io_in_control_0_dataflow_b;
	reg mesh_5_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_2_io_in_control_0_shift_b;
	reg mesh_6_2_io_in_control_0_dataflow_b;
	reg mesh_6_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_2_io_in_control_0_shift_b;
	reg mesh_7_2_io_in_control_0_dataflow_b;
	reg mesh_7_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_2_io_in_control_0_shift_b;
	reg mesh_8_2_io_in_control_0_dataflow_b;
	reg mesh_8_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_2_io_in_control_0_shift_b;
	reg mesh_9_2_io_in_control_0_dataflow_b;
	reg mesh_9_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_2_io_in_control_0_shift_b;
	reg mesh_10_2_io_in_control_0_dataflow_b;
	reg mesh_10_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_2_io_in_control_0_shift_b;
	reg mesh_11_2_io_in_control_0_dataflow_b;
	reg mesh_11_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_2_io_in_control_0_shift_b;
	reg mesh_12_2_io_in_control_0_dataflow_b;
	reg mesh_12_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_2_io_in_control_0_shift_b;
	reg mesh_13_2_io_in_control_0_dataflow_b;
	reg mesh_13_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_2_io_in_control_0_shift_b;
	reg mesh_14_2_io_in_control_0_dataflow_b;
	reg mesh_14_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_2_io_in_control_0_shift_b;
	reg mesh_15_2_io_in_control_0_dataflow_b;
	reg mesh_15_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_3_io_in_control_0_shift_b;
	reg mesh_0_3_io_in_control_0_dataflow_b;
	reg mesh_0_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_3_io_in_control_0_shift_b;
	reg mesh_1_3_io_in_control_0_dataflow_b;
	reg mesh_1_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_3_io_in_control_0_shift_b;
	reg mesh_2_3_io_in_control_0_dataflow_b;
	reg mesh_2_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_3_io_in_control_0_shift_b;
	reg mesh_3_3_io_in_control_0_dataflow_b;
	reg mesh_3_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_3_io_in_control_0_shift_b;
	reg mesh_4_3_io_in_control_0_dataflow_b;
	reg mesh_4_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_3_io_in_control_0_shift_b;
	reg mesh_5_3_io_in_control_0_dataflow_b;
	reg mesh_5_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_3_io_in_control_0_shift_b;
	reg mesh_6_3_io_in_control_0_dataflow_b;
	reg mesh_6_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_3_io_in_control_0_shift_b;
	reg mesh_7_3_io_in_control_0_dataflow_b;
	reg mesh_7_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_3_io_in_control_0_shift_b;
	reg mesh_8_3_io_in_control_0_dataflow_b;
	reg mesh_8_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_3_io_in_control_0_shift_b;
	reg mesh_9_3_io_in_control_0_dataflow_b;
	reg mesh_9_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_3_io_in_control_0_shift_b;
	reg mesh_10_3_io_in_control_0_dataflow_b;
	reg mesh_10_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_3_io_in_control_0_shift_b;
	reg mesh_11_3_io_in_control_0_dataflow_b;
	reg mesh_11_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_3_io_in_control_0_shift_b;
	reg mesh_12_3_io_in_control_0_dataflow_b;
	reg mesh_12_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_3_io_in_control_0_shift_b;
	reg mesh_13_3_io_in_control_0_dataflow_b;
	reg mesh_13_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_3_io_in_control_0_shift_b;
	reg mesh_14_3_io_in_control_0_dataflow_b;
	reg mesh_14_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_3_io_in_control_0_shift_b;
	reg mesh_15_3_io_in_control_0_dataflow_b;
	reg mesh_15_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_4_io_in_control_0_shift_b;
	reg mesh_0_4_io_in_control_0_dataflow_b;
	reg mesh_0_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_4_io_in_control_0_shift_b;
	reg mesh_1_4_io_in_control_0_dataflow_b;
	reg mesh_1_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_4_io_in_control_0_shift_b;
	reg mesh_2_4_io_in_control_0_dataflow_b;
	reg mesh_2_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_4_io_in_control_0_shift_b;
	reg mesh_3_4_io_in_control_0_dataflow_b;
	reg mesh_3_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_4_io_in_control_0_shift_b;
	reg mesh_4_4_io_in_control_0_dataflow_b;
	reg mesh_4_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_4_io_in_control_0_shift_b;
	reg mesh_5_4_io_in_control_0_dataflow_b;
	reg mesh_5_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_4_io_in_control_0_shift_b;
	reg mesh_6_4_io_in_control_0_dataflow_b;
	reg mesh_6_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_4_io_in_control_0_shift_b;
	reg mesh_7_4_io_in_control_0_dataflow_b;
	reg mesh_7_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_4_io_in_control_0_shift_b;
	reg mesh_8_4_io_in_control_0_dataflow_b;
	reg mesh_8_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_4_io_in_control_0_shift_b;
	reg mesh_9_4_io_in_control_0_dataflow_b;
	reg mesh_9_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_4_io_in_control_0_shift_b;
	reg mesh_10_4_io_in_control_0_dataflow_b;
	reg mesh_10_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_4_io_in_control_0_shift_b;
	reg mesh_11_4_io_in_control_0_dataflow_b;
	reg mesh_11_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_4_io_in_control_0_shift_b;
	reg mesh_12_4_io_in_control_0_dataflow_b;
	reg mesh_12_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_4_io_in_control_0_shift_b;
	reg mesh_13_4_io_in_control_0_dataflow_b;
	reg mesh_13_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_4_io_in_control_0_shift_b;
	reg mesh_14_4_io_in_control_0_dataflow_b;
	reg mesh_14_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_4_io_in_control_0_shift_b;
	reg mesh_15_4_io_in_control_0_dataflow_b;
	reg mesh_15_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_5_io_in_control_0_shift_b;
	reg mesh_0_5_io_in_control_0_dataflow_b;
	reg mesh_0_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_5_io_in_control_0_shift_b;
	reg mesh_1_5_io_in_control_0_dataflow_b;
	reg mesh_1_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_5_io_in_control_0_shift_b;
	reg mesh_2_5_io_in_control_0_dataflow_b;
	reg mesh_2_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_5_io_in_control_0_shift_b;
	reg mesh_3_5_io_in_control_0_dataflow_b;
	reg mesh_3_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_5_io_in_control_0_shift_b;
	reg mesh_4_5_io_in_control_0_dataflow_b;
	reg mesh_4_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_5_io_in_control_0_shift_b;
	reg mesh_5_5_io_in_control_0_dataflow_b;
	reg mesh_5_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_5_io_in_control_0_shift_b;
	reg mesh_6_5_io_in_control_0_dataflow_b;
	reg mesh_6_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_5_io_in_control_0_shift_b;
	reg mesh_7_5_io_in_control_0_dataflow_b;
	reg mesh_7_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_5_io_in_control_0_shift_b;
	reg mesh_8_5_io_in_control_0_dataflow_b;
	reg mesh_8_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_5_io_in_control_0_shift_b;
	reg mesh_9_5_io_in_control_0_dataflow_b;
	reg mesh_9_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_5_io_in_control_0_shift_b;
	reg mesh_10_5_io_in_control_0_dataflow_b;
	reg mesh_10_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_5_io_in_control_0_shift_b;
	reg mesh_11_5_io_in_control_0_dataflow_b;
	reg mesh_11_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_5_io_in_control_0_shift_b;
	reg mesh_12_5_io_in_control_0_dataflow_b;
	reg mesh_12_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_5_io_in_control_0_shift_b;
	reg mesh_13_5_io_in_control_0_dataflow_b;
	reg mesh_13_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_5_io_in_control_0_shift_b;
	reg mesh_14_5_io_in_control_0_dataflow_b;
	reg mesh_14_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_5_io_in_control_0_shift_b;
	reg mesh_15_5_io_in_control_0_dataflow_b;
	reg mesh_15_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_6_io_in_control_0_shift_b;
	reg mesh_0_6_io_in_control_0_dataflow_b;
	reg mesh_0_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_6_io_in_control_0_shift_b;
	reg mesh_1_6_io_in_control_0_dataflow_b;
	reg mesh_1_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_6_io_in_control_0_shift_b;
	reg mesh_2_6_io_in_control_0_dataflow_b;
	reg mesh_2_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_6_io_in_control_0_shift_b;
	reg mesh_3_6_io_in_control_0_dataflow_b;
	reg mesh_3_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_6_io_in_control_0_shift_b;
	reg mesh_4_6_io_in_control_0_dataflow_b;
	reg mesh_4_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_6_io_in_control_0_shift_b;
	reg mesh_5_6_io_in_control_0_dataflow_b;
	reg mesh_5_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_6_io_in_control_0_shift_b;
	reg mesh_6_6_io_in_control_0_dataflow_b;
	reg mesh_6_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_6_io_in_control_0_shift_b;
	reg mesh_7_6_io_in_control_0_dataflow_b;
	reg mesh_7_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_6_io_in_control_0_shift_b;
	reg mesh_8_6_io_in_control_0_dataflow_b;
	reg mesh_8_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_6_io_in_control_0_shift_b;
	reg mesh_9_6_io_in_control_0_dataflow_b;
	reg mesh_9_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_6_io_in_control_0_shift_b;
	reg mesh_10_6_io_in_control_0_dataflow_b;
	reg mesh_10_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_6_io_in_control_0_shift_b;
	reg mesh_11_6_io_in_control_0_dataflow_b;
	reg mesh_11_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_6_io_in_control_0_shift_b;
	reg mesh_12_6_io_in_control_0_dataflow_b;
	reg mesh_12_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_6_io_in_control_0_shift_b;
	reg mesh_13_6_io_in_control_0_dataflow_b;
	reg mesh_13_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_6_io_in_control_0_shift_b;
	reg mesh_14_6_io_in_control_0_dataflow_b;
	reg mesh_14_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_6_io_in_control_0_shift_b;
	reg mesh_15_6_io_in_control_0_dataflow_b;
	reg mesh_15_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_7_io_in_control_0_shift_b;
	reg mesh_0_7_io_in_control_0_dataflow_b;
	reg mesh_0_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_7_io_in_control_0_shift_b;
	reg mesh_1_7_io_in_control_0_dataflow_b;
	reg mesh_1_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_7_io_in_control_0_shift_b;
	reg mesh_2_7_io_in_control_0_dataflow_b;
	reg mesh_2_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_7_io_in_control_0_shift_b;
	reg mesh_3_7_io_in_control_0_dataflow_b;
	reg mesh_3_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_7_io_in_control_0_shift_b;
	reg mesh_4_7_io_in_control_0_dataflow_b;
	reg mesh_4_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_7_io_in_control_0_shift_b;
	reg mesh_5_7_io_in_control_0_dataflow_b;
	reg mesh_5_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_7_io_in_control_0_shift_b;
	reg mesh_6_7_io_in_control_0_dataflow_b;
	reg mesh_6_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_7_io_in_control_0_shift_b;
	reg mesh_7_7_io_in_control_0_dataflow_b;
	reg mesh_7_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_7_io_in_control_0_shift_b;
	reg mesh_8_7_io_in_control_0_dataflow_b;
	reg mesh_8_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_7_io_in_control_0_shift_b;
	reg mesh_9_7_io_in_control_0_dataflow_b;
	reg mesh_9_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_7_io_in_control_0_shift_b;
	reg mesh_10_7_io_in_control_0_dataflow_b;
	reg mesh_10_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_7_io_in_control_0_shift_b;
	reg mesh_11_7_io_in_control_0_dataflow_b;
	reg mesh_11_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_7_io_in_control_0_shift_b;
	reg mesh_12_7_io_in_control_0_dataflow_b;
	reg mesh_12_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_7_io_in_control_0_shift_b;
	reg mesh_13_7_io_in_control_0_dataflow_b;
	reg mesh_13_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_7_io_in_control_0_shift_b;
	reg mesh_14_7_io_in_control_0_dataflow_b;
	reg mesh_14_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_7_io_in_control_0_shift_b;
	reg mesh_15_7_io_in_control_0_dataflow_b;
	reg mesh_15_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_8_io_in_control_0_shift_b;
	reg mesh_0_8_io_in_control_0_dataflow_b;
	reg mesh_0_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_8_io_in_control_0_shift_b;
	reg mesh_1_8_io_in_control_0_dataflow_b;
	reg mesh_1_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_8_io_in_control_0_shift_b;
	reg mesh_2_8_io_in_control_0_dataflow_b;
	reg mesh_2_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_8_io_in_control_0_shift_b;
	reg mesh_3_8_io_in_control_0_dataflow_b;
	reg mesh_3_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_8_io_in_control_0_shift_b;
	reg mesh_4_8_io_in_control_0_dataflow_b;
	reg mesh_4_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_8_io_in_control_0_shift_b;
	reg mesh_5_8_io_in_control_0_dataflow_b;
	reg mesh_5_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_8_io_in_control_0_shift_b;
	reg mesh_6_8_io_in_control_0_dataflow_b;
	reg mesh_6_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_8_io_in_control_0_shift_b;
	reg mesh_7_8_io_in_control_0_dataflow_b;
	reg mesh_7_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_8_io_in_control_0_shift_b;
	reg mesh_8_8_io_in_control_0_dataflow_b;
	reg mesh_8_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_8_io_in_control_0_shift_b;
	reg mesh_9_8_io_in_control_0_dataflow_b;
	reg mesh_9_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_8_io_in_control_0_shift_b;
	reg mesh_10_8_io_in_control_0_dataflow_b;
	reg mesh_10_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_8_io_in_control_0_shift_b;
	reg mesh_11_8_io_in_control_0_dataflow_b;
	reg mesh_11_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_8_io_in_control_0_shift_b;
	reg mesh_12_8_io_in_control_0_dataflow_b;
	reg mesh_12_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_8_io_in_control_0_shift_b;
	reg mesh_13_8_io_in_control_0_dataflow_b;
	reg mesh_13_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_8_io_in_control_0_shift_b;
	reg mesh_14_8_io_in_control_0_dataflow_b;
	reg mesh_14_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_8_io_in_control_0_shift_b;
	reg mesh_15_8_io_in_control_0_dataflow_b;
	reg mesh_15_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_9_io_in_control_0_shift_b;
	reg mesh_0_9_io_in_control_0_dataflow_b;
	reg mesh_0_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_9_io_in_control_0_shift_b;
	reg mesh_1_9_io_in_control_0_dataflow_b;
	reg mesh_1_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_9_io_in_control_0_shift_b;
	reg mesh_2_9_io_in_control_0_dataflow_b;
	reg mesh_2_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_9_io_in_control_0_shift_b;
	reg mesh_3_9_io_in_control_0_dataflow_b;
	reg mesh_3_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_9_io_in_control_0_shift_b;
	reg mesh_4_9_io_in_control_0_dataflow_b;
	reg mesh_4_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_9_io_in_control_0_shift_b;
	reg mesh_5_9_io_in_control_0_dataflow_b;
	reg mesh_5_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_9_io_in_control_0_shift_b;
	reg mesh_6_9_io_in_control_0_dataflow_b;
	reg mesh_6_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_9_io_in_control_0_shift_b;
	reg mesh_7_9_io_in_control_0_dataflow_b;
	reg mesh_7_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_9_io_in_control_0_shift_b;
	reg mesh_8_9_io_in_control_0_dataflow_b;
	reg mesh_8_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_9_io_in_control_0_shift_b;
	reg mesh_9_9_io_in_control_0_dataflow_b;
	reg mesh_9_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_9_io_in_control_0_shift_b;
	reg mesh_10_9_io_in_control_0_dataflow_b;
	reg mesh_10_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_9_io_in_control_0_shift_b;
	reg mesh_11_9_io_in_control_0_dataflow_b;
	reg mesh_11_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_9_io_in_control_0_shift_b;
	reg mesh_12_9_io_in_control_0_dataflow_b;
	reg mesh_12_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_9_io_in_control_0_shift_b;
	reg mesh_13_9_io_in_control_0_dataflow_b;
	reg mesh_13_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_9_io_in_control_0_shift_b;
	reg mesh_14_9_io_in_control_0_dataflow_b;
	reg mesh_14_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_9_io_in_control_0_shift_b;
	reg mesh_15_9_io_in_control_0_dataflow_b;
	reg mesh_15_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_10_io_in_control_0_shift_b;
	reg mesh_0_10_io_in_control_0_dataflow_b;
	reg mesh_0_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_10_io_in_control_0_shift_b;
	reg mesh_1_10_io_in_control_0_dataflow_b;
	reg mesh_1_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_10_io_in_control_0_shift_b;
	reg mesh_2_10_io_in_control_0_dataflow_b;
	reg mesh_2_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_10_io_in_control_0_shift_b;
	reg mesh_3_10_io_in_control_0_dataflow_b;
	reg mesh_3_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_10_io_in_control_0_shift_b;
	reg mesh_4_10_io_in_control_0_dataflow_b;
	reg mesh_4_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_10_io_in_control_0_shift_b;
	reg mesh_5_10_io_in_control_0_dataflow_b;
	reg mesh_5_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_10_io_in_control_0_shift_b;
	reg mesh_6_10_io_in_control_0_dataflow_b;
	reg mesh_6_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_10_io_in_control_0_shift_b;
	reg mesh_7_10_io_in_control_0_dataflow_b;
	reg mesh_7_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_10_io_in_control_0_shift_b;
	reg mesh_8_10_io_in_control_0_dataflow_b;
	reg mesh_8_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_10_io_in_control_0_shift_b;
	reg mesh_9_10_io_in_control_0_dataflow_b;
	reg mesh_9_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_10_io_in_control_0_shift_b;
	reg mesh_10_10_io_in_control_0_dataflow_b;
	reg mesh_10_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_10_io_in_control_0_shift_b;
	reg mesh_11_10_io_in_control_0_dataflow_b;
	reg mesh_11_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_10_io_in_control_0_shift_b;
	reg mesh_12_10_io_in_control_0_dataflow_b;
	reg mesh_12_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_10_io_in_control_0_shift_b;
	reg mesh_13_10_io_in_control_0_dataflow_b;
	reg mesh_13_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_10_io_in_control_0_shift_b;
	reg mesh_14_10_io_in_control_0_dataflow_b;
	reg mesh_14_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_10_io_in_control_0_shift_b;
	reg mesh_15_10_io_in_control_0_dataflow_b;
	reg mesh_15_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_11_io_in_control_0_shift_b;
	reg mesh_0_11_io_in_control_0_dataflow_b;
	reg mesh_0_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_11_io_in_control_0_shift_b;
	reg mesh_1_11_io_in_control_0_dataflow_b;
	reg mesh_1_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_11_io_in_control_0_shift_b;
	reg mesh_2_11_io_in_control_0_dataflow_b;
	reg mesh_2_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_11_io_in_control_0_shift_b;
	reg mesh_3_11_io_in_control_0_dataflow_b;
	reg mesh_3_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_11_io_in_control_0_shift_b;
	reg mesh_4_11_io_in_control_0_dataflow_b;
	reg mesh_4_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_11_io_in_control_0_shift_b;
	reg mesh_5_11_io_in_control_0_dataflow_b;
	reg mesh_5_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_11_io_in_control_0_shift_b;
	reg mesh_6_11_io_in_control_0_dataflow_b;
	reg mesh_6_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_11_io_in_control_0_shift_b;
	reg mesh_7_11_io_in_control_0_dataflow_b;
	reg mesh_7_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_11_io_in_control_0_shift_b;
	reg mesh_8_11_io_in_control_0_dataflow_b;
	reg mesh_8_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_11_io_in_control_0_shift_b;
	reg mesh_9_11_io_in_control_0_dataflow_b;
	reg mesh_9_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_11_io_in_control_0_shift_b;
	reg mesh_10_11_io_in_control_0_dataflow_b;
	reg mesh_10_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_11_io_in_control_0_shift_b;
	reg mesh_11_11_io_in_control_0_dataflow_b;
	reg mesh_11_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_11_io_in_control_0_shift_b;
	reg mesh_12_11_io_in_control_0_dataflow_b;
	reg mesh_12_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_11_io_in_control_0_shift_b;
	reg mesh_13_11_io_in_control_0_dataflow_b;
	reg mesh_13_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_11_io_in_control_0_shift_b;
	reg mesh_14_11_io_in_control_0_dataflow_b;
	reg mesh_14_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_11_io_in_control_0_shift_b;
	reg mesh_15_11_io_in_control_0_dataflow_b;
	reg mesh_15_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_12_io_in_control_0_shift_b;
	reg mesh_0_12_io_in_control_0_dataflow_b;
	reg mesh_0_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_12_io_in_control_0_shift_b;
	reg mesh_1_12_io_in_control_0_dataflow_b;
	reg mesh_1_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_12_io_in_control_0_shift_b;
	reg mesh_2_12_io_in_control_0_dataflow_b;
	reg mesh_2_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_12_io_in_control_0_shift_b;
	reg mesh_3_12_io_in_control_0_dataflow_b;
	reg mesh_3_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_12_io_in_control_0_shift_b;
	reg mesh_4_12_io_in_control_0_dataflow_b;
	reg mesh_4_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_12_io_in_control_0_shift_b;
	reg mesh_5_12_io_in_control_0_dataflow_b;
	reg mesh_5_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_12_io_in_control_0_shift_b;
	reg mesh_6_12_io_in_control_0_dataflow_b;
	reg mesh_6_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_12_io_in_control_0_shift_b;
	reg mesh_7_12_io_in_control_0_dataflow_b;
	reg mesh_7_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_12_io_in_control_0_shift_b;
	reg mesh_8_12_io_in_control_0_dataflow_b;
	reg mesh_8_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_12_io_in_control_0_shift_b;
	reg mesh_9_12_io_in_control_0_dataflow_b;
	reg mesh_9_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_12_io_in_control_0_shift_b;
	reg mesh_10_12_io_in_control_0_dataflow_b;
	reg mesh_10_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_12_io_in_control_0_shift_b;
	reg mesh_11_12_io_in_control_0_dataflow_b;
	reg mesh_11_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_12_io_in_control_0_shift_b;
	reg mesh_12_12_io_in_control_0_dataflow_b;
	reg mesh_12_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_12_io_in_control_0_shift_b;
	reg mesh_13_12_io_in_control_0_dataflow_b;
	reg mesh_13_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_12_io_in_control_0_shift_b;
	reg mesh_14_12_io_in_control_0_dataflow_b;
	reg mesh_14_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_12_io_in_control_0_shift_b;
	reg mesh_15_12_io_in_control_0_dataflow_b;
	reg mesh_15_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_13_io_in_control_0_shift_b;
	reg mesh_0_13_io_in_control_0_dataflow_b;
	reg mesh_0_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_13_io_in_control_0_shift_b;
	reg mesh_1_13_io_in_control_0_dataflow_b;
	reg mesh_1_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_13_io_in_control_0_shift_b;
	reg mesh_2_13_io_in_control_0_dataflow_b;
	reg mesh_2_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_13_io_in_control_0_shift_b;
	reg mesh_3_13_io_in_control_0_dataflow_b;
	reg mesh_3_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_13_io_in_control_0_shift_b;
	reg mesh_4_13_io_in_control_0_dataflow_b;
	reg mesh_4_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_13_io_in_control_0_shift_b;
	reg mesh_5_13_io_in_control_0_dataflow_b;
	reg mesh_5_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_13_io_in_control_0_shift_b;
	reg mesh_6_13_io_in_control_0_dataflow_b;
	reg mesh_6_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_13_io_in_control_0_shift_b;
	reg mesh_7_13_io_in_control_0_dataflow_b;
	reg mesh_7_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_13_io_in_control_0_shift_b;
	reg mesh_8_13_io_in_control_0_dataflow_b;
	reg mesh_8_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_13_io_in_control_0_shift_b;
	reg mesh_9_13_io_in_control_0_dataflow_b;
	reg mesh_9_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_13_io_in_control_0_shift_b;
	reg mesh_10_13_io_in_control_0_dataflow_b;
	reg mesh_10_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_13_io_in_control_0_shift_b;
	reg mesh_11_13_io_in_control_0_dataflow_b;
	reg mesh_11_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_13_io_in_control_0_shift_b;
	reg mesh_12_13_io_in_control_0_dataflow_b;
	reg mesh_12_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_13_io_in_control_0_shift_b;
	reg mesh_13_13_io_in_control_0_dataflow_b;
	reg mesh_13_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_13_io_in_control_0_shift_b;
	reg mesh_14_13_io_in_control_0_dataflow_b;
	reg mesh_14_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_13_io_in_control_0_shift_b;
	reg mesh_15_13_io_in_control_0_dataflow_b;
	reg mesh_15_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_14_io_in_control_0_shift_b;
	reg mesh_0_14_io_in_control_0_dataflow_b;
	reg mesh_0_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_14_io_in_control_0_shift_b;
	reg mesh_1_14_io_in_control_0_dataflow_b;
	reg mesh_1_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_14_io_in_control_0_shift_b;
	reg mesh_2_14_io_in_control_0_dataflow_b;
	reg mesh_2_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_14_io_in_control_0_shift_b;
	reg mesh_3_14_io_in_control_0_dataflow_b;
	reg mesh_3_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_14_io_in_control_0_shift_b;
	reg mesh_4_14_io_in_control_0_dataflow_b;
	reg mesh_4_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_14_io_in_control_0_shift_b;
	reg mesh_5_14_io_in_control_0_dataflow_b;
	reg mesh_5_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_14_io_in_control_0_shift_b;
	reg mesh_6_14_io_in_control_0_dataflow_b;
	reg mesh_6_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_14_io_in_control_0_shift_b;
	reg mesh_7_14_io_in_control_0_dataflow_b;
	reg mesh_7_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_14_io_in_control_0_shift_b;
	reg mesh_8_14_io_in_control_0_dataflow_b;
	reg mesh_8_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_14_io_in_control_0_shift_b;
	reg mesh_9_14_io_in_control_0_dataflow_b;
	reg mesh_9_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_14_io_in_control_0_shift_b;
	reg mesh_10_14_io_in_control_0_dataflow_b;
	reg mesh_10_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_14_io_in_control_0_shift_b;
	reg mesh_11_14_io_in_control_0_dataflow_b;
	reg mesh_11_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_14_io_in_control_0_shift_b;
	reg mesh_12_14_io_in_control_0_dataflow_b;
	reg mesh_12_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_14_io_in_control_0_shift_b;
	reg mesh_13_14_io_in_control_0_dataflow_b;
	reg mesh_13_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_14_io_in_control_0_shift_b;
	reg mesh_14_14_io_in_control_0_dataflow_b;
	reg mesh_14_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_14_io_in_control_0_shift_b;
	reg mesh_15_14_io_in_control_0_dataflow_b;
	reg mesh_15_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_15_io_in_control_0_shift_b;
	reg mesh_0_15_io_in_control_0_dataflow_b;
	reg mesh_0_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_15_io_in_control_0_shift_b;
	reg mesh_1_15_io_in_control_0_dataflow_b;
	reg mesh_1_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_15_io_in_control_0_shift_b;
	reg mesh_2_15_io_in_control_0_dataflow_b;
	reg mesh_2_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_15_io_in_control_0_shift_b;
	reg mesh_3_15_io_in_control_0_dataflow_b;
	reg mesh_3_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_15_io_in_control_0_shift_b;
	reg mesh_4_15_io_in_control_0_dataflow_b;
	reg mesh_4_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_15_io_in_control_0_shift_b;
	reg mesh_5_15_io_in_control_0_dataflow_b;
	reg mesh_5_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_15_io_in_control_0_shift_b;
	reg mesh_6_15_io_in_control_0_dataflow_b;
	reg mesh_6_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_15_io_in_control_0_shift_b;
	reg mesh_7_15_io_in_control_0_dataflow_b;
	reg mesh_7_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_15_io_in_control_0_shift_b;
	reg mesh_8_15_io_in_control_0_dataflow_b;
	reg mesh_8_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_15_io_in_control_0_shift_b;
	reg mesh_9_15_io_in_control_0_dataflow_b;
	reg mesh_9_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_15_io_in_control_0_shift_b;
	reg mesh_10_15_io_in_control_0_dataflow_b;
	reg mesh_10_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_15_io_in_control_0_shift_b;
	reg mesh_11_15_io_in_control_0_dataflow_b;
	reg mesh_11_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_15_io_in_control_0_shift_b;
	reg mesh_12_15_io_in_control_0_dataflow_b;
	reg mesh_12_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_15_io_in_control_0_shift_b;
	reg mesh_13_15_io_in_control_0_dataflow_b;
	reg mesh_13_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_15_io_in_control_0_shift_b;
	reg mesh_14_15_io_in_control_0_dataflow_b;
	reg mesh_14_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_15_io_in_control_0_shift_b;
	reg mesh_15_15_io_in_control_0_dataflow_b;
	reg mesh_15_15_io_in_control_0_propagate_b;
	reg r_256_0;
	reg r_257_0;
	reg r_258_0;
	reg r_259_0;
	reg r_260_0;
	reg r_261_0;
	reg r_262_0;
	reg r_263_0;
	reg r_264_0;
	reg r_265_0;
	reg r_266_0;
	reg r_267_0;
	reg r_268_0;
	reg r_269_0;
	reg r_270_0;
	reg r_271_0;
	reg r_272_0;
	reg r_273_0;
	reg r_274_0;
	reg r_275_0;
	reg r_276_0;
	reg r_277_0;
	reg r_278_0;
	reg r_279_0;
	reg r_280_0;
	reg r_281_0;
	reg r_282_0;
	reg r_283_0;
	reg r_284_0;
	reg r_285_0;
	reg r_286_0;
	reg r_287_0;
	reg r_288_0;
	reg r_289_0;
	reg r_290_0;
	reg r_291_0;
	reg r_292_0;
	reg r_293_0;
	reg r_294_0;
	reg r_295_0;
	reg r_296_0;
	reg r_297_0;
	reg r_298_0;
	reg r_299_0;
	reg r_300_0;
	reg r_301_0;
	reg r_302_0;
	reg r_303_0;
	reg r_304_0;
	reg r_305_0;
	reg r_306_0;
	reg r_307_0;
	reg r_308_0;
	reg r_309_0;
	reg r_310_0;
	reg r_311_0;
	reg r_312_0;
	reg r_313_0;
	reg r_314_0;
	reg r_315_0;
	reg r_316_0;
	reg r_317_0;
	reg r_318_0;
	reg r_319_0;
	reg r_320_0;
	reg r_321_0;
	reg r_322_0;
	reg r_323_0;
	reg r_324_0;
	reg r_325_0;
	reg r_326_0;
	reg r_327_0;
	reg r_328_0;
	reg r_329_0;
	reg r_330_0;
	reg r_331_0;
	reg r_332_0;
	reg r_333_0;
	reg r_334_0;
	reg r_335_0;
	reg r_336_0;
	reg r_337_0;
	reg r_338_0;
	reg r_339_0;
	reg r_340_0;
	reg r_341_0;
	reg r_342_0;
	reg r_343_0;
	reg r_344_0;
	reg r_345_0;
	reg r_346_0;
	reg r_347_0;
	reg r_348_0;
	reg r_349_0;
	reg r_350_0;
	reg r_351_0;
	reg r_352_0;
	reg r_353_0;
	reg r_354_0;
	reg r_355_0;
	reg r_356_0;
	reg r_357_0;
	reg r_358_0;
	reg r_359_0;
	reg r_360_0;
	reg r_361_0;
	reg r_362_0;
	reg r_363_0;
	reg r_364_0;
	reg r_365_0;
	reg r_366_0;
	reg r_367_0;
	reg r_368_0;
	reg r_369_0;
	reg r_370_0;
	reg r_371_0;
	reg r_372_0;
	reg r_373_0;
	reg r_374_0;
	reg r_375_0;
	reg r_376_0;
	reg r_377_0;
	reg r_378_0;
	reg r_379_0;
	reg r_380_0;
	reg r_381_0;
	reg r_382_0;
	reg r_383_0;
	reg r_384_0;
	reg r_385_0;
	reg r_386_0;
	reg r_387_0;
	reg r_388_0;
	reg r_389_0;
	reg r_390_0;
	reg r_391_0;
	reg r_392_0;
	reg r_393_0;
	reg r_394_0;
	reg r_395_0;
	reg r_396_0;
	reg r_397_0;
	reg r_398_0;
	reg r_399_0;
	reg r_400_0;
	reg r_401_0;
	reg r_402_0;
	reg r_403_0;
	reg r_404_0;
	reg r_405_0;
	reg r_406_0;
	reg r_407_0;
	reg r_408_0;
	reg r_409_0;
	reg r_410_0;
	reg r_411_0;
	reg r_412_0;
	reg r_413_0;
	reg r_414_0;
	reg r_415_0;
	reg r_416_0;
	reg r_417_0;
	reg r_418_0;
	reg r_419_0;
	reg r_420_0;
	reg r_421_0;
	reg r_422_0;
	reg r_423_0;
	reg r_424_0;
	reg r_425_0;
	reg r_426_0;
	reg r_427_0;
	reg r_428_0;
	reg r_429_0;
	reg r_430_0;
	reg r_431_0;
	reg r_432_0;
	reg r_433_0;
	reg r_434_0;
	reg r_435_0;
	reg r_436_0;
	reg r_437_0;
	reg r_438_0;
	reg r_439_0;
	reg r_440_0;
	reg r_441_0;
	reg r_442_0;
	reg r_443_0;
	reg r_444_0;
	reg r_445_0;
	reg r_446_0;
	reg r_447_0;
	reg r_448_0;
	reg r_449_0;
	reg r_450_0;
	reg r_451_0;
	reg r_452_0;
	reg r_453_0;
	reg r_454_0;
	reg r_455_0;
	reg r_456_0;
	reg r_457_0;
	reg r_458_0;
	reg r_459_0;
	reg r_460_0;
	reg r_461_0;
	reg r_462_0;
	reg r_463_0;
	reg r_464_0;
	reg r_465_0;
	reg r_466_0;
	reg r_467_0;
	reg r_468_0;
	reg r_469_0;
	reg r_470_0;
	reg r_471_0;
	reg r_472_0;
	reg r_473_0;
	reg r_474_0;
	reg r_475_0;
	reg r_476_0;
	reg r_477_0;
	reg r_478_0;
	reg r_479_0;
	reg r_480_0;
	reg r_481_0;
	reg r_482_0;
	reg r_483_0;
	reg r_484_0;
	reg r_485_0;
	reg r_486_0;
	reg r_487_0;
	reg r_488_0;
	reg r_489_0;
	reg r_490_0;
	reg r_491_0;
	reg r_492_0;
	reg r_493_0;
	reg r_494_0;
	reg r_495_0;
	reg r_496_0;
	reg r_497_0;
	reg r_498_0;
	reg r_499_0;
	reg r_500_0;
	reg r_501_0;
	reg r_502_0;
	reg r_503_0;
	reg r_504_0;
	reg r_505_0;
	reg r_506_0;
	reg r_507_0;
	reg r_508_0;
	reg r_509_0;
	reg r_510_0;
	reg r_511_0;
	reg [2:0] r_512_0;
	reg [2:0] r_513_0;
	reg [2:0] r_514_0;
	reg [2:0] r_515_0;
	reg [2:0] r_516_0;
	reg [2:0] r_517_0;
	reg [2:0] r_518_0;
	reg [2:0] r_519_0;
	reg [2:0] r_520_0;
	reg [2:0] r_521_0;
	reg [2:0] r_522_0;
	reg [2:0] r_523_0;
	reg [2:0] r_524_0;
	reg [2:0] r_525_0;
	reg [2:0] r_526_0;
	reg [2:0] r_527_0;
	reg [2:0] r_528_0;
	reg [2:0] r_529_0;
	reg [2:0] r_530_0;
	reg [2:0] r_531_0;
	reg [2:0] r_532_0;
	reg [2:0] r_533_0;
	reg [2:0] r_534_0;
	reg [2:0] r_535_0;
	reg [2:0] r_536_0;
	reg [2:0] r_537_0;
	reg [2:0] r_538_0;
	reg [2:0] r_539_0;
	reg [2:0] r_540_0;
	reg [2:0] r_541_0;
	reg [2:0] r_542_0;
	reg [2:0] r_543_0;
	reg [2:0] r_544_0;
	reg [2:0] r_545_0;
	reg [2:0] r_546_0;
	reg [2:0] r_547_0;
	reg [2:0] r_548_0;
	reg [2:0] r_549_0;
	reg [2:0] r_550_0;
	reg [2:0] r_551_0;
	reg [2:0] r_552_0;
	reg [2:0] r_553_0;
	reg [2:0] r_554_0;
	reg [2:0] r_555_0;
	reg [2:0] r_556_0;
	reg [2:0] r_557_0;
	reg [2:0] r_558_0;
	reg [2:0] r_559_0;
	reg [2:0] r_560_0;
	reg [2:0] r_561_0;
	reg [2:0] r_562_0;
	reg [2:0] r_563_0;
	reg [2:0] r_564_0;
	reg [2:0] r_565_0;
	reg [2:0] r_566_0;
	reg [2:0] r_567_0;
	reg [2:0] r_568_0;
	reg [2:0] r_569_0;
	reg [2:0] r_570_0;
	reg [2:0] r_571_0;
	reg [2:0] r_572_0;
	reg [2:0] r_573_0;
	reg [2:0] r_574_0;
	reg [2:0] r_575_0;
	reg [2:0] r_576_0;
	reg [2:0] r_577_0;
	reg [2:0] r_578_0;
	reg [2:0] r_579_0;
	reg [2:0] r_580_0;
	reg [2:0] r_581_0;
	reg [2:0] r_582_0;
	reg [2:0] r_583_0;
	reg [2:0] r_584_0;
	reg [2:0] r_585_0;
	reg [2:0] r_586_0;
	reg [2:0] r_587_0;
	reg [2:0] r_588_0;
	reg [2:0] r_589_0;
	reg [2:0] r_590_0;
	reg [2:0] r_591_0;
	reg [2:0] r_592_0;
	reg [2:0] r_593_0;
	reg [2:0] r_594_0;
	reg [2:0] r_595_0;
	reg [2:0] r_596_0;
	reg [2:0] r_597_0;
	reg [2:0] r_598_0;
	reg [2:0] r_599_0;
	reg [2:0] r_600_0;
	reg [2:0] r_601_0;
	reg [2:0] r_602_0;
	reg [2:0] r_603_0;
	reg [2:0] r_604_0;
	reg [2:0] r_605_0;
	reg [2:0] r_606_0;
	reg [2:0] r_607_0;
	reg [2:0] r_608_0;
	reg [2:0] r_609_0;
	reg [2:0] r_610_0;
	reg [2:0] r_611_0;
	reg [2:0] r_612_0;
	reg [2:0] r_613_0;
	reg [2:0] r_614_0;
	reg [2:0] r_615_0;
	reg [2:0] r_616_0;
	reg [2:0] r_617_0;
	reg [2:0] r_618_0;
	reg [2:0] r_619_0;
	reg [2:0] r_620_0;
	reg [2:0] r_621_0;
	reg [2:0] r_622_0;
	reg [2:0] r_623_0;
	reg [2:0] r_624_0;
	reg [2:0] r_625_0;
	reg [2:0] r_626_0;
	reg [2:0] r_627_0;
	reg [2:0] r_628_0;
	reg [2:0] r_629_0;
	reg [2:0] r_630_0;
	reg [2:0] r_631_0;
	reg [2:0] r_632_0;
	reg [2:0] r_633_0;
	reg [2:0] r_634_0;
	reg [2:0] r_635_0;
	reg [2:0] r_636_0;
	reg [2:0] r_637_0;
	reg [2:0] r_638_0;
	reg [2:0] r_639_0;
	reg [2:0] r_640_0;
	reg [2:0] r_641_0;
	reg [2:0] r_642_0;
	reg [2:0] r_643_0;
	reg [2:0] r_644_0;
	reg [2:0] r_645_0;
	reg [2:0] r_646_0;
	reg [2:0] r_647_0;
	reg [2:0] r_648_0;
	reg [2:0] r_649_0;
	reg [2:0] r_650_0;
	reg [2:0] r_651_0;
	reg [2:0] r_652_0;
	reg [2:0] r_653_0;
	reg [2:0] r_654_0;
	reg [2:0] r_655_0;
	reg [2:0] r_656_0;
	reg [2:0] r_657_0;
	reg [2:0] r_658_0;
	reg [2:0] r_659_0;
	reg [2:0] r_660_0;
	reg [2:0] r_661_0;
	reg [2:0] r_662_0;
	reg [2:0] r_663_0;
	reg [2:0] r_664_0;
	reg [2:0] r_665_0;
	reg [2:0] r_666_0;
	reg [2:0] r_667_0;
	reg [2:0] r_668_0;
	reg [2:0] r_669_0;
	reg [2:0] r_670_0;
	reg [2:0] r_671_0;
	reg [2:0] r_672_0;
	reg [2:0] r_673_0;
	reg [2:0] r_674_0;
	reg [2:0] r_675_0;
	reg [2:0] r_676_0;
	reg [2:0] r_677_0;
	reg [2:0] r_678_0;
	reg [2:0] r_679_0;
	reg [2:0] r_680_0;
	reg [2:0] r_681_0;
	reg [2:0] r_682_0;
	reg [2:0] r_683_0;
	reg [2:0] r_684_0;
	reg [2:0] r_685_0;
	reg [2:0] r_686_0;
	reg [2:0] r_687_0;
	reg [2:0] r_688_0;
	reg [2:0] r_689_0;
	reg [2:0] r_690_0;
	reg [2:0] r_691_0;
	reg [2:0] r_692_0;
	reg [2:0] r_693_0;
	reg [2:0] r_694_0;
	reg [2:0] r_695_0;
	reg [2:0] r_696_0;
	reg [2:0] r_697_0;
	reg [2:0] r_698_0;
	reg [2:0] r_699_0;
	reg [2:0] r_700_0;
	reg [2:0] r_701_0;
	reg [2:0] r_702_0;
	reg [2:0] r_703_0;
	reg [2:0] r_704_0;
	reg [2:0] r_705_0;
	reg [2:0] r_706_0;
	reg [2:0] r_707_0;
	reg [2:0] r_708_0;
	reg [2:0] r_709_0;
	reg [2:0] r_710_0;
	reg [2:0] r_711_0;
	reg [2:0] r_712_0;
	reg [2:0] r_713_0;
	reg [2:0] r_714_0;
	reg [2:0] r_715_0;
	reg [2:0] r_716_0;
	reg [2:0] r_717_0;
	reg [2:0] r_718_0;
	reg [2:0] r_719_0;
	reg [2:0] r_720_0;
	reg [2:0] r_721_0;
	reg [2:0] r_722_0;
	reg [2:0] r_723_0;
	reg [2:0] r_724_0;
	reg [2:0] r_725_0;
	reg [2:0] r_726_0;
	reg [2:0] r_727_0;
	reg [2:0] r_728_0;
	reg [2:0] r_729_0;
	reg [2:0] r_730_0;
	reg [2:0] r_731_0;
	reg [2:0] r_732_0;
	reg [2:0] r_733_0;
	reg [2:0] r_734_0;
	reg [2:0] r_735_0;
	reg [2:0] r_736_0;
	reg [2:0] r_737_0;
	reg [2:0] r_738_0;
	reg [2:0] r_739_0;
	reg [2:0] r_740_0;
	reg [2:0] r_741_0;
	reg [2:0] r_742_0;
	reg [2:0] r_743_0;
	reg [2:0] r_744_0;
	reg [2:0] r_745_0;
	reg [2:0] r_746_0;
	reg [2:0] r_747_0;
	reg [2:0] r_748_0;
	reg [2:0] r_749_0;
	reg [2:0] r_750_0;
	reg [2:0] r_751_0;
	reg [2:0] r_752_0;
	reg [2:0] r_753_0;
	reg [2:0] r_754_0;
	reg [2:0] r_755_0;
	reg [2:0] r_756_0;
	reg [2:0] r_757_0;
	reg [2:0] r_758_0;
	reg [2:0] r_759_0;
	reg [2:0] r_760_0;
	reg [2:0] r_761_0;
	reg [2:0] r_762_0;
	reg [2:0] r_763_0;
	reg [2:0] r_764_0;
	reg [2:0] r_765_0;
	reg [2:0] r_766_0;
	reg [2:0] r_767_0;
	reg r_768_0;
	reg r_769_0;
	reg r_770_0;
	reg r_771_0;
	reg r_772_0;
	reg r_773_0;
	reg r_774_0;
	reg r_775_0;
	reg r_776_0;
	reg r_777_0;
	reg r_778_0;
	reg r_779_0;
	reg r_780_0;
	reg r_781_0;
	reg r_782_0;
	reg r_783_0;
	reg r_784_0;
	reg r_785_0;
	reg r_786_0;
	reg r_787_0;
	reg r_788_0;
	reg r_789_0;
	reg r_790_0;
	reg r_791_0;
	reg r_792_0;
	reg r_793_0;
	reg r_794_0;
	reg r_795_0;
	reg r_796_0;
	reg r_797_0;
	reg r_798_0;
	reg r_799_0;
	reg r_800_0;
	reg r_801_0;
	reg r_802_0;
	reg r_803_0;
	reg r_804_0;
	reg r_805_0;
	reg r_806_0;
	reg r_807_0;
	reg r_808_0;
	reg r_809_0;
	reg r_810_0;
	reg r_811_0;
	reg r_812_0;
	reg r_813_0;
	reg r_814_0;
	reg r_815_0;
	reg r_816_0;
	reg r_817_0;
	reg r_818_0;
	reg r_819_0;
	reg r_820_0;
	reg r_821_0;
	reg r_822_0;
	reg r_823_0;
	reg r_824_0;
	reg r_825_0;
	reg r_826_0;
	reg r_827_0;
	reg r_828_0;
	reg r_829_0;
	reg r_830_0;
	reg r_831_0;
	reg r_832_0;
	reg r_833_0;
	reg r_834_0;
	reg r_835_0;
	reg r_836_0;
	reg r_837_0;
	reg r_838_0;
	reg r_839_0;
	reg r_840_0;
	reg r_841_0;
	reg r_842_0;
	reg r_843_0;
	reg r_844_0;
	reg r_845_0;
	reg r_846_0;
	reg r_847_0;
	reg r_848_0;
	reg r_849_0;
	reg r_850_0;
	reg r_851_0;
	reg r_852_0;
	reg r_853_0;
	reg r_854_0;
	reg r_855_0;
	reg r_856_0;
	reg r_857_0;
	reg r_858_0;
	reg r_859_0;
	reg r_860_0;
	reg r_861_0;
	reg r_862_0;
	reg r_863_0;
	reg r_864_0;
	reg r_865_0;
	reg r_866_0;
	reg r_867_0;
	reg r_868_0;
	reg r_869_0;
	reg r_870_0;
	reg r_871_0;
	reg r_872_0;
	reg r_873_0;
	reg r_874_0;
	reg r_875_0;
	reg r_876_0;
	reg r_877_0;
	reg r_878_0;
	reg r_879_0;
	reg r_880_0;
	reg r_881_0;
	reg r_882_0;
	reg r_883_0;
	reg r_884_0;
	reg r_885_0;
	reg r_886_0;
	reg r_887_0;
	reg r_888_0;
	reg r_889_0;
	reg r_890_0;
	reg r_891_0;
	reg r_892_0;
	reg r_893_0;
	reg r_894_0;
	reg r_895_0;
	reg r_896_0;
	reg r_897_0;
	reg r_898_0;
	reg r_899_0;
	reg r_900_0;
	reg r_901_0;
	reg r_902_0;
	reg r_903_0;
	reg r_904_0;
	reg r_905_0;
	reg r_906_0;
	reg r_907_0;
	reg r_908_0;
	reg r_909_0;
	reg r_910_0;
	reg r_911_0;
	reg r_912_0;
	reg r_913_0;
	reg r_914_0;
	reg r_915_0;
	reg r_916_0;
	reg r_917_0;
	reg r_918_0;
	reg r_919_0;
	reg r_920_0;
	reg r_921_0;
	reg r_922_0;
	reg r_923_0;
	reg r_924_0;
	reg r_925_0;
	reg r_926_0;
	reg r_927_0;
	reg r_928_0;
	reg r_929_0;
	reg r_930_0;
	reg r_931_0;
	reg r_932_0;
	reg r_933_0;
	reg r_934_0;
	reg r_935_0;
	reg r_936_0;
	reg r_937_0;
	reg r_938_0;
	reg r_939_0;
	reg r_940_0;
	reg r_941_0;
	reg r_942_0;
	reg r_943_0;
	reg r_944_0;
	reg r_945_0;
	reg r_946_0;
	reg r_947_0;
	reg r_948_0;
	reg r_949_0;
	reg r_950_0;
	reg r_951_0;
	reg r_952_0;
	reg r_953_0;
	reg r_954_0;
	reg r_955_0;
	reg r_956_0;
	reg r_957_0;
	reg r_958_0;
	reg r_959_0;
	reg r_960_0;
	reg r_961_0;
	reg r_962_0;
	reg r_963_0;
	reg r_964_0;
	reg r_965_0;
	reg r_966_0;
	reg r_967_0;
	reg r_968_0;
	reg r_969_0;
	reg r_970_0;
	reg r_971_0;
	reg r_972_0;
	reg r_973_0;
	reg r_974_0;
	reg r_975_0;
	reg r_976_0;
	reg r_977_0;
	reg r_978_0;
	reg r_979_0;
	reg r_980_0;
	reg r_981_0;
	reg r_982_0;
	reg r_983_0;
	reg r_984_0;
	reg r_985_0;
	reg r_986_0;
	reg r_987_0;
	reg r_988_0;
	reg r_989_0;
	reg r_990_0;
	reg r_991_0;
	reg r_992_0;
	reg r_993_0;
	reg r_994_0;
	reg r_995_0;
	reg r_996_0;
	reg r_997_0;
	reg r_998_0;
	reg r_999_0;
	reg r_1000_0;
	reg r_1001_0;
	reg r_1002_0;
	reg r_1003_0;
	reg r_1004_0;
	reg r_1005_0;
	reg r_1006_0;
	reg r_1007_0;
	reg r_1008_0;
	reg r_1009_0;
	reg r_1010_0;
	reg r_1011_0;
	reg r_1012_0;
	reg r_1013_0;
	reg r_1014_0;
	reg r_1015_0;
	reg r_1016_0;
	reg r_1017_0;
	reg r_1018_0;
	reg r_1019_0;
	reg r_1020_0;
	reg r_1021_0;
	reg r_1022_0;
	reg r_1023_0;
	reg [31:0] r_1024_0;
	reg [31:0] r_1025_0;
	reg r_1026_0;
	reg r_1027_0_dataflow;
	reg [2:0] r_1028_0;
	reg r_1029_0;
	reg [31:0] r_1030_0;
	reg [31:0] r_1031_0;
	reg [31:0] r_1036_0;
	reg [31:0] r_1037_0;
	reg [31:0] r_1042_0;
	reg [31:0] r_1043_0;
	reg [31:0] r_1048_0;
	reg [31:0] r_1049_0;
	reg [31:0] r_1054_0;
	reg [31:0] r_1055_0;
	reg [31:0] r_1060_0;
	reg [31:0] r_1061_0;
	reg [31:0] r_1066_0;
	reg [31:0] r_1067_0;
	reg [31:0] r_1072_0;
	reg [31:0] r_1073_0;
	reg [31:0] r_1078_0;
	reg [31:0] r_1079_0;
	reg [31:0] r_1084_0;
	reg [31:0] r_1085_0;
	reg [31:0] r_1090_0;
	reg [31:0] r_1091_0;
	reg [31:0] r_1096_0;
	reg [31:0] r_1097_0;
	reg [31:0] r_1102_0;
	reg [31:0] r_1103_0;
	reg [31:0] r_1108_0;
	reg [31:0] r_1109_0;
	reg [31:0] r_1114_0;
	reg [31:0] r_1115_0;
	always @(posedge clock) begin
		r_0 <=( io_in_a_0_0) ^ ((fiEnable && (17 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1_0 <=( _mesh_0_0_io_out_a_0) ^ ((fiEnable && (18 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_2_0 <=( _mesh_0_1_io_out_a_0) ^ ((fiEnable && (19 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_3_0 <=( _mesh_0_2_io_out_a_0) ^ ((fiEnable && (20 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4_0 <=( _mesh_0_3_io_out_a_0) ^ ((fiEnable && (21 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_5_0 <=( _mesh_0_4_io_out_a_0) ^ ((fiEnable && (22 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_6_0 <=( _mesh_0_5_io_out_a_0) ^ ((fiEnable && (23 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_7_0 <=( _mesh_0_6_io_out_a_0) ^ ((fiEnable && (24 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_8_0 <=( _mesh_0_7_io_out_a_0) ^ ((fiEnable && (25 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_9_0 <=( _mesh_0_8_io_out_a_0) ^ ((fiEnable && (26 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_10_0 <=( _mesh_0_9_io_out_a_0) ^ ((fiEnable && (27 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_11_0 <=( _mesh_0_10_io_out_a_0) ^ ((fiEnable && (28 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_12_0 <=( _mesh_0_11_io_out_a_0) ^ ((fiEnable && (29 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_13_0 <=( _mesh_0_12_io_out_a_0) ^ ((fiEnable && (30 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_14_0 <=( _mesh_0_13_io_out_a_0) ^ ((fiEnable && (31 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_15_0 <=( _mesh_0_14_io_out_a_0) ^ ((fiEnable && (32 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_16_0 <=( io_in_a_1_0) ^ ((fiEnable && (33 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_17_0 <=( _mesh_1_0_io_out_a_0) ^ ((fiEnable && (34 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_18_0 <=( _mesh_1_1_io_out_a_0) ^ ((fiEnable && (35 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_19_0 <=( _mesh_1_2_io_out_a_0) ^ ((fiEnable && (36 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_20_0 <=( _mesh_1_3_io_out_a_0) ^ ((fiEnable && (37 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_21_0 <=( _mesh_1_4_io_out_a_0) ^ ((fiEnable && (38 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_22_0 <=( _mesh_1_5_io_out_a_0) ^ ((fiEnable && (39 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_23_0 <=( _mesh_1_6_io_out_a_0) ^ ((fiEnable && (40 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_24_0 <=( _mesh_1_7_io_out_a_0) ^ ((fiEnable && (41 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_25_0 <=( _mesh_1_8_io_out_a_0) ^ ((fiEnable && (42 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_26_0 <=( _mesh_1_9_io_out_a_0) ^ ((fiEnable && (43 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_27_0 <=( _mesh_1_10_io_out_a_0) ^ ((fiEnable && (44 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_28_0 <=( _mesh_1_11_io_out_a_0) ^ ((fiEnable && (45 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_29_0 <=( _mesh_1_12_io_out_a_0) ^ ((fiEnable && (46 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_30_0 <=( _mesh_1_13_io_out_a_0) ^ ((fiEnable && (47 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_31_0 <=( _mesh_1_14_io_out_a_0) ^ ((fiEnable && (48 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_32_0 <=( io_in_a_2_0) ^ ((fiEnable && (49 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_33_0 <=( _mesh_2_0_io_out_a_0) ^ ((fiEnable && (50 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_34_0 <=( _mesh_2_1_io_out_a_0) ^ ((fiEnable && (51 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_35_0 <=( _mesh_2_2_io_out_a_0) ^ ((fiEnable && (52 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_36_0 <=( _mesh_2_3_io_out_a_0) ^ ((fiEnable && (53 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_37_0 <=( _mesh_2_4_io_out_a_0) ^ ((fiEnable && (54 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_38_0 <=( _mesh_2_5_io_out_a_0) ^ ((fiEnable && (55 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_39_0 <=( _mesh_2_6_io_out_a_0) ^ ((fiEnable && (56 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_40_0 <=( _mesh_2_7_io_out_a_0) ^ ((fiEnable && (57 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_41_0 <=( _mesh_2_8_io_out_a_0) ^ ((fiEnable && (58 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_42_0 <=( _mesh_2_9_io_out_a_0) ^ ((fiEnable && (59 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_43_0 <=( _mesh_2_10_io_out_a_0) ^ ((fiEnable && (60 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_44_0 <=( _mesh_2_11_io_out_a_0) ^ ((fiEnable && (61 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_45_0 <=( _mesh_2_12_io_out_a_0) ^ ((fiEnable && (62 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_46_0 <=( _mesh_2_13_io_out_a_0) ^ ((fiEnable && (63 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_47_0 <=( _mesh_2_14_io_out_a_0) ^ ((fiEnable && (64 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_48_0 <=( io_in_a_3_0) ^ ((fiEnable && (65 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_49_0 <=( _mesh_3_0_io_out_a_0) ^ ((fiEnable && (66 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_50_0 <=( _mesh_3_1_io_out_a_0) ^ ((fiEnable && (67 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_51_0 <=( _mesh_3_2_io_out_a_0) ^ ((fiEnable && (68 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_52_0 <=( _mesh_3_3_io_out_a_0) ^ ((fiEnable && (69 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_53_0 <=( _mesh_3_4_io_out_a_0) ^ ((fiEnable && (70 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_54_0 <=( _mesh_3_5_io_out_a_0) ^ ((fiEnable && (71 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_55_0 <=( _mesh_3_6_io_out_a_0) ^ ((fiEnable && (72 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_56_0 <=( _mesh_3_7_io_out_a_0) ^ ((fiEnable && (73 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_57_0 <=( _mesh_3_8_io_out_a_0) ^ ((fiEnable && (74 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_58_0 <=( _mesh_3_9_io_out_a_0) ^ ((fiEnable && (75 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_59_0 <=( _mesh_3_10_io_out_a_0) ^ ((fiEnable && (76 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_60_0 <=( _mesh_3_11_io_out_a_0) ^ ((fiEnable && (77 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_61_0 <=( _mesh_3_12_io_out_a_0) ^ ((fiEnable && (78 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_62_0 <=( _mesh_3_13_io_out_a_0) ^ ((fiEnable && (79 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_63_0 <=( _mesh_3_14_io_out_a_0) ^ ((fiEnable && (80 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_64_0 <=( io_in_a_4_0) ^ ((fiEnable && (81 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_65_0 <=( _mesh_4_0_io_out_a_0) ^ ((fiEnable && (82 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_66_0 <=( _mesh_4_1_io_out_a_0) ^ ((fiEnable && (83 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_67_0 <=( _mesh_4_2_io_out_a_0) ^ ((fiEnable && (84 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_68_0 <=( _mesh_4_3_io_out_a_0) ^ ((fiEnable && (85 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_69_0 <=( _mesh_4_4_io_out_a_0) ^ ((fiEnable && (86 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_70_0 <=( _mesh_4_5_io_out_a_0) ^ ((fiEnable && (87 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_71_0 <=( _mesh_4_6_io_out_a_0) ^ ((fiEnable && (88 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_72_0 <=( _mesh_4_7_io_out_a_0) ^ ((fiEnable && (89 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_73_0 <=( _mesh_4_8_io_out_a_0) ^ ((fiEnable && (90 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_74_0 <=( _mesh_4_9_io_out_a_0) ^ ((fiEnable && (91 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_75_0 <=( _mesh_4_10_io_out_a_0) ^ ((fiEnable && (92 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_76_0 <=( _mesh_4_11_io_out_a_0) ^ ((fiEnable && (93 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_77_0 <=( _mesh_4_12_io_out_a_0) ^ ((fiEnable && (94 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_78_0 <=( _mesh_4_13_io_out_a_0) ^ ((fiEnable && (95 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_79_0 <=( _mesh_4_14_io_out_a_0) ^ ((fiEnable && (96 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_80_0 <=( io_in_a_5_0) ^ ((fiEnable && (97 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_81_0 <=( _mesh_5_0_io_out_a_0) ^ ((fiEnable && (98 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_82_0 <=( _mesh_5_1_io_out_a_0) ^ ((fiEnable && (99 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_83_0 <=( _mesh_5_2_io_out_a_0) ^ ((fiEnable && (100 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_84_0 <=( _mesh_5_3_io_out_a_0) ^ ((fiEnable && (101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_85_0 <=( _mesh_5_4_io_out_a_0) ^ ((fiEnable && (102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_86_0 <=( _mesh_5_5_io_out_a_0) ^ ((fiEnable && (103 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_87_0 <=( _mesh_5_6_io_out_a_0) ^ ((fiEnable && (104 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_88_0 <=( _mesh_5_7_io_out_a_0) ^ ((fiEnable && (105 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_89_0 <=( _mesh_5_8_io_out_a_0) ^ ((fiEnable && (106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_90_0 <=( _mesh_5_9_io_out_a_0) ^ ((fiEnable && (107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_91_0 <=( _mesh_5_10_io_out_a_0) ^ ((fiEnable && (108 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_92_0 <=( _mesh_5_11_io_out_a_0) ^ ((fiEnable && (109 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_93_0 <=( _mesh_5_12_io_out_a_0) ^ ((fiEnable && (110 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_94_0 <=( _mesh_5_13_io_out_a_0) ^ ((fiEnable && (111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_95_0 <=( _mesh_5_14_io_out_a_0) ^ ((fiEnable && (112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_96_0 <=( io_in_a_6_0) ^ ((fiEnable && (113 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_97_0 <=( _mesh_6_0_io_out_a_0) ^ ((fiEnable && (114 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_98_0 <=( _mesh_6_1_io_out_a_0) ^ ((fiEnable && (115 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_99_0 <=( _mesh_6_2_io_out_a_0) ^ ((fiEnable && (116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_100_0 <=( _mesh_6_3_io_out_a_0) ^ ((fiEnable && (117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_101_0 <=( _mesh_6_4_io_out_a_0) ^ ((fiEnable && (118 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_102_0 <=( _mesh_6_5_io_out_a_0) ^ ((fiEnable && (119 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_103_0 <=( _mesh_6_6_io_out_a_0) ^ ((fiEnable && (120 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_104_0 <=( _mesh_6_7_io_out_a_0) ^ ((fiEnable && (121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_105_0 <=( _mesh_6_8_io_out_a_0) ^ ((fiEnable && (122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_106_0 <=( _mesh_6_9_io_out_a_0) ^ ((fiEnable && (123 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_107_0 <=( _mesh_6_10_io_out_a_0) ^ ((fiEnable && (124 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_108_0 <=( _mesh_6_11_io_out_a_0) ^ ((fiEnable && (125 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_109_0 <=( _mesh_6_12_io_out_a_0) ^ ((fiEnable && (126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_110_0 <=( _mesh_6_13_io_out_a_0) ^ ((fiEnable && (127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_111_0 <=( _mesh_6_14_io_out_a_0) ^ ((fiEnable && (128 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_112_0 <=( io_in_a_7_0) ^ ((fiEnable && (129 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_113_0 <=( _mesh_7_0_io_out_a_0) ^ ((fiEnable && (130 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_114_0 <=( _mesh_7_1_io_out_a_0) ^ ((fiEnable && (131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_115_0 <=( _mesh_7_2_io_out_a_0) ^ ((fiEnable && (132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_116_0 <=( _mesh_7_3_io_out_a_0) ^ ((fiEnable && (133 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_117_0 <=( _mesh_7_4_io_out_a_0) ^ ((fiEnable && (134 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_118_0 <=( _mesh_7_5_io_out_a_0) ^ ((fiEnable && (135 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_119_0 <=( _mesh_7_6_io_out_a_0) ^ ((fiEnable && (136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_120_0 <=( _mesh_7_7_io_out_a_0) ^ ((fiEnable && (137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_121_0 <=( _mesh_7_8_io_out_a_0) ^ ((fiEnable && (138 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_122_0 <=( _mesh_7_9_io_out_a_0) ^ ((fiEnable && (139 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_123_0 <=( _mesh_7_10_io_out_a_0) ^ ((fiEnable && (140 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_124_0 <=( _mesh_7_11_io_out_a_0) ^ ((fiEnable && (141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_125_0 <=( _mesh_7_12_io_out_a_0) ^ ((fiEnable && (142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_126_0 <=( _mesh_7_13_io_out_a_0) ^ ((fiEnable && (143 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_127_0 <=( _mesh_7_14_io_out_a_0) ^ ((fiEnable && (144 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_128_0 <=( io_in_a_8_0) ^ ((fiEnable && (145 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_129_0 <=( _mesh_8_0_io_out_a_0) ^ ((fiEnable && (146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_130_0 <=( _mesh_8_1_io_out_a_0) ^ ((fiEnable && (147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_131_0 <=( _mesh_8_2_io_out_a_0) ^ ((fiEnable && (148 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_132_0 <=( _mesh_8_3_io_out_a_0) ^ ((fiEnable && (149 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_133_0 <=( _mesh_8_4_io_out_a_0) ^ ((fiEnable && (150 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_134_0 <=( _mesh_8_5_io_out_a_0) ^ ((fiEnable && (151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_135_0 <=( _mesh_8_6_io_out_a_0) ^ ((fiEnable && (152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_136_0 <=( _mesh_8_7_io_out_a_0) ^ ((fiEnable && (153 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_137_0 <=( _mesh_8_8_io_out_a_0) ^ ((fiEnable && (154 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_138_0 <=( _mesh_8_9_io_out_a_0) ^ ((fiEnable && (155 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_139_0 <=( _mesh_8_10_io_out_a_0) ^ ((fiEnable && (156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_140_0 <=( _mesh_8_11_io_out_a_0) ^ ((fiEnable && (157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_141_0 <=( _mesh_8_12_io_out_a_0) ^ ((fiEnable && (158 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_142_0 <=( _mesh_8_13_io_out_a_0) ^ ((fiEnable && (159 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_143_0 <=( _mesh_8_14_io_out_a_0) ^ ((fiEnable && (160 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_144_0 <=( io_in_a_9_0) ^ ((fiEnable && (161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_145_0 <=( _mesh_9_0_io_out_a_0) ^ ((fiEnable && (162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_146_0 <=( _mesh_9_1_io_out_a_0) ^ ((fiEnable && (163 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_147_0 <=( _mesh_9_2_io_out_a_0) ^ ((fiEnable && (164 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_148_0 <=( _mesh_9_3_io_out_a_0) ^ ((fiEnable && (165 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_149_0 <=( _mesh_9_4_io_out_a_0) ^ ((fiEnable && (166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_150_0 <=( _mesh_9_5_io_out_a_0) ^ ((fiEnable && (167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_151_0 <=( _mesh_9_6_io_out_a_0) ^ ((fiEnable && (168 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_152_0 <=( _mesh_9_7_io_out_a_0) ^ ((fiEnable && (169 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_153_0 <=( _mesh_9_8_io_out_a_0) ^ ((fiEnable && (170 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_154_0 <=( _mesh_9_9_io_out_a_0) ^ ((fiEnable && (171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_155_0 <=( _mesh_9_10_io_out_a_0) ^ ((fiEnable && (172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_156_0 <=( _mesh_9_11_io_out_a_0) ^ ((fiEnable && (173 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_157_0 <=( _mesh_9_12_io_out_a_0) ^ ((fiEnable && (174 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_158_0 <=( _mesh_9_13_io_out_a_0) ^ ((fiEnable && (175 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_159_0 <=( _mesh_9_14_io_out_a_0) ^ ((fiEnable && (176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_160_0 <=( io_in_a_10_0) ^ ((fiEnable && (177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_161_0 <=( _mesh_10_0_io_out_a_0) ^ ((fiEnable && (178 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_162_0 <=( _mesh_10_1_io_out_a_0) ^ ((fiEnable && (179 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_163_0 <=( _mesh_10_2_io_out_a_0) ^ ((fiEnable && (180 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_164_0 <=( _mesh_10_3_io_out_a_0) ^ ((fiEnable && (181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_165_0 <=( _mesh_10_4_io_out_a_0) ^ ((fiEnable && (182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_166_0 <=( _mesh_10_5_io_out_a_0) ^ ((fiEnable && (183 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_167_0 <=( _mesh_10_6_io_out_a_0) ^ ((fiEnable && (184 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_168_0 <=( _mesh_10_7_io_out_a_0) ^ ((fiEnable && (185 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_169_0 <=( _mesh_10_8_io_out_a_0) ^ ((fiEnable && (186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_170_0 <=( _mesh_10_9_io_out_a_0) ^ ((fiEnable && (187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_171_0 <=( _mesh_10_10_io_out_a_0) ^ ((fiEnable && (188 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_172_0 <=( _mesh_10_11_io_out_a_0) ^ ((fiEnable && (189 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_173_0 <=( _mesh_10_12_io_out_a_0) ^ ((fiEnable && (190 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_174_0 <=( _mesh_10_13_io_out_a_0) ^ ((fiEnable && (191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_175_0 <=( _mesh_10_14_io_out_a_0) ^ ((fiEnable && (192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_176_0 <=( io_in_a_11_0) ^ ((fiEnable && (193 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_177_0 <=( _mesh_11_0_io_out_a_0) ^ ((fiEnable && (194 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_178_0 <=( _mesh_11_1_io_out_a_0) ^ ((fiEnable && (195 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_179_0 <=( _mesh_11_2_io_out_a_0) ^ ((fiEnable && (196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_180_0 <=( _mesh_11_3_io_out_a_0) ^ ((fiEnable && (197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_181_0 <=( _mesh_11_4_io_out_a_0) ^ ((fiEnable && (198 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_182_0 <=( _mesh_11_5_io_out_a_0) ^ ((fiEnable && (199 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_183_0 <=( _mesh_11_6_io_out_a_0) ^ ((fiEnable && (200 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_184_0 <=( _mesh_11_7_io_out_a_0) ^ ((fiEnable && (201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_185_0 <=( _mesh_11_8_io_out_a_0) ^ ((fiEnable && (202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_186_0 <=( _mesh_11_9_io_out_a_0) ^ ((fiEnable && (203 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_187_0 <=( _mesh_11_10_io_out_a_0) ^ ((fiEnable && (204 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_188_0 <=( _mesh_11_11_io_out_a_0) ^ ((fiEnable && (205 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_189_0 <=( _mesh_11_12_io_out_a_0) ^ ((fiEnable && (206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_190_0 <=( _mesh_11_13_io_out_a_0) ^ ((fiEnable && (207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_191_0 <=( _mesh_11_14_io_out_a_0) ^ ((fiEnable && (208 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_192_0 <=( io_in_a_12_0) ^ ((fiEnable && (209 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_193_0 <=( _mesh_12_0_io_out_a_0) ^ ((fiEnable && (210 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_194_0 <=( _mesh_12_1_io_out_a_0) ^ ((fiEnable && (211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_195_0 <=( _mesh_12_2_io_out_a_0) ^ ((fiEnable && (212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_196_0 <=( _mesh_12_3_io_out_a_0) ^ ((fiEnable && (213 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_197_0 <=( _mesh_12_4_io_out_a_0) ^ ((fiEnable && (214 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_198_0 <=( _mesh_12_5_io_out_a_0) ^ ((fiEnable && (215 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_199_0 <=( _mesh_12_6_io_out_a_0) ^ ((fiEnable && (216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_200_0 <=( _mesh_12_7_io_out_a_0) ^ ((fiEnable && (217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_201_0 <=( _mesh_12_8_io_out_a_0) ^ ((fiEnable && (218 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_202_0 <=( _mesh_12_9_io_out_a_0) ^ ((fiEnable && (219 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_203_0 <=( _mesh_12_10_io_out_a_0) ^ ((fiEnable && (220 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_204_0 <=( _mesh_12_11_io_out_a_0) ^ ((fiEnable && (221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_205_0 <=( _mesh_12_12_io_out_a_0) ^ ((fiEnable && (222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_206_0 <=( _mesh_12_13_io_out_a_0) ^ ((fiEnable && (223 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_207_0 <=( _mesh_12_14_io_out_a_0) ^ ((fiEnable && (224 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_208_0 <=( io_in_a_13_0) ^ ((fiEnable && (225 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_209_0 <=( _mesh_13_0_io_out_a_0) ^ ((fiEnable && (226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_210_0 <=( _mesh_13_1_io_out_a_0) ^ ((fiEnable && (227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_211_0 <=( _mesh_13_2_io_out_a_0) ^ ((fiEnable && (228 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_212_0 <=( _mesh_13_3_io_out_a_0) ^ ((fiEnable && (229 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_213_0 <=( _mesh_13_4_io_out_a_0) ^ ((fiEnable && (230 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_214_0 <=( _mesh_13_5_io_out_a_0) ^ ((fiEnable && (231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_215_0 <=( _mesh_13_6_io_out_a_0) ^ ((fiEnable && (232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_216_0 <=( _mesh_13_7_io_out_a_0) ^ ((fiEnable && (233 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_217_0 <=( _mesh_13_8_io_out_a_0) ^ ((fiEnable && (234 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_218_0 <=( _mesh_13_9_io_out_a_0) ^ ((fiEnable && (235 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_219_0 <=( _mesh_13_10_io_out_a_0) ^ ((fiEnable && (236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_220_0 <=( _mesh_13_11_io_out_a_0) ^ ((fiEnable && (237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_221_0 <=( _mesh_13_12_io_out_a_0) ^ ((fiEnable && (238 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_222_0 <=( _mesh_13_13_io_out_a_0) ^ ((fiEnable && (239 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_223_0 <=( _mesh_13_14_io_out_a_0) ^ ((fiEnable && (240 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_224_0 <=( io_in_a_14_0) ^ ((fiEnable && (241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_225_0 <=( _mesh_14_0_io_out_a_0) ^ ((fiEnable && (242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_226_0 <=( _mesh_14_1_io_out_a_0) ^ ((fiEnable && (243 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_227_0 <=( _mesh_14_2_io_out_a_0) ^ ((fiEnable && (244 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_228_0 <=( _mesh_14_3_io_out_a_0) ^ ((fiEnable && (245 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_229_0 <=( _mesh_14_4_io_out_a_0) ^ ((fiEnable && (246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_230_0 <=( _mesh_14_5_io_out_a_0) ^ ((fiEnable && (247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_231_0 <=( _mesh_14_6_io_out_a_0) ^ ((fiEnable && (248 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_232_0 <=( _mesh_14_7_io_out_a_0) ^ ((fiEnable && (249 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_233_0 <=( _mesh_14_8_io_out_a_0) ^ ((fiEnable && (250 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_234_0 <=( _mesh_14_9_io_out_a_0) ^ ((fiEnable && (251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_235_0 <=( _mesh_14_10_io_out_a_0) ^ ((fiEnable && (252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_236_0 <=( _mesh_14_11_io_out_a_0) ^ ((fiEnable && (253 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_237_0 <=( _mesh_14_12_io_out_a_0) ^ ((fiEnable && (254 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_238_0 <=( _mesh_14_13_io_out_a_0) ^ ((fiEnable && (255 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_239_0 <=( _mesh_14_14_io_out_a_0) ^ ((fiEnable && (256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_240_0 <=( io_in_a_15_0) ^ ((fiEnable && (257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_241_0 <=( _mesh_15_0_io_out_a_0) ^ ((fiEnable && (258 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_242_0 <=( _mesh_15_1_io_out_a_0) ^ ((fiEnable && (259 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_243_0 <=( _mesh_15_2_io_out_a_0) ^ ((fiEnable && (260 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_244_0 <=( _mesh_15_3_io_out_a_0) ^ ((fiEnable && (261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_245_0 <=( _mesh_15_4_io_out_a_0) ^ ((fiEnable && (262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_246_0 <=( _mesh_15_5_io_out_a_0) ^ ((fiEnable && (263 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_247_0 <=( _mesh_15_6_io_out_a_0) ^ ((fiEnable && (264 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_248_0 <=( _mesh_15_7_io_out_a_0) ^ ((fiEnable && (265 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_249_0 <=( _mesh_15_8_io_out_a_0) ^ ((fiEnable && (266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_250_0 <=( _mesh_15_9_io_out_a_0) ^ ((fiEnable && (267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_251_0 <=( _mesh_15_10_io_out_a_0) ^ ((fiEnable && (268 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_252_0 <=( _mesh_15_11_io_out_a_0) ^ ((fiEnable && (269 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_253_0 <=( _mesh_15_12_io_out_a_0) ^ ((fiEnable && (270 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_254_0 <=( _mesh_15_13_io_out_a_0) ^ ((fiEnable && (271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_255_0 <=( _mesh_15_14_io_out_a_0) ^ ((fiEnable && (272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		if (io_in_valid_0_0) begin
			b_0 <=( io_in_b_0_0) ^ ((fiEnable && (273 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_256_0 <=( io_in_d_0_0) ^ ((fiEnable && (274 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_0_io_in_control_0_shift_b <=( io_in_control_0_0_shift) ^ ((fiEnable && (275 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_0_io_in_control_0_dataflow_b <=( io_in_control_0_0_dataflow) ^ ((fiEnable && (276 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_0_io_in_control_0_propagate_b <=( io_in_control_0_0_propagate) ^ ((fiEnable && (277 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_0_io_out_valid_0) begin
			b_1_0 <=( _mesh_0_0_io_out_b_0) ^ ((fiEnable && (278 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_257_0 <=( _mesh_0_0_io_out_c_0) ^ ((fiEnable && (279 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_0_io_in_control_0_shift_b <=( _mesh_0_0_io_out_control_0_shift) ^ ((fiEnable && (280 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_0_io_in_control_0_dataflow_b <=( _mesh_0_0_io_out_control_0_dataflow) ^ ((fiEnable && (281 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_0_io_in_control_0_propagate_b <=( _mesh_0_0_io_out_control_0_propagate) ^ ((fiEnable && (282 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_0_io_out_valid_0) begin
			b_2_0 <=( _mesh_1_0_io_out_b_0) ^ ((fiEnable && (283 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_258_0 <=( _mesh_1_0_io_out_c_0) ^ ((fiEnable && (284 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_0_io_in_control_0_shift_b <=( _mesh_1_0_io_out_control_0_shift) ^ ((fiEnable && (285 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_0_io_in_control_0_dataflow_b <=( _mesh_1_0_io_out_control_0_dataflow) ^ ((fiEnable && (286 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_0_io_in_control_0_propagate_b <=( _mesh_1_0_io_out_control_0_propagate) ^ ((fiEnable && (287 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_0_io_out_valid_0) begin
			b_3_0 <=( _mesh_2_0_io_out_b_0) ^ ((fiEnable && (288 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_259_0 <=( _mesh_2_0_io_out_c_0) ^ ((fiEnable && (289 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_0_io_in_control_0_shift_b <=( _mesh_2_0_io_out_control_0_shift) ^ ((fiEnable && (290 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_0_io_in_control_0_dataflow_b <=( _mesh_2_0_io_out_control_0_dataflow) ^ ((fiEnable && (291 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_0_io_in_control_0_propagate_b <=( _mesh_2_0_io_out_control_0_propagate) ^ ((fiEnable && (292 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_0_io_out_valid_0) begin
			b_4_0 <=( _mesh_3_0_io_out_b_0) ^ ((fiEnable && (293 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_260_0 <=( _mesh_3_0_io_out_c_0) ^ ((fiEnable && (294 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_0_io_in_control_0_shift_b <=( _mesh_3_0_io_out_control_0_shift) ^ ((fiEnable && (295 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_0_io_in_control_0_dataflow_b <=( _mesh_3_0_io_out_control_0_dataflow) ^ ((fiEnable && (296 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_0_io_in_control_0_propagate_b <=( _mesh_3_0_io_out_control_0_propagate) ^ ((fiEnable && (297 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_0_io_out_valid_0) begin
			b_5_0 <=( _mesh_4_0_io_out_b_0) ^ ((fiEnable && (298 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_261_0 <=( _mesh_4_0_io_out_c_0) ^ ((fiEnable && (299 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_0_io_in_control_0_shift_b <=( _mesh_4_0_io_out_control_0_shift) ^ ((fiEnable && (300 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_0_io_in_control_0_dataflow_b <=( _mesh_4_0_io_out_control_0_dataflow) ^ ((fiEnable && (301 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_0_io_in_control_0_propagate_b <=( _mesh_4_0_io_out_control_0_propagate) ^ ((fiEnable && (302 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_0_io_out_valid_0) begin
			b_6_0 <=( _mesh_5_0_io_out_b_0) ^ ((fiEnable && (303 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_262_0 <=( _mesh_5_0_io_out_c_0) ^ ((fiEnable && (304 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_0_io_in_control_0_shift_b <=( _mesh_5_0_io_out_control_0_shift) ^ ((fiEnable && (305 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_0_io_in_control_0_dataflow_b <=( _mesh_5_0_io_out_control_0_dataflow) ^ ((fiEnable && (306 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_0_io_in_control_0_propagate_b <=( _mesh_5_0_io_out_control_0_propagate) ^ ((fiEnable && (307 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_0_io_out_valid_0) begin
			b_7_0 <=( _mesh_6_0_io_out_b_0) ^ ((fiEnable && (308 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_263_0 <=( _mesh_6_0_io_out_c_0) ^ ((fiEnable && (309 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_0_io_in_control_0_shift_b <=( _mesh_6_0_io_out_control_0_shift) ^ ((fiEnable && (310 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_0_io_in_control_0_dataflow_b <=( _mesh_6_0_io_out_control_0_dataflow) ^ ((fiEnable && (311 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_0_io_in_control_0_propagate_b <=( _mesh_6_0_io_out_control_0_propagate) ^ ((fiEnable && (312 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_0_io_out_valid_0) begin
			b_8_0 <=( _mesh_7_0_io_out_b_0) ^ ((fiEnable && (313 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_264_0 <=( _mesh_7_0_io_out_c_0) ^ ((fiEnable && (314 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_0_io_in_control_0_shift_b <=( _mesh_7_0_io_out_control_0_shift) ^ ((fiEnable && (315 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_0_io_in_control_0_dataflow_b <=( _mesh_7_0_io_out_control_0_dataflow) ^ ((fiEnable && (316 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_0_io_in_control_0_propagate_b <=( _mesh_7_0_io_out_control_0_propagate) ^ ((fiEnable && (317 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_0_io_out_valid_0) begin
			b_9_0 <=( _mesh_8_0_io_out_b_0) ^ ((fiEnable && (318 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_265_0 <=( _mesh_8_0_io_out_c_0) ^ ((fiEnable && (319 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_0_io_in_control_0_shift_b <=( _mesh_8_0_io_out_control_0_shift) ^ ((fiEnable && (320 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_0_io_in_control_0_dataflow_b <=( _mesh_8_0_io_out_control_0_dataflow) ^ ((fiEnable && (321 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_0_io_in_control_0_propagate_b <=( _mesh_8_0_io_out_control_0_propagate) ^ ((fiEnable && (322 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_0_io_out_valid_0) begin
			b_10_0 <=( _mesh_9_0_io_out_b_0) ^ ((fiEnable && (323 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_266_0 <=( _mesh_9_0_io_out_c_0) ^ ((fiEnable && (324 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_0_io_in_control_0_shift_b <=( _mesh_9_0_io_out_control_0_shift) ^ ((fiEnable && (325 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_0_io_in_control_0_dataflow_b <=( _mesh_9_0_io_out_control_0_dataflow) ^ ((fiEnable && (326 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_0_io_in_control_0_propagate_b <=( _mesh_9_0_io_out_control_0_propagate) ^ ((fiEnable && (327 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_0_io_out_valid_0) begin
			b_11_0 <=( _mesh_10_0_io_out_b_0) ^ ((fiEnable && (328 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_267_0 <=( _mesh_10_0_io_out_c_0) ^ ((fiEnable && (329 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_0_io_in_control_0_shift_b <=( _mesh_10_0_io_out_control_0_shift) ^ ((fiEnable && (330 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_0_io_in_control_0_dataflow_b <=( _mesh_10_0_io_out_control_0_dataflow) ^ ((fiEnable && (331 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_0_io_in_control_0_propagate_b <=( _mesh_10_0_io_out_control_0_propagate) ^ ((fiEnable && (332 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_0_io_out_valid_0) begin
			b_12_0 <=( _mesh_11_0_io_out_b_0) ^ ((fiEnable && (333 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_268_0 <=( _mesh_11_0_io_out_c_0) ^ ((fiEnable && (334 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_0_io_in_control_0_shift_b <=( _mesh_11_0_io_out_control_0_shift) ^ ((fiEnable && (335 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_0_io_in_control_0_dataflow_b <=( _mesh_11_0_io_out_control_0_dataflow) ^ ((fiEnable && (336 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_0_io_in_control_0_propagate_b <=( _mesh_11_0_io_out_control_0_propagate) ^ ((fiEnable && (337 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_0_io_out_valid_0) begin
			b_13_0 <=( _mesh_12_0_io_out_b_0) ^ ((fiEnable && (338 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_269_0 <=( _mesh_12_0_io_out_c_0) ^ ((fiEnable && (339 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_0_io_in_control_0_shift_b <=( _mesh_12_0_io_out_control_0_shift) ^ ((fiEnable && (340 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_0_io_in_control_0_dataflow_b <=( _mesh_12_0_io_out_control_0_dataflow) ^ ((fiEnable && (341 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_0_io_in_control_0_propagate_b <=( _mesh_12_0_io_out_control_0_propagate) ^ ((fiEnable && (342 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_0_io_out_valid_0) begin
			b_14_0 <=( _mesh_13_0_io_out_b_0) ^ ((fiEnable && (343 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_270_0 <=( _mesh_13_0_io_out_c_0) ^ ((fiEnable && (344 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_0_io_in_control_0_shift_b <=( _mesh_13_0_io_out_control_0_shift) ^ ((fiEnable && (345 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_0_io_in_control_0_dataflow_b <=( _mesh_13_0_io_out_control_0_dataflow) ^ ((fiEnable && (346 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_0_io_in_control_0_propagate_b <=( _mesh_13_0_io_out_control_0_propagate) ^ ((fiEnable && (347 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_0_io_out_valid_0) begin
			b_15_0 <=( _mesh_14_0_io_out_b_0) ^ ((fiEnable && (348 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_271_0 <=( _mesh_14_0_io_out_c_0) ^ ((fiEnable && (349 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_0_io_in_control_0_shift_b <=( _mesh_14_0_io_out_control_0_shift) ^ ((fiEnable && (350 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_0_io_in_control_0_dataflow_b <=( _mesh_14_0_io_out_control_0_dataflow) ^ ((fiEnable && (351 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_0_io_in_control_0_propagate_b <=( _mesh_14_0_io_out_control_0_propagate) ^ ((fiEnable && (352 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_1_0) begin
			b_16_0 <=( io_in_b_1_0) ^ ((fiEnable && (353 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_272_0 <=( io_in_d_1_0) ^ ((fiEnable && (354 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_1_io_in_control_0_shift_b <=( io_in_control_1_0_shift) ^ ((fiEnable && (355 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_1_io_in_control_0_dataflow_b <=( io_in_control_1_0_dataflow) ^ ((fiEnable && (356 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_1_io_in_control_0_propagate_b <=( io_in_control_1_0_propagate) ^ ((fiEnable && (357 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_1_io_out_valid_0) begin
			b_17_0 <=( _mesh_0_1_io_out_b_0) ^ ((fiEnable && (358 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_273_0 <=( _mesh_0_1_io_out_c_0) ^ ((fiEnable && (359 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_1_io_in_control_0_shift_b <=( _mesh_0_1_io_out_control_0_shift) ^ ((fiEnable && (360 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_1_io_in_control_0_dataflow_b <=( _mesh_0_1_io_out_control_0_dataflow) ^ ((fiEnable && (361 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_1_io_in_control_0_propagate_b <=( _mesh_0_1_io_out_control_0_propagate) ^ ((fiEnable && (362 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_1_io_out_valid_0) begin
			b_18_0 <=( _mesh_1_1_io_out_b_0) ^ ((fiEnable && (363 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_274_0 <=( _mesh_1_1_io_out_c_0) ^ ((fiEnable && (364 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_1_io_in_control_0_shift_b <=( _mesh_1_1_io_out_control_0_shift) ^ ((fiEnable && (365 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_1_io_in_control_0_dataflow_b <=( _mesh_1_1_io_out_control_0_dataflow) ^ ((fiEnable && (366 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_1_io_in_control_0_propagate_b <=( _mesh_1_1_io_out_control_0_propagate) ^ ((fiEnable && (367 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_1_io_out_valid_0) begin
			b_19_0 <=( _mesh_2_1_io_out_b_0) ^ ((fiEnable && (368 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_275_0 <=( _mesh_2_1_io_out_c_0) ^ ((fiEnable && (369 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_1_io_in_control_0_shift_b <=( _mesh_2_1_io_out_control_0_shift) ^ ((fiEnable && (370 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_1_io_in_control_0_dataflow_b <=( _mesh_2_1_io_out_control_0_dataflow) ^ ((fiEnable && (371 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_1_io_in_control_0_propagate_b <=( _mesh_2_1_io_out_control_0_propagate) ^ ((fiEnable && (372 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_1_io_out_valid_0) begin
			b_20_0 <=( _mesh_3_1_io_out_b_0) ^ ((fiEnable && (373 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_276_0 <=( _mesh_3_1_io_out_c_0) ^ ((fiEnable && (374 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_1_io_in_control_0_shift_b <=( _mesh_3_1_io_out_control_0_shift) ^ ((fiEnable && (375 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_1_io_in_control_0_dataflow_b <=( _mesh_3_1_io_out_control_0_dataflow) ^ ((fiEnable && (376 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_1_io_in_control_0_propagate_b <=( _mesh_3_1_io_out_control_0_propagate) ^ ((fiEnable && (377 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_1_io_out_valid_0) begin
			b_21_0 <=( _mesh_4_1_io_out_b_0) ^ ((fiEnable && (378 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_277_0 <=( _mesh_4_1_io_out_c_0) ^ ((fiEnable && (379 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_1_io_in_control_0_shift_b <=( _mesh_4_1_io_out_control_0_shift) ^ ((fiEnable && (380 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_1_io_in_control_0_dataflow_b <=( _mesh_4_1_io_out_control_0_dataflow) ^ ((fiEnable && (381 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_1_io_in_control_0_propagate_b <=( _mesh_4_1_io_out_control_0_propagate) ^ ((fiEnable && (382 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_1_io_out_valid_0) begin
			b_22_0 <=( _mesh_5_1_io_out_b_0) ^ ((fiEnable && (383 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_278_0 <=( _mesh_5_1_io_out_c_0) ^ ((fiEnable && (384 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_1_io_in_control_0_shift_b <=( _mesh_5_1_io_out_control_0_shift) ^ ((fiEnable && (385 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_1_io_in_control_0_dataflow_b <=( _mesh_5_1_io_out_control_0_dataflow) ^ ((fiEnable && (386 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_1_io_in_control_0_propagate_b <=( _mesh_5_1_io_out_control_0_propagate) ^ ((fiEnable && (387 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_1_io_out_valid_0) begin
			b_23_0 <=( _mesh_6_1_io_out_b_0) ^ ((fiEnable && (388 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_279_0 <=( _mesh_6_1_io_out_c_0) ^ ((fiEnable && (389 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_1_io_in_control_0_shift_b <=( _mesh_6_1_io_out_control_0_shift) ^ ((fiEnable && (390 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_1_io_in_control_0_dataflow_b <=( _mesh_6_1_io_out_control_0_dataflow) ^ ((fiEnable && (391 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_1_io_in_control_0_propagate_b <=( _mesh_6_1_io_out_control_0_propagate) ^ ((fiEnable && (392 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_1_io_out_valid_0) begin
			b_24_0 <=( _mesh_7_1_io_out_b_0) ^ ((fiEnable && (393 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_280_0 <=( _mesh_7_1_io_out_c_0) ^ ((fiEnable && (394 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_1_io_in_control_0_shift_b <=( _mesh_7_1_io_out_control_0_shift) ^ ((fiEnable && (395 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_1_io_in_control_0_dataflow_b <=( _mesh_7_1_io_out_control_0_dataflow) ^ ((fiEnable && (396 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_1_io_in_control_0_propagate_b <=( _mesh_7_1_io_out_control_0_propagate) ^ ((fiEnable && (397 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_1_io_out_valid_0) begin
			b_25_0 <=( _mesh_8_1_io_out_b_0) ^ ((fiEnable && (398 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_281_0 <=( _mesh_8_1_io_out_c_0) ^ ((fiEnable && (399 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_1_io_in_control_0_shift_b <=( _mesh_8_1_io_out_control_0_shift) ^ ((fiEnable && (400 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_1_io_in_control_0_dataflow_b <=( _mesh_8_1_io_out_control_0_dataflow) ^ ((fiEnable && (401 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_1_io_in_control_0_propagate_b <=( _mesh_8_1_io_out_control_0_propagate) ^ ((fiEnable && (402 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_1_io_out_valid_0) begin
			b_26_0 <=( _mesh_9_1_io_out_b_0) ^ ((fiEnable && (403 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_282_0 <=( _mesh_9_1_io_out_c_0) ^ ((fiEnable && (404 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_1_io_in_control_0_shift_b <=( _mesh_9_1_io_out_control_0_shift) ^ ((fiEnable && (405 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_1_io_in_control_0_dataflow_b <=( _mesh_9_1_io_out_control_0_dataflow) ^ ((fiEnable && (406 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_1_io_in_control_0_propagate_b <=( _mesh_9_1_io_out_control_0_propagate) ^ ((fiEnable && (407 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_1_io_out_valid_0) begin
			b_27_0 <=( _mesh_10_1_io_out_b_0) ^ ((fiEnable && (408 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_283_0 <=( _mesh_10_1_io_out_c_0) ^ ((fiEnable && (409 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_1_io_in_control_0_shift_b <=( _mesh_10_1_io_out_control_0_shift) ^ ((fiEnable && (410 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_1_io_in_control_0_dataflow_b <=( _mesh_10_1_io_out_control_0_dataflow) ^ ((fiEnable && (411 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_1_io_in_control_0_propagate_b <=( _mesh_10_1_io_out_control_0_propagate) ^ ((fiEnable && (412 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_1_io_out_valid_0) begin
			b_28_0 <=( _mesh_11_1_io_out_b_0) ^ ((fiEnable && (413 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_284_0 <=( _mesh_11_1_io_out_c_0) ^ ((fiEnable && (414 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_1_io_in_control_0_shift_b <=( _mesh_11_1_io_out_control_0_shift) ^ ((fiEnable && (415 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_1_io_in_control_0_dataflow_b <=( _mesh_11_1_io_out_control_0_dataflow) ^ ((fiEnable && (416 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_1_io_in_control_0_propagate_b <=( _mesh_11_1_io_out_control_0_propagate) ^ ((fiEnable && (417 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_1_io_out_valid_0) begin
			b_29_0 <=( _mesh_12_1_io_out_b_0) ^ ((fiEnable && (418 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_285_0 <=( _mesh_12_1_io_out_c_0) ^ ((fiEnable && (419 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_1_io_in_control_0_shift_b <=( _mesh_12_1_io_out_control_0_shift) ^ ((fiEnable && (420 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_1_io_in_control_0_dataflow_b <=( _mesh_12_1_io_out_control_0_dataflow) ^ ((fiEnable && (421 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_1_io_in_control_0_propagate_b <=( _mesh_12_1_io_out_control_0_propagate) ^ ((fiEnable && (422 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_1_io_out_valid_0) begin
			b_30_0 <=( _mesh_13_1_io_out_b_0) ^ ((fiEnable && (423 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_286_0 <=( _mesh_13_1_io_out_c_0) ^ ((fiEnable && (424 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_1_io_in_control_0_shift_b <=( _mesh_13_1_io_out_control_0_shift) ^ ((fiEnable && (425 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_1_io_in_control_0_dataflow_b <=( _mesh_13_1_io_out_control_0_dataflow) ^ ((fiEnable && (426 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_1_io_in_control_0_propagate_b <=( _mesh_13_1_io_out_control_0_propagate) ^ ((fiEnable && (427 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_1_io_out_valid_0) begin
			b_31_0 <=( _mesh_14_1_io_out_b_0) ^ ((fiEnable && (428 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_287_0 <=( _mesh_14_1_io_out_c_0) ^ ((fiEnable && (429 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_1_io_in_control_0_shift_b <=( _mesh_14_1_io_out_control_0_shift) ^ ((fiEnable && (430 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_1_io_in_control_0_dataflow_b <=( _mesh_14_1_io_out_control_0_dataflow) ^ ((fiEnable && (431 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_1_io_in_control_0_propagate_b <=( _mesh_14_1_io_out_control_0_propagate) ^ ((fiEnable && (432 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_2_0) begin
			b_32_0 <=( io_in_b_2_0) ^ ((fiEnable && (433 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_288_0 <=( io_in_d_2_0) ^ ((fiEnable && (434 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_2_io_in_control_0_shift_b <=( io_in_control_2_0_shift) ^ ((fiEnable && (435 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_2_io_in_control_0_dataflow_b <=( io_in_control_2_0_dataflow) ^ ((fiEnable && (436 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_2_io_in_control_0_propagate_b <=( io_in_control_2_0_propagate) ^ ((fiEnable && (437 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_2_io_out_valid_0) begin
			b_33_0 <=( _mesh_0_2_io_out_b_0) ^ ((fiEnable && (438 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_289_0 <=( _mesh_0_2_io_out_c_0) ^ ((fiEnable && (439 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_2_io_in_control_0_shift_b <=( _mesh_0_2_io_out_control_0_shift) ^ ((fiEnable && (440 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_2_io_in_control_0_dataflow_b <=( _mesh_0_2_io_out_control_0_dataflow) ^ ((fiEnable && (441 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_2_io_in_control_0_propagate_b <=( _mesh_0_2_io_out_control_0_propagate) ^ ((fiEnable && (442 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_2_io_out_valid_0) begin
			b_34_0 <=( _mesh_1_2_io_out_b_0) ^ ((fiEnable && (443 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_290_0 <=( _mesh_1_2_io_out_c_0) ^ ((fiEnable && (444 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_2_io_in_control_0_shift_b <=( _mesh_1_2_io_out_control_0_shift) ^ ((fiEnable && (445 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_2_io_in_control_0_dataflow_b <=( _mesh_1_2_io_out_control_0_dataflow) ^ ((fiEnable && (446 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_2_io_in_control_0_propagate_b <=( _mesh_1_2_io_out_control_0_propagate) ^ ((fiEnable && (447 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_2_io_out_valid_0) begin
			b_35_0 <=( _mesh_2_2_io_out_b_0) ^ ((fiEnable && (448 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_291_0 <=( _mesh_2_2_io_out_c_0) ^ ((fiEnable && (449 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_2_io_in_control_0_shift_b <=( _mesh_2_2_io_out_control_0_shift) ^ ((fiEnable && (450 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_2_io_in_control_0_dataflow_b <=( _mesh_2_2_io_out_control_0_dataflow) ^ ((fiEnable && (451 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_2_io_in_control_0_propagate_b <=( _mesh_2_2_io_out_control_0_propagate) ^ ((fiEnable && (452 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_2_io_out_valid_0) begin
			b_36_0 <=( _mesh_3_2_io_out_b_0) ^ ((fiEnable && (453 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_292_0 <=( _mesh_3_2_io_out_c_0) ^ ((fiEnable && (454 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_2_io_in_control_0_shift_b <=( _mesh_3_2_io_out_control_0_shift) ^ ((fiEnable && (455 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_2_io_in_control_0_dataflow_b <=( _mesh_3_2_io_out_control_0_dataflow) ^ ((fiEnable && (456 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_2_io_in_control_0_propagate_b <=( _mesh_3_2_io_out_control_0_propagate) ^ ((fiEnable && (457 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_2_io_out_valid_0) begin
			b_37_0 <=( _mesh_4_2_io_out_b_0) ^ ((fiEnable && (458 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_293_0 <=( _mesh_4_2_io_out_c_0) ^ ((fiEnable && (459 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_2_io_in_control_0_shift_b <=( _mesh_4_2_io_out_control_0_shift) ^ ((fiEnable && (460 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_2_io_in_control_0_dataflow_b <=( _mesh_4_2_io_out_control_0_dataflow) ^ ((fiEnable && (461 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_2_io_in_control_0_propagate_b <=( _mesh_4_2_io_out_control_0_propagate) ^ ((fiEnable && (462 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_2_io_out_valid_0) begin
			b_38_0 <=( _mesh_5_2_io_out_b_0) ^ ((fiEnable && (463 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_294_0 <=( _mesh_5_2_io_out_c_0) ^ ((fiEnable && (464 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_2_io_in_control_0_shift_b <=( _mesh_5_2_io_out_control_0_shift) ^ ((fiEnable && (465 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_2_io_in_control_0_dataflow_b <=( _mesh_5_2_io_out_control_0_dataflow) ^ ((fiEnable && (466 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_2_io_in_control_0_propagate_b <=( _mesh_5_2_io_out_control_0_propagate) ^ ((fiEnable && (467 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_2_io_out_valid_0) begin
			b_39_0 <=( _mesh_6_2_io_out_b_0) ^ ((fiEnable && (468 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_295_0 <=( _mesh_6_2_io_out_c_0) ^ ((fiEnable && (469 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_2_io_in_control_0_shift_b <=( _mesh_6_2_io_out_control_0_shift) ^ ((fiEnable && (470 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_2_io_in_control_0_dataflow_b <=( _mesh_6_2_io_out_control_0_dataflow) ^ ((fiEnable && (471 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_2_io_in_control_0_propagate_b <=( _mesh_6_2_io_out_control_0_propagate) ^ ((fiEnable && (472 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_2_io_out_valid_0) begin
			b_40_0 <=( _mesh_7_2_io_out_b_0) ^ ((fiEnable && (473 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_296_0 <=( _mesh_7_2_io_out_c_0) ^ ((fiEnable && (474 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_2_io_in_control_0_shift_b <=( _mesh_7_2_io_out_control_0_shift) ^ ((fiEnable && (475 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_2_io_in_control_0_dataflow_b <=( _mesh_7_2_io_out_control_0_dataflow) ^ ((fiEnable && (476 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_2_io_in_control_0_propagate_b <=( _mesh_7_2_io_out_control_0_propagate) ^ ((fiEnable && (477 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_2_io_out_valid_0) begin
			b_41_0 <=( _mesh_8_2_io_out_b_0) ^ ((fiEnable && (478 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_297_0 <=( _mesh_8_2_io_out_c_0) ^ ((fiEnable && (479 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_2_io_in_control_0_shift_b <=( _mesh_8_2_io_out_control_0_shift) ^ ((fiEnable && (480 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_2_io_in_control_0_dataflow_b <=( _mesh_8_2_io_out_control_0_dataflow) ^ ((fiEnable && (481 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_2_io_in_control_0_propagate_b <=( _mesh_8_2_io_out_control_0_propagate) ^ ((fiEnable && (482 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_2_io_out_valid_0) begin
			b_42_0 <=( _mesh_9_2_io_out_b_0) ^ ((fiEnable && (483 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_298_0 <=( _mesh_9_2_io_out_c_0) ^ ((fiEnable && (484 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_2_io_in_control_0_shift_b <=( _mesh_9_2_io_out_control_0_shift) ^ ((fiEnable && (485 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_2_io_in_control_0_dataflow_b <=( _mesh_9_2_io_out_control_0_dataflow) ^ ((fiEnable && (486 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_2_io_in_control_0_propagate_b <=( _mesh_9_2_io_out_control_0_propagate) ^ ((fiEnable && (487 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_2_io_out_valid_0) begin
			b_43_0 <=( _mesh_10_2_io_out_b_0) ^ ((fiEnable && (488 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_299_0 <=( _mesh_10_2_io_out_c_0) ^ ((fiEnable && (489 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_2_io_in_control_0_shift_b <=( _mesh_10_2_io_out_control_0_shift) ^ ((fiEnable && (490 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_2_io_in_control_0_dataflow_b <=( _mesh_10_2_io_out_control_0_dataflow) ^ ((fiEnable && (491 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_2_io_in_control_0_propagate_b <=( _mesh_10_2_io_out_control_0_propagate) ^ ((fiEnable && (492 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_2_io_out_valid_0) begin
			b_44_0 <=( _mesh_11_2_io_out_b_0) ^ ((fiEnable && (493 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_300_0 <=( _mesh_11_2_io_out_c_0) ^ ((fiEnable && (494 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_2_io_in_control_0_shift_b <=( _mesh_11_2_io_out_control_0_shift) ^ ((fiEnable && (495 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_2_io_in_control_0_dataflow_b <=( _mesh_11_2_io_out_control_0_dataflow) ^ ((fiEnable && (496 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_2_io_in_control_0_propagate_b <=( _mesh_11_2_io_out_control_0_propagate) ^ ((fiEnable && (497 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_2_io_out_valid_0) begin
			b_45_0 <=( _mesh_12_2_io_out_b_0) ^ ((fiEnable && (498 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_301_0 <=( _mesh_12_2_io_out_c_0) ^ ((fiEnable && (499 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_2_io_in_control_0_shift_b <=( _mesh_12_2_io_out_control_0_shift) ^ ((fiEnable && (500 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_2_io_in_control_0_dataflow_b <=( _mesh_12_2_io_out_control_0_dataflow) ^ ((fiEnable && (501 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_2_io_in_control_0_propagate_b <=( _mesh_12_2_io_out_control_0_propagate) ^ ((fiEnable && (502 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_2_io_out_valid_0) begin
			b_46_0 <=( _mesh_13_2_io_out_b_0) ^ ((fiEnable && (503 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_302_0 <=( _mesh_13_2_io_out_c_0) ^ ((fiEnable && (504 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_2_io_in_control_0_shift_b <=( _mesh_13_2_io_out_control_0_shift) ^ ((fiEnable && (505 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_2_io_in_control_0_dataflow_b <=( _mesh_13_2_io_out_control_0_dataflow) ^ ((fiEnable && (506 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_2_io_in_control_0_propagate_b <=( _mesh_13_2_io_out_control_0_propagate) ^ ((fiEnable && (507 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_2_io_out_valid_0) begin
			b_47_0 <=( _mesh_14_2_io_out_b_0) ^ ((fiEnable && (508 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_303_0 <=( _mesh_14_2_io_out_c_0) ^ ((fiEnable && (509 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_2_io_in_control_0_shift_b <=( _mesh_14_2_io_out_control_0_shift) ^ ((fiEnable && (510 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_2_io_in_control_0_dataflow_b <=( _mesh_14_2_io_out_control_0_dataflow) ^ ((fiEnable && (511 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_2_io_in_control_0_propagate_b <=( _mesh_14_2_io_out_control_0_propagate) ^ ((fiEnable && (512 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_3_0) begin
			b_48_0 <=( io_in_b_3_0) ^ ((fiEnable && (513 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_304_0 <=( io_in_d_3_0) ^ ((fiEnable && (514 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_3_io_in_control_0_shift_b <=( io_in_control_3_0_shift) ^ ((fiEnable && (515 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_3_io_in_control_0_dataflow_b <=( io_in_control_3_0_dataflow) ^ ((fiEnable && (516 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_3_io_in_control_0_propagate_b <=( io_in_control_3_0_propagate) ^ ((fiEnable && (517 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_3_io_out_valid_0) begin
			b_49_0 <=( _mesh_0_3_io_out_b_0) ^ ((fiEnable && (518 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_305_0 <=( _mesh_0_3_io_out_c_0) ^ ((fiEnable && (519 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_3_io_in_control_0_shift_b <=( _mesh_0_3_io_out_control_0_shift) ^ ((fiEnable && (520 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_3_io_in_control_0_dataflow_b <=( _mesh_0_3_io_out_control_0_dataflow) ^ ((fiEnable && (521 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_3_io_in_control_0_propagate_b <=( _mesh_0_3_io_out_control_0_propagate) ^ ((fiEnable && (522 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_3_io_out_valid_0) begin
			b_50_0 <=( _mesh_1_3_io_out_b_0) ^ ((fiEnable && (523 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_306_0 <=( _mesh_1_3_io_out_c_0) ^ ((fiEnable && (524 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_3_io_in_control_0_shift_b <=( _mesh_1_3_io_out_control_0_shift) ^ ((fiEnable && (525 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_3_io_in_control_0_dataflow_b <=( _mesh_1_3_io_out_control_0_dataflow) ^ ((fiEnable && (526 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_3_io_in_control_0_propagate_b <=( _mesh_1_3_io_out_control_0_propagate) ^ ((fiEnable && (527 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_3_io_out_valid_0) begin
			b_51_0 <=( _mesh_2_3_io_out_b_0) ^ ((fiEnable && (528 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_307_0 <=( _mesh_2_3_io_out_c_0) ^ ((fiEnable && (529 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_3_io_in_control_0_shift_b <=( _mesh_2_3_io_out_control_0_shift) ^ ((fiEnable && (530 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_3_io_in_control_0_dataflow_b <=( _mesh_2_3_io_out_control_0_dataflow) ^ ((fiEnable && (531 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_3_io_in_control_0_propagate_b <=( _mesh_2_3_io_out_control_0_propagate) ^ ((fiEnable && (532 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_3_io_out_valid_0) begin
			b_52_0 <=( _mesh_3_3_io_out_b_0) ^ ((fiEnable && (533 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_308_0 <=( _mesh_3_3_io_out_c_0) ^ ((fiEnable && (534 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_3_io_in_control_0_shift_b <=( _mesh_3_3_io_out_control_0_shift) ^ ((fiEnable && (535 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_3_io_in_control_0_dataflow_b <=( _mesh_3_3_io_out_control_0_dataflow) ^ ((fiEnable && (536 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_3_io_in_control_0_propagate_b <=( _mesh_3_3_io_out_control_0_propagate) ^ ((fiEnable && (537 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_3_io_out_valid_0) begin
			b_53_0 <=( _mesh_4_3_io_out_b_0) ^ ((fiEnable && (538 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_309_0 <=( _mesh_4_3_io_out_c_0) ^ ((fiEnable && (539 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_3_io_in_control_0_shift_b <=( _mesh_4_3_io_out_control_0_shift) ^ ((fiEnable && (540 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_3_io_in_control_0_dataflow_b <=( _mesh_4_3_io_out_control_0_dataflow) ^ ((fiEnable && (541 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_3_io_in_control_0_propagate_b <=( _mesh_4_3_io_out_control_0_propagate) ^ ((fiEnable && (542 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_3_io_out_valid_0) begin
			b_54_0 <=( _mesh_5_3_io_out_b_0) ^ ((fiEnable && (543 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_310_0 <=( _mesh_5_3_io_out_c_0) ^ ((fiEnable && (544 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_3_io_in_control_0_shift_b <=( _mesh_5_3_io_out_control_0_shift) ^ ((fiEnable && (545 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_3_io_in_control_0_dataflow_b <=( _mesh_5_3_io_out_control_0_dataflow) ^ ((fiEnable && (546 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_3_io_in_control_0_propagate_b <=( _mesh_5_3_io_out_control_0_propagate) ^ ((fiEnable && (547 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_3_io_out_valid_0) begin
			b_55_0 <=( _mesh_6_3_io_out_b_0) ^ ((fiEnable && (548 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_311_0 <=( _mesh_6_3_io_out_c_0) ^ ((fiEnable && (549 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_3_io_in_control_0_shift_b <=( _mesh_6_3_io_out_control_0_shift) ^ ((fiEnable && (550 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_3_io_in_control_0_dataflow_b <=( _mesh_6_3_io_out_control_0_dataflow) ^ ((fiEnable && (551 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_3_io_in_control_0_propagate_b <=( _mesh_6_3_io_out_control_0_propagate) ^ ((fiEnable && (552 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_3_io_out_valid_0) begin
			b_56_0 <=( _mesh_7_3_io_out_b_0) ^ ((fiEnable && (553 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_312_0 <=( _mesh_7_3_io_out_c_0) ^ ((fiEnable && (554 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_3_io_in_control_0_shift_b <=( _mesh_7_3_io_out_control_0_shift) ^ ((fiEnable && (555 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_3_io_in_control_0_dataflow_b <=( _mesh_7_3_io_out_control_0_dataflow) ^ ((fiEnable && (556 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_3_io_in_control_0_propagate_b <=( _mesh_7_3_io_out_control_0_propagate) ^ ((fiEnable && (557 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_3_io_out_valid_0) begin
			b_57_0 <=( _mesh_8_3_io_out_b_0) ^ ((fiEnable && (558 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_313_0 <=( _mesh_8_3_io_out_c_0) ^ ((fiEnable && (559 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_3_io_in_control_0_shift_b <=( _mesh_8_3_io_out_control_0_shift) ^ ((fiEnable && (560 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_3_io_in_control_0_dataflow_b <=( _mesh_8_3_io_out_control_0_dataflow) ^ ((fiEnable && (561 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_3_io_in_control_0_propagate_b <=( _mesh_8_3_io_out_control_0_propagate) ^ ((fiEnable && (562 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_3_io_out_valid_0) begin
			b_58_0 <=( _mesh_9_3_io_out_b_0) ^ ((fiEnable && (563 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_314_0 <=( _mesh_9_3_io_out_c_0) ^ ((fiEnable && (564 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_3_io_in_control_0_shift_b <=( _mesh_9_3_io_out_control_0_shift) ^ ((fiEnable && (565 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_3_io_in_control_0_dataflow_b <=( _mesh_9_3_io_out_control_0_dataflow) ^ ((fiEnable && (566 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_3_io_in_control_0_propagate_b <=( _mesh_9_3_io_out_control_0_propagate) ^ ((fiEnable && (567 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_3_io_out_valid_0) begin
			b_59_0 <=( _mesh_10_3_io_out_b_0) ^ ((fiEnable && (568 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_315_0 <=( _mesh_10_3_io_out_c_0) ^ ((fiEnable && (569 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_3_io_in_control_0_shift_b <=( _mesh_10_3_io_out_control_0_shift) ^ ((fiEnable && (570 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_3_io_in_control_0_dataflow_b <=( _mesh_10_3_io_out_control_0_dataflow) ^ ((fiEnable && (571 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_3_io_in_control_0_propagate_b <=( _mesh_10_3_io_out_control_0_propagate) ^ ((fiEnable && (572 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_3_io_out_valid_0) begin
			b_60_0 <=( _mesh_11_3_io_out_b_0) ^ ((fiEnable && (573 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_316_0 <=( _mesh_11_3_io_out_c_0) ^ ((fiEnable && (574 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_3_io_in_control_0_shift_b <=( _mesh_11_3_io_out_control_0_shift) ^ ((fiEnable && (575 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_3_io_in_control_0_dataflow_b <=( _mesh_11_3_io_out_control_0_dataflow) ^ ((fiEnable && (576 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_3_io_in_control_0_propagate_b <=( _mesh_11_3_io_out_control_0_propagate) ^ ((fiEnable && (577 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_3_io_out_valid_0) begin
			b_61_0 <=( _mesh_12_3_io_out_b_0) ^ ((fiEnable && (578 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_317_0 <=( _mesh_12_3_io_out_c_0) ^ ((fiEnable && (579 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_3_io_in_control_0_shift_b <=( _mesh_12_3_io_out_control_0_shift) ^ ((fiEnable && (580 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_3_io_in_control_0_dataflow_b <=( _mesh_12_3_io_out_control_0_dataflow) ^ ((fiEnable && (581 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_3_io_in_control_0_propagate_b <=( _mesh_12_3_io_out_control_0_propagate) ^ ((fiEnable && (582 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_3_io_out_valid_0) begin
			b_62_0 <=( _mesh_13_3_io_out_b_0) ^ ((fiEnable && (583 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_318_0 <=( _mesh_13_3_io_out_c_0) ^ ((fiEnable && (584 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_3_io_in_control_0_shift_b <=( _mesh_13_3_io_out_control_0_shift) ^ ((fiEnable && (585 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_3_io_in_control_0_dataflow_b <=( _mesh_13_3_io_out_control_0_dataflow) ^ ((fiEnable && (586 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_3_io_in_control_0_propagate_b <=( _mesh_13_3_io_out_control_0_propagate) ^ ((fiEnable && (587 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_3_io_out_valid_0) begin
			b_63_0 <=( _mesh_14_3_io_out_b_0) ^ ((fiEnable && (588 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_319_0 <=( _mesh_14_3_io_out_c_0) ^ ((fiEnable && (589 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_3_io_in_control_0_shift_b <=( _mesh_14_3_io_out_control_0_shift) ^ ((fiEnable && (590 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_3_io_in_control_0_dataflow_b <=( _mesh_14_3_io_out_control_0_dataflow) ^ ((fiEnable && (591 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_3_io_in_control_0_propagate_b <=( _mesh_14_3_io_out_control_0_propagate) ^ ((fiEnable && (592 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_4_0) begin
			b_64_0 <=( io_in_b_4_0) ^ ((fiEnable && (593 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_320_0 <=( io_in_d_4_0) ^ ((fiEnable && (594 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_4_io_in_control_0_shift_b <=( io_in_control_4_0_shift) ^ ((fiEnable && (595 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_4_io_in_control_0_dataflow_b <=( io_in_control_4_0_dataflow) ^ ((fiEnable && (596 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_4_io_in_control_0_propagate_b <=( io_in_control_4_0_propagate) ^ ((fiEnable && (597 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_4_io_out_valid_0) begin
			b_65_0 <=( _mesh_0_4_io_out_b_0) ^ ((fiEnable && (598 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_321_0 <=( _mesh_0_4_io_out_c_0) ^ ((fiEnable && (599 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_4_io_in_control_0_shift_b <=( _mesh_0_4_io_out_control_0_shift) ^ ((fiEnable && (600 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_4_io_in_control_0_dataflow_b <=( _mesh_0_4_io_out_control_0_dataflow) ^ ((fiEnable && (601 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_4_io_in_control_0_propagate_b <=( _mesh_0_4_io_out_control_0_propagate) ^ ((fiEnable && (602 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_4_io_out_valid_0) begin
			b_66_0 <=( _mesh_1_4_io_out_b_0) ^ ((fiEnable && (603 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_322_0 <=( _mesh_1_4_io_out_c_0) ^ ((fiEnable && (604 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_4_io_in_control_0_shift_b <=( _mesh_1_4_io_out_control_0_shift) ^ ((fiEnable && (605 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_4_io_in_control_0_dataflow_b <=( _mesh_1_4_io_out_control_0_dataflow) ^ ((fiEnable && (606 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_4_io_in_control_0_propagate_b <=( _mesh_1_4_io_out_control_0_propagate) ^ ((fiEnable && (607 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_4_io_out_valid_0) begin
			b_67_0 <=( _mesh_2_4_io_out_b_0) ^ ((fiEnable && (608 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_323_0 <=( _mesh_2_4_io_out_c_0) ^ ((fiEnable && (609 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_4_io_in_control_0_shift_b <=( _mesh_2_4_io_out_control_0_shift) ^ ((fiEnable && (610 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_4_io_in_control_0_dataflow_b <=( _mesh_2_4_io_out_control_0_dataflow) ^ ((fiEnable && (611 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_4_io_in_control_0_propagate_b <=( _mesh_2_4_io_out_control_0_propagate) ^ ((fiEnable && (612 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_4_io_out_valid_0) begin
			b_68_0 <=( _mesh_3_4_io_out_b_0) ^ ((fiEnable && (613 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_324_0 <=( _mesh_3_4_io_out_c_0) ^ ((fiEnable && (614 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_4_io_in_control_0_shift_b <=( _mesh_3_4_io_out_control_0_shift) ^ ((fiEnable && (615 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_4_io_in_control_0_dataflow_b <=( _mesh_3_4_io_out_control_0_dataflow) ^ ((fiEnable && (616 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_4_io_in_control_0_propagate_b <=( _mesh_3_4_io_out_control_0_propagate) ^ ((fiEnable && (617 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_4_io_out_valid_0) begin
			b_69_0 <=( _mesh_4_4_io_out_b_0) ^ ((fiEnable && (618 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_325_0 <=( _mesh_4_4_io_out_c_0) ^ ((fiEnable && (619 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_4_io_in_control_0_shift_b <=( _mesh_4_4_io_out_control_0_shift) ^ ((fiEnable && (620 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_4_io_in_control_0_dataflow_b <=( _mesh_4_4_io_out_control_0_dataflow) ^ ((fiEnable && (621 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_4_io_in_control_0_propagate_b <=( _mesh_4_4_io_out_control_0_propagate) ^ ((fiEnable && (622 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_4_io_out_valid_0) begin
			b_70_0 <=( _mesh_5_4_io_out_b_0) ^ ((fiEnable && (623 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_326_0 <=( _mesh_5_4_io_out_c_0) ^ ((fiEnable && (624 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_4_io_in_control_0_shift_b <=( _mesh_5_4_io_out_control_0_shift) ^ ((fiEnable && (625 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_4_io_in_control_0_dataflow_b <=( _mesh_5_4_io_out_control_0_dataflow) ^ ((fiEnable && (626 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_4_io_in_control_0_propagate_b <=( _mesh_5_4_io_out_control_0_propagate) ^ ((fiEnable && (627 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_4_io_out_valid_0) begin
			b_71_0 <=( _mesh_6_4_io_out_b_0) ^ ((fiEnable && (628 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_327_0 <=( _mesh_6_4_io_out_c_0) ^ ((fiEnable && (629 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_4_io_in_control_0_shift_b <=( _mesh_6_4_io_out_control_0_shift) ^ ((fiEnable && (630 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_4_io_in_control_0_dataflow_b <=( _mesh_6_4_io_out_control_0_dataflow) ^ ((fiEnable && (631 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_4_io_in_control_0_propagate_b <=( _mesh_6_4_io_out_control_0_propagate) ^ ((fiEnable && (632 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_4_io_out_valid_0) begin
			b_72_0 <=( _mesh_7_4_io_out_b_0) ^ ((fiEnable && (633 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_328_0 <=( _mesh_7_4_io_out_c_0) ^ ((fiEnable && (634 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_4_io_in_control_0_shift_b <=( _mesh_7_4_io_out_control_0_shift) ^ ((fiEnable && (635 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_4_io_in_control_0_dataflow_b <=( _mesh_7_4_io_out_control_0_dataflow) ^ ((fiEnable && (636 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_4_io_in_control_0_propagate_b <=( _mesh_7_4_io_out_control_0_propagate) ^ ((fiEnable && (637 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_4_io_out_valid_0) begin
			b_73_0 <=( _mesh_8_4_io_out_b_0) ^ ((fiEnable && (638 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_329_0 <=( _mesh_8_4_io_out_c_0) ^ ((fiEnable && (639 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_4_io_in_control_0_shift_b <=( _mesh_8_4_io_out_control_0_shift) ^ ((fiEnable && (640 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_4_io_in_control_0_dataflow_b <=( _mesh_8_4_io_out_control_0_dataflow) ^ ((fiEnable && (641 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_4_io_in_control_0_propagate_b <=( _mesh_8_4_io_out_control_0_propagate) ^ ((fiEnable && (642 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_4_io_out_valid_0) begin
			b_74_0 <=( _mesh_9_4_io_out_b_0) ^ ((fiEnable && (643 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_330_0 <=( _mesh_9_4_io_out_c_0) ^ ((fiEnable && (644 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_4_io_in_control_0_shift_b <=( _mesh_9_4_io_out_control_0_shift) ^ ((fiEnable && (645 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_4_io_in_control_0_dataflow_b <=( _mesh_9_4_io_out_control_0_dataflow) ^ ((fiEnable && (646 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_4_io_in_control_0_propagate_b <=( _mesh_9_4_io_out_control_0_propagate) ^ ((fiEnable && (647 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_4_io_out_valid_0) begin
			b_75_0 <=( _mesh_10_4_io_out_b_0) ^ ((fiEnable && (648 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_331_0 <=( _mesh_10_4_io_out_c_0) ^ ((fiEnable && (649 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_4_io_in_control_0_shift_b <=( _mesh_10_4_io_out_control_0_shift) ^ ((fiEnable && (650 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_4_io_in_control_0_dataflow_b <=( _mesh_10_4_io_out_control_0_dataflow) ^ ((fiEnable && (651 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_4_io_in_control_0_propagate_b <=( _mesh_10_4_io_out_control_0_propagate) ^ ((fiEnable && (652 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_4_io_out_valid_0) begin
			b_76_0 <=( _mesh_11_4_io_out_b_0) ^ ((fiEnable && (653 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_332_0 <=( _mesh_11_4_io_out_c_0) ^ ((fiEnable && (654 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_4_io_in_control_0_shift_b <=( _mesh_11_4_io_out_control_0_shift) ^ ((fiEnable && (655 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_4_io_in_control_0_dataflow_b <=( _mesh_11_4_io_out_control_0_dataflow) ^ ((fiEnable && (656 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_4_io_in_control_0_propagate_b <=( _mesh_11_4_io_out_control_0_propagate) ^ ((fiEnable && (657 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_4_io_out_valid_0) begin
			b_77_0 <=( _mesh_12_4_io_out_b_0) ^ ((fiEnable && (658 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_333_0 <=( _mesh_12_4_io_out_c_0) ^ ((fiEnable && (659 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_4_io_in_control_0_shift_b <=( _mesh_12_4_io_out_control_0_shift) ^ ((fiEnable && (660 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_4_io_in_control_0_dataflow_b <=( _mesh_12_4_io_out_control_0_dataflow) ^ ((fiEnable && (661 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_4_io_in_control_0_propagate_b <=( _mesh_12_4_io_out_control_0_propagate) ^ ((fiEnable && (662 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_4_io_out_valid_0) begin
			b_78_0 <=( _mesh_13_4_io_out_b_0) ^ ((fiEnable && (663 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_334_0 <=( _mesh_13_4_io_out_c_0) ^ ((fiEnable && (664 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_4_io_in_control_0_shift_b <=( _mesh_13_4_io_out_control_0_shift) ^ ((fiEnable && (665 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_4_io_in_control_0_dataflow_b <=( _mesh_13_4_io_out_control_0_dataflow) ^ ((fiEnable && (666 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_4_io_in_control_0_propagate_b <=( _mesh_13_4_io_out_control_0_propagate) ^ ((fiEnable && (667 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_4_io_out_valid_0) begin
			b_79_0 <=( _mesh_14_4_io_out_b_0) ^ ((fiEnable && (668 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_335_0 <=( _mesh_14_4_io_out_c_0) ^ ((fiEnable && (669 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_4_io_in_control_0_shift_b <=( _mesh_14_4_io_out_control_0_shift) ^ ((fiEnable && (670 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_4_io_in_control_0_dataflow_b <=( _mesh_14_4_io_out_control_0_dataflow) ^ ((fiEnable && (671 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_4_io_in_control_0_propagate_b <=( _mesh_14_4_io_out_control_0_propagate) ^ ((fiEnable && (672 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_5_0) begin
			b_80_0 <=( io_in_b_5_0) ^ ((fiEnable && (673 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_336_0 <=( io_in_d_5_0) ^ ((fiEnable && (674 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_5_io_in_control_0_shift_b <=( io_in_control_5_0_shift) ^ ((fiEnable && (675 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_5_io_in_control_0_dataflow_b <=( io_in_control_5_0_dataflow) ^ ((fiEnable && (676 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_5_io_in_control_0_propagate_b <=( io_in_control_5_0_propagate) ^ ((fiEnable && (677 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_5_io_out_valid_0) begin
			b_81_0 <=( _mesh_0_5_io_out_b_0) ^ ((fiEnable && (678 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_337_0 <=( _mesh_0_5_io_out_c_0) ^ ((fiEnable && (679 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_5_io_in_control_0_shift_b <=( _mesh_0_5_io_out_control_0_shift) ^ ((fiEnable && (680 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_5_io_in_control_0_dataflow_b <=( _mesh_0_5_io_out_control_0_dataflow) ^ ((fiEnable && (681 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_5_io_in_control_0_propagate_b <=( _mesh_0_5_io_out_control_0_propagate) ^ ((fiEnable && (682 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_5_io_out_valid_0) begin
			b_82_0 <=( _mesh_1_5_io_out_b_0) ^ ((fiEnable && (683 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_338_0 <=( _mesh_1_5_io_out_c_0) ^ ((fiEnable && (684 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_5_io_in_control_0_shift_b <=( _mesh_1_5_io_out_control_0_shift) ^ ((fiEnable && (685 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_5_io_in_control_0_dataflow_b <=( _mesh_1_5_io_out_control_0_dataflow) ^ ((fiEnable && (686 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_5_io_in_control_0_propagate_b <=( _mesh_1_5_io_out_control_0_propagate) ^ ((fiEnable && (687 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_5_io_out_valid_0) begin
			b_83_0 <=( _mesh_2_5_io_out_b_0) ^ ((fiEnable && (688 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_339_0 <=( _mesh_2_5_io_out_c_0) ^ ((fiEnable && (689 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_5_io_in_control_0_shift_b <=( _mesh_2_5_io_out_control_0_shift) ^ ((fiEnable && (690 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_5_io_in_control_0_dataflow_b <=( _mesh_2_5_io_out_control_0_dataflow) ^ ((fiEnable && (691 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_5_io_in_control_0_propagate_b <=( _mesh_2_5_io_out_control_0_propagate) ^ ((fiEnable && (692 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_5_io_out_valid_0) begin
			b_84_0 <=( _mesh_3_5_io_out_b_0) ^ ((fiEnable && (693 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_340_0 <=( _mesh_3_5_io_out_c_0) ^ ((fiEnable && (694 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_5_io_in_control_0_shift_b <=( _mesh_3_5_io_out_control_0_shift) ^ ((fiEnable && (695 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_5_io_in_control_0_dataflow_b <=( _mesh_3_5_io_out_control_0_dataflow) ^ ((fiEnable && (696 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_5_io_in_control_0_propagate_b <=( _mesh_3_5_io_out_control_0_propagate) ^ ((fiEnable && (697 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_5_io_out_valid_0) begin
			b_85_0 <=( _mesh_4_5_io_out_b_0) ^ ((fiEnable && (698 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_341_0 <=( _mesh_4_5_io_out_c_0) ^ ((fiEnable && (699 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_5_io_in_control_0_shift_b <=( _mesh_4_5_io_out_control_0_shift) ^ ((fiEnable && (700 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_5_io_in_control_0_dataflow_b <=( _mesh_4_5_io_out_control_0_dataflow) ^ ((fiEnable && (701 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_5_io_in_control_0_propagate_b <=( _mesh_4_5_io_out_control_0_propagate) ^ ((fiEnable && (702 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_5_io_out_valid_0) begin
			b_86_0 <=( _mesh_5_5_io_out_b_0) ^ ((fiEnable && (703 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_342_0 <=( _mesh_5_5_io_out_c_0) ^ ((fiEnable && (704 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_5_io_in_control_0_shift_b <=( _mesh_5_5_io_out_control_0_shift) ^ ((fiEnable && (705 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_5_io_in_control_0_dataflow_b <=( _mesh_5_5_io_out_control_0_dataflow) ^ ((fiEnable && (706 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_5_io_in_control_0_propagate_b <=( _mesh_5_5_io_out_control_0_propagate) ^ ((fiEnable && (707 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_5_io_out_valid_0) begin
			b_87_0 <=( _mesh_6_5_io_out_b_0) ^ ((fiEnable && (708 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_343_0 <=( _mesh_6_5_io_out_c_0) ^ ((fiEnable && (709 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_5_io_in_control_0_shift_b <=( _mesh_6_5_io_out_control_0_shift) ^ ((fiEnable && (710 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_5_io_in_control_0_dataflow_b <=( _mesh_6_5_io_out_control_0_dataflow) ^ ((fiEnable && (711 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_5_io_in_control_0_propagate_b <=( _mesh_6_5_io_out_control_0_propagate) ^ ((fiEnable && (712 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_5_io_out_valid_0) begin
			b_88_0 <=( _mesh_7_5_io_out_b_0) ^ ((fiEnable && (713 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_344_0 <=( _mesh_7_5_io_out_c_0) ^ ((fiEnable && (714 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_5_io_in_control_0_shift_b <=( _mesh_7_5_io_out_control_0_shift) ^ ((fiEnable && (715 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_5_io_in_control_0_dataflow_b <=( _mesh_7_5_io_out_control_0_dataflow) ^ ((fiEnable && (716 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_5_io_in_control_0_propagate_b <=( _mesh_7_5_io_out_control_0_propagate) ^ ((fiEnable && (717 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_5_io_out_valid_0) begin
			b_89_0 <=( _mesh_8_5_io_out_b_0) ^ ((fiEnable && (718 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_345_0 <=( _mesh_8_5_io_out_c_0) ^ ((fiEnable && (719 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_5_io_in_control_0_shift_b <=( _mesh_8_5_io_out_control_0_shift) ^ ((fiEnable && (720 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_5_io_in_control_0_dataflow_b <=( _mesh_8_5_io_out_control_0_dataflow) ^ ((fiEnable && (721 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_5_io_in_control_0_propagate_b <=( _mesh_8_5_io_out_control_0_propagate) ^ ((fiEnable && (722 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_5_io_out_valid_0) begin
			b_90_0 <=( _mesh_9_5_io_out_b_0) ^ ((fiEnable && (723 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_346_0 <=( _mesh_9_5_io_out_c_0) ^ ((fiEnable && (724 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_5_io_in_control_0_shift_b <=( _mesh_9_5_io_out_control_0_shift) ^ ((fiEnable && (725 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_5_io_in_control_0_dataflow_b <=( _mesh_9_5_io_out_control_0_dataflow) ^ ((fiEnable && (726 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_5_io_in_control_0_propagate_b <=( _mesh_9_5_io_out_control_0_propagate) ^ ((fiEnable && (727 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_5_io_out_valid_0) begin
			b_91_0 <=( _mesh_10_5_io_out_b_0) ^ ((fiEnable && (728 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_347_0 <=( _mesh_10_5_io_out_c_0) ^ ((fiEnable && (729 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_5_io_in_control_0_shift_b <=( _mesh_10_5_io_out_control_0_shift) ^ ((fiEnable && (730 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_5_io_in_control_0_dataflow_b <=( _mesh_10_5_io_out_control_0_dataflow) ^ ((fiEnable && (731 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_5_io_in_control_0_propagate_b <=( _mesh_10_5_io_out_control_0_propagate) ^ ((fiEnable && (732 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_5_io_out_valid_0) begin
			b_92_0 <=( _mesh_11_5_io_out_b_0) ^ ((fiEnable && (733 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_348_0 <=( _mesh_11_5_io_out_c_0) ^ ((fiEnable && (734 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_5_io_in_control_0_shift_b <=( _mesh_11_5_io_out_control_0_shift) ^ ((fiEnable && (735 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_5_io_in_control_0_dataflow_b <=( _mesh_11_5_io_out_control_0_dataflow) ^ ((fiEnable && (736 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_5_io_in_control_0_propagate_b <=( _mesh_11_5_io_out_control_0_propagate) ^ ((fiEnable && (737 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_5_io_out_valid_0) begin
			b_93_0 <=( _mesh_12_5_io_out_b_0) ^ ((fiEnable && (738 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_349_0 <=( _mesh_12_5_io_out_c_0) ^ ((fiEnable && (739 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_5_io_in_control_0_shift_b <=( _mesh_12_5_io_out_control_0_shift) ^ ((fiEnable && (740 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_5_io_in_control_0_dataflow_b <=( _mesh_12_5_io_out_control_0_dataflow) ^ ((fiEnable && (741 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_5_io_in_control_0_propagate_b <=( _mesh_12_5_io_out_control_0_propagate) ^ ((fiEnable && (742 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_5_io_out_valid_0) begin
			b_94_0 <=( _mesh_13_5_io_out_b_0) ^ ((fiEnable && (743 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_350_0 <=( _mesh_13_5_io_out_c_0) ^ ((fiEnable && (744 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_5_io_in_control_0_shift_b <=( _mesh_13_5_io_out_control_0_shift) ^ ((fiEnable && (745 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_5_io_in_control_0_dataflow_b <=( _mesh_13_5_io_out_control_0_dataflow) ^ ((fiEnable && (746 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_5_io_in_control_0_propagate_b <=( _mesh_13_5_io_out_control_0_propagate) ^ ((fiEnable && (747 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_5_io_out_valid_0) begin
			b_95_0 <=( _mesh_14_5_io_out_b_0) ^ ((fiEnable && (748 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_351_0 <=( _mesh_14_5_io_out_c_0) ^ ((fiEnable && (749 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_5_io_in_control_0_shift_b <=( _mesh_14_5_io_out_control_0_shift) ^ ((fiEnable && (750 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_5_io_in_control_0_dataflow_b <=( _mesh_14_5_io_out_control_0_dataflow) ^ ((fiEnable && (751 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_5_io_in_control_0_propagate_b <=( _mesh_14_5_io_out_control_0_propagate) ^ ((fiEnable && (752 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_6_0) begin
			b_96_0 <=( io_in_b_6_0) ^ ((fiEnable && (753 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_352_0 <=( io_in_d_6_0) ^ ((fiEnable && (754 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_6_io_in_control_0_shift_b <=( io_in_control_6_0_shift) ^ ((fiEnable && (755 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_6_io_in_control_0_dataflow_b <=( io_in_control_6_0_dataflow) ^ ((fiEnable && (756 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_6_io_in_control_0_propagate_b <=( io_in_control_6_0_propagate) ^ ((fiEnable && (757 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_6_io_out_valid_0) begin
			b_97_0 <=( _mesh_0_6_io_out_b_0) ^ ((fiEnable && (758 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_353_0 <=( _mesh_0_6_io_out_c_0) ^ ((fiEnable && (759 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_6_io_in_control_0_shift_b <=( _mesh_0_6_io_out_control_0_shift) ^ ((fiEnable && (760 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_6_io_in_control_0_dataflow_b <=( _mesh_0_6_io_out_control_0_dataflow) ^ ((fiEnable && (761 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_6_io_in_control_0_propagate_b <=( _mesh_0_6_io_out_control_0_propagate) ^ ((fiEnable && (762 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_6_io_out_valid_0) begin
			b_98_0 <=( _mesh_1_6_io_out_b_0) ^ ((fiEnable && (763 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_354_0 <=( _mesh_1_6_io_out_c_0) ^ ((fiEnable && (764 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_6_io_in_control_0_shift_b <=( _mesh_1_6_io_out_control_0_shift) ^ ((fiEnable && (765 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_6_io_in_control_0_dataflow_b <=( _mesh_1_6_io_out_control_0_dataflow) ^ ((fiEnable && (766 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_6_io_in_control_0_propagate_b <=( _mesh_1_6_io_out_control_0_propagate) ^ ((fiEnable && (767 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_6_io_out_valid_0) begin
			b_99_0 <=( _mesh_2_6_io_out_b_0) ^ ((fiEnable && (768 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_355_0 <=( _mesh_2_6_io_out_c_0) ^ ((fiEnable && (769 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_6_io_in_control_0_shift_b <=( _mesh_2_6_io_out_control_0_shift) ^ ((fiEnable && (770 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_6_io_in_control_0_dataflow_b <=( _mesh_2_6_io_out_control_0_dataflow) ^ ((fiEnable && (771 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_6_io_in_control_0_propagate_b <=( _mesh_2_6_io_out_control_0_propagate) ^ ((fiEnable && (772 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_6_io_out_valid_0) begin
			b_100_0 <=( _mesh_3_6_io_out_b_0) ^ ((fiEnable && (773 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_356_0 <=( _mesh_3_6_io_out_c_0) ^ ((fiEnable && (774 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_6_io_in_control_0_shift_b <=( _mesh_3_6_io_out_control_0_shift) ^ ((fiEnable && (775 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_6_io_in_control_0_dataflow_b <=( _mesh_3_6_io_out_control_0_dataflow) ^ ((fiEnable && (776 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_6_io_in_control_0_propagate_b <=( _mesh_3_6_io_out_control_0_propagate) ^ ((fiEnable && (777 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_6_io_out_valid_0) begin
			b_101_0 <=( _mesh_4_6_io_out_b_0) ^ ((fiEnable && (778 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_357_0 <=( _mesh_4_6_io_out_c_0) ^ ((fiEnable && (779 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_6_io_in_control_0_shift_b <=( _mesh_4_6_io_out_control_0_shift) ^ ((fiEnable && (780 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_6_io_in_control_0_dataflow_b <=( _mesh_4_6_io_out_control_0_dataflow) ^ ((fiEnable && (781 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_6_io_in_control_0_propagate_b <=( _mesh_4_6_io_out_control_0_propagate) ^ ((fiEnable && (782 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_6_io_out_valid_0) begin
			b_102_0 <=( _mesh_5_6_io_out_b_0) ^ ((fiEnable && (783 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_358_0 <=( _mesh_5_6_io_out_c_0) ^ ((fiEnable && (784 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_6_io_in_control_0_shift_b <=( _mesh_5_6_io_out_control_0_shift) ^ ((fiEnable && (785 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_6_io_in_control_0_dataflow_b <=( _mesh_5_6_io_out_control_0_dataflow) ^ ((fiEnable && (786 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_6_io_in_control_0_propagate_b <=( _mesh_5_6_io_out_control_0_propagate) ^ ((fiEnable && (787 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_6_io_out_valid_0) begin
			b_103_0 <=( _mesh_6_6_io_out_b_0) ^ ((fiEnable && (788 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_359_0 <=( _mesh_6_6_io_out_c_0) ^ ((fiEnable && (789 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_6_io_in_control_0_shift_b <=( _mesh_6_6_io_out_control_0_shift) ^ ((fiEnable && (790 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_6_io_in_control_0_dataflow_b <=( _mesh_6_6_io_out_control_0_dataflow) ^ ((fiEnable && (791 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_6_io_in_control_0_propagate_b <=( _mesh_6_6_io_out_control_0_propagate) ^ ((fiEnable && (792 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_6_io_out_valid_0) begin
			b_104_0 <=( _mesh_7_6_io_out_b_0) ^ ((fiEnable && (793 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_360_0 <=( _mesh_7_6_io_out_c_0) ^ ((fiEnable && (794 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_6_io_in_control_0_shift_b <=( _mesh_7_6_io_out_control_0_shift) ^ ((fiEnable && (795 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_6_io_in_control_0_dataflow_b <=( _mesh_7_6_io_out_control_0_dataflow) ^ ((fiEnable && (796 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_6_io_in_control_0_propagate_b <=( _mesh_7_6_io_out_control_0_propagate) ^ ((fiEnable && (797 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_6_io_out_valid_0) begin
			b_105_0 <=( _mesh_8_6_io_out_b_0) ^ ((fiEnable && (798 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_361_0 <=( _mesh_8_6_io_out_c_0) ^ ((fiEnable && (799 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_6_io_in_control_0_shift_b <=( _mesh_8_6_io_out_control_0_shift) ^ ((fiEnable && (800 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_6_io_in_control_0_dataflow_b <=( _mesh_8_6_io_out_control_0_dataflow) ^ ((fiEnable && (801 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_6_io_in_control_0_propagate_b <=( _mesh_8_6_io_out_control_0_propagate) ^ ((fiEnable && (802 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_6_io_out_valid_0) begin
			b_106_0 <=( _mesh_9_6_io_out_b_0) ^ ((fiEnable && (803 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_362_0 <=( _mesh_9_6_io_out_c_0) ^ ((fiEnable && (804 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_6_io_in_control_0_shift_b <=( _mesh_9_6_io_out_control_0_shift) ^ ((fiEnable && (805 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_6_io_in_control_0_dataflow_b <=( _mesh_9_6_io_out_control_0_dataflow) ^ ((fiEnable && (806 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_6_io_in_control_0_propagate_b <=( _mesh_9_6_io_out_control_0_propagate) ^ ((fiEnable && (807 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_6_io_out_valid_0) begin
			b_107_0 <=( _mesh_10_6_io_out_b_0) ^ ((fiEnable && (808 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_363_0 <=( _mesh_10_6_io_out_c_0) ^ ((fiEnable && (809 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_6_io_in_control_0_shift_b <=( _mesh_10_6_io_out_control_0_shift) ^ ((fiEnable && (810 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_6_io_in_control_0_dataflow_b <=( _mesh_10_6_io_out_control_0_dataflow) ^ ((fiEnable && (811 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_6_io_in_control_0_propagate_b <=( _mesh_10_6_io_out_control_0_propagate) ^ ((fiEnable && (812 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_6_io_out_valid_0) begin
			b_108_0 <=( _mesh_11_6_io_out_b_0) ^ ((fiEnable && (813 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_364_0 <=( _mesh_11_6_io_out_c_0) ^ ((fiEnable && (814 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_6_io_in_control_0_shift_b <=( _mesh_11_6_io_out_control_0_shift) ^ ((fiEnable && (815 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_6_io_in_control_0_dataflow_b <=( _mesh_11_6_io_out_control_0_dataflow) ^ ((fiEnable && (816 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_6_io_in_control_0_propagate_b <=( _mesh_11_6_io_out_control_0_propagate) ^ ((fiEnable && (817 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_6_io_out_valid_0) begin
			b_109_0 <=( _mesh_12_6_io_out_b_0) ^ ((fiEnable && (818 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_365_0 <=( _mesh_12_6_io_out_c_0) ^ ((fiEnable && (819 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_6_io_in_control_0_shift_b <=( _mesh_12_6_io_out_control_0_shift) ^ ((fiEnable && (820 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_6_io_in_control_0_dataflow_b <=( _mesh_12_6_io_out_control_0_dataflow) ^ ((fiEnable && (821 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_6_io_in_control_0_propagate_b <=( _mesh_12_6_io_out_control_0_propagate) ^ ((fiEnable && (822 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_6_io_out_valid_0) begin
			b_110_0 <=( _mesh_13_6_io_out_b_0) ^ ((fiEnable && (823 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_366_0 <=( _mesh_13_6_io_out_c_0) ^ ((fiEnable && (824 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_6_io_in_control_0_shift_b <=( _mesh_13_6_io_out_control_0_shift) ^ ((fiEnable && (825 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_6_io_in_control_0_dataflow_b <=( _mesh_13_6_io_out_control_0_dataflow) ^ ((fiEnable && (826 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_6_io_in_control_0_propagate_b <=( _mesh_13_6_io_out_control_0_propagate) ^ ((fiEnable && (827 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_6_io_out_valid_0) begin
			b_111_0 <=( _mesh_14_6_io_out_b_0) ^ ((fiEnable && (828 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_367_0 <=( _mesh_14_6_io_out_c_0) ^ ((fiEnable && (829 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_6_io_in_control_0_shift_b <=( _mesh_14_6_io_out_control_0_shift) ^ ((fiEnable && (830 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_6_io_in_control_0_dataflow_b <=( _mesh_14_6_io_out_control_0_dataflow) ^ ((fiEnable && (831 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_6_io_in_control_0_propagate_b <=( _mesh_14_6_io_out_control_0_propagate) ^ ((fiEnable && (832 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_7_0) begin
			b_112_0 <=( io_in_b_7_0) ^ ((fiEnable && (833 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_368_0 <=( io_in_d_7_0) ^ ((fiEnable && (834 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_7_io_in_control_0_shift_b <=( io_in_control_7_0_shift) ^ ((fiEnable && (835 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_7_io_in_control_0_dataflow_b <=( io_in_control_7_0_dataflow) ^ ((fiEnable && (836 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_7_io_in_control_0_propagate_b <=( io_in_control_7_0_propagate) ^ ((fiEnable && (837 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_7_io_out_valid_0) begin
			b_113_0 <=( _mesh_0_7_io_out_b_0) ^ ((fiEnable && (838 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_369_0 <=( _mesh_0_7_io_out_c_0) ^ ((fiEnable && (839 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_7_io_in_control_0_shift_b <=( _mesh_0_7_io_out_control_0_shift) ^ ((fiEnable && (840 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_7_io_in_control_0_dataflow_b <=( _mesh_0_7_io_out_control_0_dataflow) ^ ((fiEnable && (841 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_7_io_in_control_0_propagate_b <=( _mesh_0_7_io_out_control_0_propagate) ^ ((fiEnable && (842 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_7_io_out_valid_0) begin
			b_114_0 <=( _mesh_1_7_io_out_b_0) ^ ((fiEnable && (843 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_370_0 <=( _mesh_1_7_io_out_c_0) ^ ((fiEnable && (844 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_7_io_in_control_0_shift_b <=( _mesh_1_7_io_out_control_0_shift) ^ ((fiEnable && (845 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_7_io_in_control_0_dataflow_b <=( _mesh_1_7_io_out_control_0_dataflow) ^ ((fiEnable && (846 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_7_io_in_control_0_propagate_b <=( _mesh_1_7_io_out_control_0_propagate) ^ ((fiEnable && (847 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_7_io_out_valid_0) begin
			b_115_0 <=( _mesh_2_7_io_out_b_0) ^ ((fiEnable && (848 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_371_0 <=( _mesh_2_7_io_out_c_0) ^ ((fiEnable && (849 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_7_io_in_control_0_shift_b <=( _mesh_2_7_io_out_control_0_shift) ^ ((fiEnable && (850 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_7_io_in_control_0_dataflow_b <=( _mesh_2_7_io_out_control_0_dataflow) ^ ((fiEnable && (851 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_7_io_in_control_0_propagate_b <=( _mesh_2_7_io_out_control_0_propagate) ^ ((fiEnable && (852 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_7_io_out_valid_0) begin
			b_116_0 <=( _mesh_3_7_io_out_b_0) ^ ((fiEnable && (853 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_372_0 <=( _mesh_3_7_io_out_c_0) ^ ((fiEnable && (854 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_7_io_in_control_0_shift_b <=( _mesh_3_7_io_out_control_0_shift) ^ ((fiEnable && (855 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_7_io_in_control_0_dataflow_b <=( _mesh_3_7_io_out_control_0_dataflow) ^ ((fiEnable && (856 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_7_io_in_control_0_propagate_b <=( _mesh_3_7_io_out_control_0_propagate) ^ ((fiEnable && (857 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_7_io_out_valid_0) begin
			b_117_0 <=( _mesh_4_7_io_out_b_0) ^ ((fiEnable && (858 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_373_0 <=( _mesh_4_7_io_out_c_0) ^ ((fiEnable && (859 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_7_io_in_control_0_shift_b <=( _mesh_4_7_io_out_control_0_shift) ^ ((fiEnable && (860 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_7_io_in_control_0_dataflow_b <=( _mesh_4_7_io_out_control_0_dataflow) ^ ((fiEnable && (861 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_7_io_in_control_0_propagate_b <=( _mesh_4_7_io_out_control_0_propagate) ^ ((fiEnable && (862 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_7_io_out_valid_0) begin
			b_118_0 <=( _mesh_5_7_io_out_b_0) ^ ((fiEnable && (863 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_374_0 <=( _mesh_5_7_io_out_c_0) ^ ((fiEnable && (864 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_7_io_in_control_0_shift_b <=( _mesh_5_7_io_out_control_0_shift) ^ ((fiEnable && (865 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_7_io_in_control_0_dataflow_b <=( _mesh_5_7_io_out_control_0_dataflow) ^ ((fiEnable && (866 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_7_io_in_control_0_propagate_b <=( _mesh_5_7_io_out_control_0_propagate) ^ ((fiEnable && (867 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_7_io_out_valid_0) begin
			b_119_0 <=( _mesh_6_7_io_out_b_0) ^ ((fiEnable && (868 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_375_0 <=( _mesh_6_7_io_out_c_0) ^ ((fiEnable && (869 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_7_io_in_control_0_shift_b <=( _mesh_6_7_io_out_control_0_shift) ^ ((fiEnable && (870 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_7_io_in_control_0_dataflow_b <=( _mesh_6_7_io_out_control_0_dataflow) ^ ((fiEnable && (871 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_7_io_in_control_0_propagate_b <=( _mesh_6_7_io_out_control_0_propagate) ^ ((fiEnable && (872 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_7_io_out_valid_0) begin
			b_120_0 <=( _mesh_7_7_io_out_b_0) ^ ((fiEnable && (873 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_376_0 <=( _mesh_7_7_io_out_c_0) ^ ((fiEnable && (874 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_7_io_in_control_0_shift_b <=( _mesh_7_7_io_out_control_0_shift) ^ ((fiEnable && (875 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_7_io_in_control_0_dataflow_b <=( _mesh_7_7_io_out_control_0_dataflow) ^ ((fiEnable && (876 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_7_io_in_control_0_propagate_b <=( _mesh_7_7_io_out_control_0_propagate) ^ ((fiEnable && (877 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_7_io_out_valid_0) begin
			b_121_0 <=( _mesh_8_7_io_out_b_0) ^ ((fiEnable && (878 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_377_0 <=( _mesh_8_7_io_out_c_0) ^ ((fiEnable && (879 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_7_io_in_control_0_shift_b <=( _mesh_8_7_io_out_control_0_shift) ^ ((fiEnable && (880 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_7_io_in_control_0_dataflow_b <=( _mesh_8_7_io_out_control_0_dataflow) ^ ((fiEnable && (881 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_7_io_in_control_0_propagate_b <=( _mesh_8_7_io_out_control_0_propagate) ^ ((fiEnable && (882 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_7_io_out_valid_0) begin
			b_122_0 <=( _mesh_9_7_io_out_b_0) ^ ((fiEnable && (883 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_378_0 <=( _mesh_9_7_io_out_c_0) ^ ((fiEnable && (884 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_7_io_in_control_0_shift_b <=( _mesh_9_7_io_out_control_0_shift) ^ ((fiEnable && (885 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_7_io_in_control_0_dataflow_b <=( _mesh_9_7_io_out_control_0_dataflow) ^ ((fiEnable && (886 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_7_io_in_control_0_propagate_b <=( _mesh_9_7_io_out_control_0_propagate) ^ ((fiEnable && (887 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_7_io_out_valid_0) begin
			b_123_0 <=( _mesh_10_7_io_out_b_0) ^ ((fiEnable && (888 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_379_0 <=( _mesh_10_7_io_out_c_0) ^ ((fiEnable && (889 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_7_io_in_control_0_shift_b <=( _mesh_10_7_io_out_control_0_shift) ^ ((fiEnable && (890 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_7_io_in_control_0_dataflow_b <=( _mesh_10_7_io_out_control_0_dataflow) ^ ((fiEnable && (891 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_7_io_in_control_0_propagate_b <=( _mesh_10_7_io_out_control_0_propagate) ^ ((fiEnable && (892 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_7_io_out_valid_0) begin
			b_124_0 <=( _mesh_11_7_io_out_b_0) ^ ((fiEnable && (893 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_380_0 <=( _mesh_11_7_io_out_c_0) ^ ((fiEnable && (894 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_7_io_in_control_0_shift_b <=( _mesh_11_7_io_out_control_0_shift) ^ ((fiEnable && (895 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_7_io_in_control_0_dataflow_b <=( _mesh_11_7_io_out_control_0_dataflow) ^ ((fiEnable && (896 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_7_io_in_control_0_propagate_b <=( _mesh_11_7_io_out_control_0_propagate) ^ ((fiEnable && (897 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_7_io_out_valid_0) begin
			b_125_0 <=( _mesh_12_7_io_out_b_0) ^ ((fiEnable && (898 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_381_0 <=( _mesh_12_7_io_out_c_0) ^ ((fiEnable && (899 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_7_io_in_control_0_shift_b <=( _mesh_12_7_io_out_control_0_shift) ^ ((fiEnable && (900 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_7_io_in_control_0_dataflow_b <=( _mesh_12_7_io_out_control_0_dataflow) ^ ((fiEnable && (901 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_7_io_in_control_0_propagate_b <=( _mesh_12_7_io_out_control_0_propagate) ^ ((fiEnable && (902 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_7_io_out_valid_0) begin
			b_126_0 <=( _mesh_13_7_io_out_b_0) ^ ((fiEnable && (903 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_382_0 <=( _mesh_13_7_io_out_c_0) ^ ((fiEnable && (904 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_7_io_in_control_0_shift_b <=( _mesh_13_7_io_out_control_0_shift) ^ ((fiEnable && (905 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_7_io_in_control_0_dataflow_b <=( _mesh_13_7_io_out_control_0_dataflow) ^ ((fiEnable && (906 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_7_io_in_control_0_propagate_b <=( _mesh_13_7_io_out_control_0_propagate) ^ ((fiEnable && (907 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_7_io_out_valid_0) begin
			b_127_0 <=( _mesh_14_7_io_out_b_0) ^ ((fiEnable && (908 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_383_0 <=( _mesh_14_7_io_out_c_0) ^ ((fiEnable && (909 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_7_io_in_control_0_shift_b <=( _mesh_14_7_io_out_control_0_shift) ^ ((fiEnable && (910 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_7_io_in_control_0_dataflow_b <=( _mesh_14_7_io_out_control_0_dataflow) ^ ((fiEnable && (911 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_7_io_in_control_0_propagate_b <=( _mesh_14_7_io_out_control_0_propagate) ^ ((fiEnable && (912 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_8_0) begin
			b_128_0 <=( io_in_b_8_0) ^ ((fiEnable && (913 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_384_0 <=( io_in_d_8_0) ^ ((fiEnable && (914 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_8_io_in_control_0_shift_b <=( io_in_control_8_0_shift) ^ ((fiEnable && (915 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_8_io_in_control_0_dataflow_b <=( io_in_control_8_0_dataflow) ^ ((fiEnable && (916 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_8_io_in_control_0_propagate_b <=( io_in_control_8_0_propagate) ^ ((fiEnable && (917 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_8_io_out_valid_0) begin
			b_129_0 <=( _mesh_0_8_io_out_b_0) ^ ((fiEnable && (918 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_385_0 <=( _mesh_0_8_io_out_c_0) ^ ((fiEnable && (919 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_8_io_in_control_0_shift_b <=( _mesh_0_8_io_out_control_0_shift) ^ ((fiEnable && (920 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_8_io_in_control_0_dataflow_b <=( _mesh_0_8_io_out_control_0_dataflow) ^ ((fiEnable && (921 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_8_io_in_control_0_propagate_b <=( _mesh_0_8_io_out_control_0_propagate) ^ ((fiEnable && (922 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_8_io_out_valid_0) begin
			b_130_0 <=( _mesh_1_8_io_out_b_0) ^ ((fiEnable && (923 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_386_0 <=( _mesh_1_8_io_out_c_0) ^ ((fiEnable && (924 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_8_io_in_control_0_shift_b <=( _mesh_1_8_io_out_control_0_shift) ^ ((fiEnable && (925 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_8_io_in_control_0_dataflow_b <=( _mesh_1_8_io_out_control_0_dataflow) ^ ((fiEnable && (926 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_8_io_in_control_0_propagate_b <=( _mesh_1_8_io_out_control_0_propagate) ^ ((fiEnable && (927 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_8_io_out_valid_0) begin
			b_131_0 <=( _mesh_2_8_io_out_b_0) ^ ((fiEnable && (928 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_387_0 <=( _mesh_2_8_io_out_c_0) ^ ((fiEnable && (929 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_8_io_in_control_0_shift_b <=( _mesh_2_8_io_out_control_0_shift) ^ ((fiEnable && (930 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_8_io_in_control_0_dataflow_b <=( _mesh_2_8_io_out_control_0_dataflow) ^ ((fiEnable && (931 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_8_io_in_control_0_propagate_b <=( _mesh_2_8_io_out_control_0_propagate) ^ ((fiEnable && (932 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_8_io_out_valid_0) begin
			b_132_0 <=( _mesh_3_8_io_out_b_0) ^ ((fiEnable && (933 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_388_0 <=( _mesh_3_8_io_out_c_0) ^ ((fiEnable && (934 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_8_io_in_control_0_shift_b <=( _mesh_3_8_io_out_control_0_shift) ^ ((fiEnable && (935 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_8_io_in_control_0_dataflow_b <=( _mesh_3_8_io_out_control_0_dataflow) ^ ((fiEnable && (936 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_8_io_in_control_0_propagate_b <=( _mesh_3_8_io_out_control_0_propagate) ^ ((fiEnable && (937 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_8_io_out_valid_0) begin
			b_133_0 <=( _mesh_4_8_io_out_b_0) ^ ((fiEnable && (938 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_389_0 <=( _mesh_4_8_io_out_c_0) ^ ((fiEnable && (939 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_8_io_in_control_0_shift_b <=( _mesh_4_8_io_out_control_0_shift) ^ ((fiEnable && (940 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_8_io_in_control_0_dataflow_b <=( _mesh_4_8_io_out_control_0_dataflow) ^ ((fiEnable && (941 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_8_io_in_control_0_propagate_b <=( _mesh_4_8_io_out_control_0_propagate) ^ ((fiEnable && (942 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_8_io_out_valid_0) begin
			b_134_0 <=( _mesh_5_8_io_out_b_0) ^ ((fiEnable && (943 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_390_0 <=( _mesh_5_8_io_out_c_0) ^ ((fiEnable && (944 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_8_io_in_control_0_shift_b <=( _mesh_5_8_io_out_control_0_shift) ^ ((fiEnable && (945 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_8_io_in_control_0_dataflow_b <=( _mesh_5_8_io_out_control_0_dataflow) ^ ((fiEnable && (946 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_8_io_in_control_0_propagate_b <=( _mesh_5_8_io_out_control_0_propagate) ^ ((fiEnable && (947 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_8_io_out_valid_0) begin
			b_135_0 <=( _mesh_6_8_io_out_b_0) ^ ((fiEnable && (948 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_391_0 <=( _mesh_6_8_io_out_c_0) ^ ((fiEnable && (949 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_8_io_in_control_0_shift_b <=( _mesh_6_8_io_out_control_0_shift) ^ ((fiEnable && (950 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_8_io_in_control_0_dataflow_b <=( _mesh_6_8_io_out_control_0_dataflow) ^ ((fiEnable && (951 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_8_io_in_control_0_propagate_b <=( _mesh_6_8_io_out_control_0_propagate) ^ ((fiEnable && (952 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_8_io_out_valid_0) begin
			b_136_0 <=( _mesh_7_8_io_out_b_0) ^ ((fiEnable && (953 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_392_0 <=( _mesh_7_8_io_out_c_0) ^ ((fiEnable && (954 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_8_io_in_control_0_shift_b <=( _mesh_7_8_io_out_control_0_shift) ^ ((fiEnable && (955 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_8_io_in_control_0_dataflow_b <=( _mesh_7_8_io_out_control_0_dataflow) ^ ((fiEnable && (956 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_8_io_in_control_0_propagate_b <=( _mesh_7_8_io_out_control_0_propagate) ^ ((fiEnable && (957 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_8_io_out_valid_0) begin
			b_137_0 <=( _mesh_8_8_io_out_b_0) ^ ((fiEnable && (958 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_393_0 <=( _mesh_8_8_io_out_c_0) ^ ((fiEnable && (959 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_8_io_in_control_0_shift_b <=( _mesh_8_8_io_out_control_0_shift) ^ ((fiEnable && (960 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_8_io_in_control_0_dataflow_b <=( _mesh_8_8_io_out_control_0_dataflow) ^ ((fiEnable && (961 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_8_io_in_control_0_propagate_b <=( _mesh_8_8_io_out_control_0_propagate) ^ ((fiEnable && (962 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_8_io_out_valid_0) begin
			b_138_0 <=( _mesh_9_8_io_out_b_0) ^ ((fiEnable && (963 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_394_0 <=( _mesh_9_8_io_out_c_0) ^ ((fiEnable && (964 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_8_io_in_control_0_shift_b <=( _mesh_9_8_io_out_control_0_shift) ^ ((fiEnable && (965 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_8_io_in_control_0_dataflow_b <=( _mesh_9_8_io_out_control_0_dataflow) ^ ((fiEnable && (966 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_8_io_in_control_0_propagate_b <=( _mesh_9_8_io_out_control_0_propagate) ^ ((fiEnable && (967 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_8_io_out_valid_0) begin
			b_139_0 <=( _mesh_10_8_io_out_b_0) ^ ((fiEnable && (968 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_395_0 <=( _mesh_10_8_io_out_c_0) ^ ((fiEnable && (969 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_8_io_in_control_0_shift_b <=( _mesh_10_8_io_out_control_0_shift) ^ ((fiEnable && (970 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_8_io_in_control_0_dataflow_b <=( _mesh_10_8_io_out_control_0_dataflow) ^ ((fiEnable && (971 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_8_io_in_control_0_propagate_b <=( _mesh_10_8_io_out_control_0_propagate) ^ ((fiEnable && (972 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_8_io_out_valid_0) begin
			b_140_0 <=( _mesh_11_8_io_out_b_0) ^ ((fiEnable && (973 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_396_0 <=( _mesh_11_8_io_out_c_0) ^ ((fiEnable && (974 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_8_io_in_control_0_shift_b <=( _mesh_11_8_io_out_control_0_shift) ^ ((fiEnable && (975 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_8_io_in_control_0_dataflow_b <=( _mesh_11_8_io_out_control_0_dataflow) ^ ((fiEnable && (976 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_8_io_in_control_0_propagate_b <=( _mesh_11_8_io_out_control_0_propagate) ^ ((fiEnable && (977 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_8_io_out_valid_0) begin
			b_141_0 <=( _mesh_12_8_io_out_b_0) ^ ((fiEnable && (978 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_397_0 <=( _mesh_12_8_io_out_c_0) ^ ((fiEnable && (979 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_8_io_in_control_0_shift_b <=( _mesh_12_8_io_out_control_0_shift) ^ ((fiEnable && (980 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_8_io_in_control_0_dataflow_b <=( _mesh_12_8_io_out_control_0_dataflow) ^ ((fiEnable && (981 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_8_io_in_control_0_propagate_b <=( _mesh_12_8_io_out_control_0_propagate) ^ ((fiEnable && (982 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_8_io_out_valid_0) begin
			b_142_0 <=( _mesh_13_8_io_out_b_0) ^ ((fiEnable && (983 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_398_0 <=( _mesh_13_8_io_out_c_0) ^ ((fiEnable && (984 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_8_io_in_control_0_shift_b <=( _mesh_13_8_io_out_control_0_shift) ^ ((fiEnable && (985 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_8_io_in_control_0_dataflow_b <=( _mesh_13_8_io_out_control_0_dataflow) ^ ((fiEnable && (986 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_8_io_in_control_0_propagate_b <=( _mesh_13_8_io_out_control_0_propagate) ^ ((fiEnable && (987 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_8_io_out_valid_0) begin
			b_143_0 <=( _mesh_14_8_io_out_b_0) ^ ((fiEnable && (988 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_399_0 <=( _mesh_14_8_io_out_c_0) ^ ((fiEnable && (989 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_8_io_in_control_0_shift_b <=( _mesh_14_8_io_out_control_0_shift) ^ ((fiEnable && (990 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_8_io_in_control_0_dataflow_b <=( _mesh_14_8_io_out_control_0_dataflow) ^ ((fiEnable && (991 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_8_io_in_control_0_propagate_b <=( _mesh_14_8_io_out_control_0_propagate) ^ ((fiEnable && (992 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_9_0) begin
			b_144_0 <=( io_in_b_9_0) ^ ((fiEnable && (993 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_400_0 <=( io_in_d_9_0) ^ ((fiEnable && (994 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_9_io_in_control_0_shift_b <=( io_in_control_9_0_shift) ^ ((fiEnable && (995 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_9_io_in_control_0_dataflow_b <=( io_in_control_9_0_dataflow) ^ ((fiEnable && (996 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_9_io_in_control_0_propagate_b <=( io_in_control_9_0_propagate) ^ ((fiEnable && (997 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_9_io_out_valid_0) begin
			b_145_0 <=( _mesh_0_9_io_out_b_0) ^ ((fiEnable && (998 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_401_0 <=( _mesh_0_9_io_out_c_0) ^ ((fiEnable && (999 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_9_io_in_control_0_shift_b <=( _mesh_0_9_io_out_control_0_shift) ^ ((fiEnable && (1000 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_9_io_in_control_0_dataflow_b <=( _mesh_0_9_io_out_control_0_dataflow) ^ ((fiEnable && (1001 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_9_io_in_control_0_propagate_b <=( _mesh_0_9_io_out_control_0_propagate) ^ ((fiEnable && (1002 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_9_io_out_valid_0) begin
			b_146_0 <=( _mesh_1_9_io_out_b_0) ^ ((fiEnable && (1003 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_402_0 <=( _mesh_1_9_io_out_c_0) ^ ((fiEnable && (1004 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_9_io_in_control_0_shift_b <=( _mesh_1_9_io_out_control_0_shift) ^ ((fiEnable && (1005 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_9_io_in_control_0_dataflow_b <=( _mesh_1_9_io_out_control_0_dataflow) ^ ((fiEnable && (1006 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_9_io_in_control_0_propagate_b <=( _mesh_1_9_io_out_control_0_propagate) ^ ((fiEnable && (1007 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_9_io_out_valid_0) begin
			b_147_0 <=( _mesh_2_9_io_out_b_0) ^ ((fiEnable && (1008 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_403_0 <=( _mesh_2_9_io_out_c_0) ^ ((fiEnable && (1009 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_9_io_in_control_0_shift_b <=( _mesh_2_9_io_out_control_0_shift) ^ ((fiEnable && (1010 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_9_io_in_control_0_dataflow_b <=( _mesh_2_9_io_out_control_0_dataflow) ^ ((fiEnable && (1011 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_9_io_in_control_0_propagate_b <=( _mesh_2_9_io_out_control_0_propagate) ^ ((fiEnable && (1012 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_9_io_out_valid_0) begin
			b_148_0 <=( _mesh_3_9_io_out_b_0) ^ ((fiEnable && (1013 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_404_0 <=( _mesh_3_9_io_out_c_0) ^ ((fiEnable && (1014 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_9_io_in_control_0_shift_b <=( _mesh_3_9_io_out_control_0_shift) ^ ((fiEnable && (1015 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_9_io_in_control_0_dataflow_b <=( _mesh_3_9_io_out_control_0_dataflow) ^ ((fiEnable && (1016 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_9_io_in_control_0_propagate_b <=( _mesh_3_9_io_out_control_0_propagate) ^ ((fiEnable && (1017 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_9_io_out_valid_0) begin
			b_149_0 <=( _mesh_4_9_io_out_b_0) ^ ((fiEnable && (1018 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_405_0 <=( _mesh_4_9_io_out_c_0) ^ ((fiEnable && (1019 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_9_io_in_control_0_shift_b <=( _mesh_4_9_io_out_control_0_shift) ^ ((fiEnable && (1020 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_9_io_in_control_0_dataflow_b <=( _mesh_4_9_io_out_control_0_dataflow) ^ ((fiEnable && (1021 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_9_io_in_control_0_propagate_b <=( _mesh_4_9_io_out_control_0_propagate) ^ ((fiEnable && (1022 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_9_io_out_valid_0) begin
			b_150_0 <=( _mesh_5_9_io_out_b_0) ^ ((fiEnable && (1023 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_406_0 <=( _mesh_5_9_io_out_c_0) ^ ((fiEnable && (1024 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_9_io_in_control_0_shift_b <=( _mesh_5_9_io_out_control_0_shift) ^ ((fiEnable && (1025 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_9_io_in_control_0_dataflow_b <=( _mesh_5_9_io_out_control_0_dataflow) ^ ((fiEnable && (1026 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_9_io_in_control_0_propagate_b <=( _mesh_5_9_io_out_control_0_propagate) ^ ((fiEnable && (1027 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_9_io_out_valid_0) begin
			b_151_0 <=( _mesh_6_9_io_out_b_0) ^ ((fiEnable && (1028 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_407_0 <=( _mesh_6_9_io_out_c_0) ^ ((fiEnable && (1029 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_9_io_in_control_0_shift_b <=( _mesh_6_9_io_out_control_0_shift) ^ ((fiEnable && (1030 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_9_io_in_control_0_dataflow_b <=( _mesh_6_9_io_out_control_0_dataflow) ^ ((fiEnable && (1031 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_9_io_in_control_0_propagate_b <=( _mesh_6_9_io_out_control_0_propagate) ^ ((fiEnable && (1032 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_9_io_out_valid_0) begin
			b_152_0 <=( _mesh_7_9_io_out_b_0) ^ ((fiEnable && (1033 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_408_0 <=( _mesh_7_9_io_out_c_0) ^ ((fiEnable && (1034 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_9_io_in_control_0_shift_b <=( _mesh_7_9_io_out_control_0_shift) ^ ((fiEnable && (1035 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_9_io_in_control_0_dataflow_b <=( _mesh_7_9_io_out_control_0_dataflow) ^ ((fiEnable && (1036 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_9_io_in_control_0_propagate_b <=( _mesh_7_9_io_out_control_0_propagate) ^ ((fiEnable && (1037 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_9_io_out_valid_0) begin
			b_153_0 <=( _mesh_8_9_io_out_b_0) ^ ((fiEnable && (1038 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_409_0 <=( _mesh_8_9_io_out_c_0) ^ ((fiEnable && (1039 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_9_io_in_control_0_shift_b <=( _mesh_8_9_io_out_control_0_shift) ^ ((fiEnable && (1040 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_9_io_in_control_0_dataflow_b <=( _mesh_8_9_io_out_control_0_dataflow) ^ ((fiEnable && (1041 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_9_io_in_control_0_propagate_b <=( _mesh_8_9_io_out_control_0_propagate) ^ ((fiEnable && (1042 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_9_io_out_valid_0) begin
			b_154_0 <=( _mesh_9_9_io_out_b_0) ^ ((fiEnable && (1043 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_410_0 <=( _mesh_9_9_io_out_c_0) ^ ((fiEnable && (1044 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_9_io_in_control_0_shift_b <=( _mesh_9_9_io_out_control_0_shift) ^ ((fiEnable && (1045 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_9_io_in_control_0_dataflow_b <=( _mesh_9_9_io_out_control_0_dataflow) ^ ((fiEnable && (1046 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_9_io_in_control_0_propagate_b <=( _mesh_9_9_io_out_control_0_propagate) ^ ((fiEnable && (1047 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_9_io_out_valid_0) begin
			b_155_0 <=( _mesh_10_9_io_out_b_0) ^ ((fiEnable && (1048 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_411_0 <=( _mesh_10_9_io_out_c_0) ^ ((fiEnable && (1049 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_9_io_in_control_0_shift_b <=( _mesh_10_9_io_out_control_0_shift) ^ ((fiEnable && (1050 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_9_io_in_control_0_dataflow_b <=( _mesh_10_9_io_out_control_0_dataflow) ^ ((fiEnable && (1051 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_9_io_in_control_0_propagate_b <=( _mesh_10_9_io_out_control_0_propagate) ^ ((fiEnable && (1052 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_9_io_out_valid_0) begin
			b_156_0 <=( _mesh_11_9_io_out_b_0) ^ ((fiEnable && (1053 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_412_0 <=( _mesh_11_9_io_out_c_0) ^ ((fiEnable && (1054 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_9_io_in_control_0_shift_b <=( _mesh_11_9_io_out_control_0_shift) ^ ((fiEnable && (1055 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_9_io_in_control_0_dataflow_b <=( _mesh_11_9_io_out_control_0_dataflow) ^ ((fiEnable && (1056 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_9_io_in_control_0_propagate_b <=( _mesh_11_9_io_out_control_0_propagate) ^ ((fiEnable && (1057 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_9_io_out_valid_0) begin
			b_157_0 <=( _mesh_12_9_io_out_b_0) ^ ((fiEnable && (1058 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_413_0 <=( _mesh_12_9_io_out_c_0) ^ ((fiEnable && (1059 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_9_io_in_control_0_shift_b <=( _mesh_12_9_io_out_control_0_shift) ^ ((fiEnable && (1060 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_9_io_in_control_0_dataflow_b <=( _mesh_12_9_io_out_control_0_dataflow) ^ ((fiEnable && (1061 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_9_io_in_control_0_propagate_b <=( _mesh_12_9_io_out_control_0_propagate) ^ ((fiEnable && (1062 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_9_io_out_valid_0) begin
			b_158_0 <=( _mesh_13_9_io_out_b_0) ^ ((fiEnable && (1063 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_414_0 <=( _mesh_13_9_io_out_c_0) ^ ((fiEnable && (1064 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_9_io_in_control_0_shift_b <=( _mesh_13_9_io_out_control_0_shift) ^ ((fiEnable && (1065 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_9_io_in_control_0_dataflow_b <=( _mesh_13_9_io_out_control_0_dataflow) ^ ((fiEnable && (1066 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_9_io_in_control_0_propagate_b <=( _mesh_13_9_io_out_control_0_propagate) ^ ((fiEnable && (1067 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_9_io_out_valid_0) begin
			b_159_0 <=( _mesh_14_9_io_out_b_0) ^ ((fiEnable && (1068 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_415_0 <=( _mesh_14_9_io_out_c_0) ^ ((fiEnable && (1069 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_9_io_in_control_0_shift_b <=( _mesh_14_9_io_out_control_0_shift) ^ ((fiEnable && (1070 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_9_io_in_control_0_dataflow_b <=( _mesh_14_9_io_out_control_0_dataflow) ^ ((fiEnable && (1071 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_9_io_in_control_0_propagate_b <=( _mesh_14_9_io_out_control_0_propagate) ^ ((fiEnable && (1072 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_10_0) begin
			b_160_0 <=( io_in_b_10_0) ^ ((fiEnable && (1073 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_416_0 <=( io_in_d_10_0) ^ ((fiEnable && (1074 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_10_io_in_control_0_shift_b <=( io_in_control_10_0_shift) ^ ((fiEnable && (1075 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_10_io_in_control_0_dataflow_b <=( io_in_control_10_0_dataflow) ^ ((fiEnable && (1076 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_10_io_in_control_0_propagate_b <=( io_in_control_10_0_propagate) ^ ((fiEnable && (1077 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_10_io_out_valid_0) begin
			b_161_0 <=( _mesh_0_10_io_out_b_0) ^ ((fiEnable && (1078 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_417_0 <=( _mesh_0_10_io_out_c_0) ^ ((fiEnable && (1079 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_10_io_in_control_0_shift_b <=( _mesh_0_10_io_out_control_0_shift) ^ ((fiEnable && (1080 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_10_io_in_control_0_dataflow_b <=( _mesh_0_10_io_out_control_0_dataflow) ^ ((fiEnable && (1081 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_10_io_in_control_0_propagate_b <=( _mesh_0_10_io_out_control_0_propagate) ^ ((fiEnable && (1082 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_10_io_out_valid_0) begin
			b_162_0 <=( _mesh_1_10_io_out_b_0) ^ ((fiEnable && (1083 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_418_0 <=( _mesh_1_10_io_out_c_0) ^ ((fiEnable && (1084 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_10_io_in_control_0_shift_b <=( _mesh_1_10_io_out_control_0_shift) ^ ((fiEnable && (1085 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_10_io_in_control_0_dataflow_b <=( _mesh_1_10_io_out_control_0_dataflow) ^ ((fiEnable && (1086 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_10_io_in_control_0_propagate_b <=( _mesh_1_10_io_out_control_0_propagate) ^ ((fiEnable && (1087 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_10_io_out_valid_0) begin
			b_163_0 <=( _mesh_2_10_io_out_b_0) ^ ((fiEnable && (1088 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_419_0 <=( _mesh_2_10_io_out_c_0) ^ ((fiEnable && (1089 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_10_io_in_control_0_shift_b <=( _mesh_2_10_io_out_control_0_shift) ^ ((fiEnable && (1090 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_10_io_in_control_0_dataflow_b <=( _mesh_2_10_io_out_control_0_dataflow) ^ ((fiEnable && (1091 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_10_io_in_control_0_propagate_b <=( _mesh_2_10_io_out_control_0_propagate) ^ ((fiEnable && (1092 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_10_io_out_valid_0) begin
			b_164_0 <=( _mesh_3_10_io_out_b_0) ^ ((fiEnable && (1093 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_420_0 <=( _mesh_3_10_io_out_c_0) ^ ((fiEnable && (1094 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_10_io_in_control_0_shift_b <=( _mesh_3_10_io_out_control_0_shift) ^ ((fiEnable && (1095 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_10_io_in_control_0_dataflow_b <=( _mesh_3_10_io_out_control_0_dataflow) ^ ((fiEnable && (1096 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_10_io_in_control_0_propagate_b <=( _mesh_3_10_io_out_control_0_propagate) ^ ((fiEnable && (1097 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_10_io_out_valid_0) begin
			b_165_0 <=( _mesh_4_10_io_out_b_0) ^ ((fiEnable && (1098 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_421_0 <=( _mesh_4_10_io_out_c_0) ^ ((fiEnable && (1099 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_10_io_in_control_0_shift_b <=( _mesh_4_10_io_out_control_0_shift) ^ ((fiEnable && (1100 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_10_io_in_control_0_dataflow_b <=( _mesh_4_10_io_out_control_0_dataflow) ^ ((fiEnable && (1101 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_10_io_in_control_0_propagate_b <=( _mesh_4_10_io_out_control_0_propagate) ^ ((fiEnable && (1102 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_10_io_out_valid_0) begin
			b_166_0 <=( _mesh_5_10_io_out_b_0) ^ ((fiEnable && (1103 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_422_0 <=( _mesh_5_10_io_out_c_0) ^ ((fiEnable && (1104 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_10_io_in_control_0_shift_b <=( _mesh_5_10_io_out_control_0_shift) ^ ((fiEnable && (1105 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_10_io_in_control_0_dataflow_b <=( _mesh_5_10_io_out_control_0_dataflow) ^ ((fiEnable && (1106 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_10_io_in_control_0_propagate_b <=( _mesh_5_10_io_out_control_0_propagate) ^ ((fiEnable && (1107 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_10_io_out_valid_0) begin
			b_167_0 <=( _mesh_6_10_io_out_b_0) ^ ((fiEnable && (1108 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_423_0 <=( _mesh_6_10_io_out_c_0) ^ ((fiEnable && (1109 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_10_io_in_control_0_shift_b <=( _mesh_6_10_io_out_control_0_shift) ^ ((fiEnable && (1110 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_10_io_in_control_0_dataflow_b <=( _mesh_6_10_io_out_control_0_dataflow) ^ ((fiEnable && (1111 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_10_io_in_control_0_propagate_b <=( _mesh_6_10_io_out_control_0_propagate) ^ ((fiEnable && (1112 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_10_io_out_valid_0) begin
			b_168_0 <=( _mesh_7_10_io_out_b_0) ^ ((fiEnable && (1113 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_424_0 <=( _mesh_7_10_io_out_c_0) ^ ((fiEnable && (1114 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_10_io_in_control_0_shift_b <=( _mesh_7_10_io_out_control_0_shift) ^ ((fiEnable && (1115 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_10_io_in_control_0_dataflow_b <=( _mesh_7_10_io_out_control_0_dataflow) ^ ((fiEnable && (1116 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_10_io_in_control_0_propagate_b <=( _mesh_7_10_io_out_control_0_propagate) ^ ((fiEnable && (1117 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_10_io_out_valid_0) begin
			b_169_0 <=( _mesh_8_10_io_out_b_0) ^ ((fiEnable && (1118 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_425_0 <=( _mesh_8_10_io_out_c_0) ^ ((fiEnable && (1119 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_10_io_in_control_0_shift_b <=( _mesh_8_10_io_out_control_0_shift) ^ ((fiEnable && (1120 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_10_io_in_control_0_dataflow_b <=( _mesh_8_10_io_out_control_0_dataflow) ^ ((fiEnable && (1121 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_10_io_in_control_0_propagate_b <=( _mesh_8_10_io_out_control_0_propagate) ^ ((fiEnable && (1122 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_10_io_out_valid_0) begin
			b_170_0 <=( _mesh_9_10_io_out_b_0) ^ ((fiEnable && (1123 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_426_0 <=( _mesh_9_10_io_out_c_0) ^ ((fiEnable && (1124 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_10_io_in_control_0_shift_b <=( _mesh_9_10_io_out_control_0_shift) ^ ((fiEnable && (1125 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_10_io_in_control_0_dataflow_b <=( _mesh_9_10_io_out_control_0_dataflow) ^ ((fiEnable && (1126 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_10_io_in_control_0_propagate_b <=( _mesh_9_10_io_out_control_0_propagate) ^ ((fiEnable && (1127 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_10_io_out_valid_0) begin
			b_171_0 <=( _mesh_10_10_io_out_b_0) ^ ((fiEnable && (1128 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_427_0 <=( _mesh_10_10_io_out_c_0) ^ ((fiEnable && (1129 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_10_io_in_control_0_shift_b <=( _mesh_10_10_io_out_control_0_shift) ^ ((fiEnable && (1130 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_10_io_in_control_0_dataflow_b <=( _mesh_10_10_io_out_control_0_dataflow) ^ ((fiEnable && (1131 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_10_io_in_control_0_propagate_b <=( _mesh_10_10_io_out_control_0_propagate) ^ ((fiEnable && (1132 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_10_io_out_valid_0) begin
			b_172_0 <=( _mesh_11_10_io_out_b_0) ^ ((fiEnable && (1133 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_428_0 <=( _mesh_11_10_io_out_c_0) ^ ((fiEnable && (1134 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_10_io_in_control_0_shift_b <=( _mesh_11_10_io_out_control_0_shift) ^ ((fiEnable && (1135 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_10_io_in_control_0_dataflow_b <=( _mesh_11_10_io_out_control_0_dataflow) ^ ((fiEnable && (1136 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_10_io_in_control_0_propagate_b <=( _mesh_11_10_io_out_control_0_propagate) ^ ((fiEnable && (1137 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_10_io_out_valid_0) begin
			b_173_0 <=( _mesh_12_10_io_out_b_0) ^ ((fiEnable && (1138 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_429_0 <=( _mesh_12_10_io_out_c_0) ^ ((fiEnable && (1139 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_10_io_in_control_0_shift_b <=( _mesh_12_10_io_out_control_0_shift) ^ ((fiEnable && (1140 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_10_io_in_control_0_dataflow_b <=( _mesh_12_10_io_out_control_0_dataflow) ^ ((fiEnable && (1141 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_10_io_in_control_0_propagate_b <=( _mesh_12_10_io_out_control_0_propagate) ^ ((fiEnable && (1142 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_10_io_out_valid_0) begin
			b_174_0 <=( _mesh_13_10_io_out_b_0) ^ ((fiEnable && (1143 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_430_0 <=( _mesh_13_10_io_out_c_0) ^ ((fiEnable && (1144 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_10_io_in_control_0_shift_b <=( _mesh_13_10_io_out_control_0_shift) ^ ((fiEnable && (1145 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_10_io_in_control_0_dataflow_b <=( _mesh_13_10_io_out_control_0_dataflow) ^ ((fiEnable && (1146 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_10_io_in_control_0_propagate_b <=( _mesh_13_10_io_out_control_0_propagate) ^ ((fiEnable && (1147 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_10_io_out_valid_0) begin
			b_175_0 <=( _mesh_14_10_io_out_b_0) ^ ((fiEnable && (1148 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_431_0 <=( _mesh_14_10_io_out_c_0) ^ ((fiEnable && (1149 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_10_io_in_control_0_shift_b <=( _mesh_14_10_io_out_control_0_shift) ^ ((fiEnable && (1150 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_10_io_in_control_0_dataflow_b <=( _mesh_14_10_io_out_control_0_dataflow) ^ ((fiEnable && (1151 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_10_io_in_control_0_propagate_b <=( _mesh_14_10_io_out_control_0_propagate) ^ ((fiEnable && (1152 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_11_0) begin
			b_176_0 <=( io_in_b_11_0) ^ ((fiEnable && (1153 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_432_0 <=( io_in_d_11_0) ^ ((fiEnable && (1154 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_11_io_in_control_0_shift_b <=( io_in_control_11_0_shift) ^ ((fiEnable && (1155 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_11_io_in_control_0_dataflow_b <=( io_in_control_11_0_dataflow) ^ ((fiEnable && (1156 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_11_io_in_control_0_propagate_b <=( io_in_control_11_0_propagate) ^ ((fiEnable && (1157 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_11_io_out_valid_0) begin
			b_177_0 <=( _mesh_0_11_io_out_b_0) ^ ((fiEnable && (1158 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_433_0 <=( _mesh_0_11_io_out_c_0) ^ ((fiEnable && (1159 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_11_io_in_control_0_shift_b <=( _mesh_0_11_io_out_control_0_shift) ^ ((fiEnable && (1160 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_11_io_in_control_0_dataflow_b <=( _mesh_0_11_io_out_control_0_dataflow) ^ ((fiEnable && (1161 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_11_io_in_control_0_propagate_b <=( _mesh_0_11_io_out_control_0_propagate) ^ ((fiEnable && (1162 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_11_io_out_valid_0) begin
			b_178_0 <=( _mesh_1_11_io_out_b_0) ^ ((fiEnable && (1163 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_434_0 <=( _mesh_1_11_io_out_c_0) ^ ((fiEnable && (1164 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_11_io_in_control_0_shift_b <=( _mesh_1_11_io_out_control_0_shift) ^ ((fiEnable && (1165 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_11_io_in_control_0_dataflow_b <=( _mesh_1_11_io_out_control_0_dataflow) ^ ((fiEnable && (1166 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_11_io_in_control_0_propagate_b <=( _mesh_1_11_io_out_control_0_propagate) ^ ((fiEnable && (1167 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_11_io_out_valid_0) begin
			b_179_0 <=( _mesh_2_11_io_out_b_0) ^ ((fiEnable && (1168 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_435_0 <=( _mesh_2_11_io_out_c_0) ^ ((fiEnable && (1169 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_11_io_in_control_0_shift_b <=( _mesh_2_11_io_out_control_0_shift) ^ ((fiEnable && (1170 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_11_io_in_control_0_dataflow_b <=( _mesh_2_11_io_out_control_0_dataflow) ^ ((fiEnable && (1171 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_11_io_in_control_0_propagate_b <=( _mesh_2_11_io_out_control_0_propagate) ^ ((fiEnable && (1172 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_11_io_out_valid_0) begin
			b_180_0 <=( _mesh_3_11_io_out_b_0) ^ ((fiEnable && (1173 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_436_0 <=( _mesh_3_11_io_out_c_0) ^ ((fiEnable && (1174 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_11_io_in_control_0_shift_b <=( _mesh_3_11_io_out_control_0_shift) ^ ((fiEnable && (1175 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_11_io_in_control_0_dataflow_b <=( _mesh_3_11_io_out_control_0_dataflow) ^ ((fiEnable && (1176 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_11_io_in_control_0_propagate_b <=( _mesh_3_11_io_out_control_0_propagate) ^ ((fiEnable && (1177 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_11_io_out_valid_0) begin
			b_181_0 <=( _mesh_4_11_io_out_b_0) ^ ((fiEnable && (1178 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_437_0 <=( _mesh_4_11_io_out_c_0) ^ ((fiEnable && (1179 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_11_io_in_control_0_shift_b <=( _mesh_4_11_io_out_control_0_shift) ^ ((fiEnable && (1180 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_11_io_in_control_0_dataflow_b <=( _mesh_4_11_io_out_control_0_dataflow) ^ ((fiEnable && (1181 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_11_io_in_control_0_propagate_b <=( _mesh_4_11_io_out_control_0_propagate) ^ ((fiEnable && (1182 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_11_io_out_valid_0) begin
			b_182_0 <=( _mesh_5_11_io_out_b_0) ^ ((fiEnable && (1183 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_438_0 <=( _mesh_5_11_io_out_c_0) ^ ((fiEnable && (1184 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_11_io_in_control_0_shift_b <=( _mesh_5_11_io_out_control_0_shift) ^ ((fiEnable && (1185 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_11_io_in_control_0_dataflow_b <=( _mesh_5_11_io_out_control_0_dataflow) ^ ((fiEnable && (1186 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_11_io_in_control_0_propagate_b <=( _mesh_5_11_io_out_control_0_propagate) ^ ((fiEnable && (1187 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_11_io_out_valid_0) begin
			b_183_0 <=( _mesh_6_11_io_out_b_0) ^ ((fiEnable && (1188 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_439_0 <=( _mesh_6_11_io_out_c_0) ^ ((fiEnable && (1189 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_11_io_in_control_0_shift_b <=( _mesh_6_11_io_out_control_0_shift) ^ ((fiEnable && (1190 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_11_io_in_control_0_dataflow_b <=( _mesh_6_11_io_out_control_0_dataflow) ^ ((fiEnable && (1191 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_11_io_in_control_0_propagate_b <=( _mesh_6_11_io_out_control_0_propagate) ^ ((fiEnable && (1192 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_11_io_out_valid_0) begin
			b_184_0 <=( _mesh_7_11_io_out_b_0) ^ ((fiEnable && (1193 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_440_0 <=( _mesh_7_11_io_out_c_0) ^ ((fiEnable && (1194 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_11_io_in_control_0_shift_b <=( _mesh_7_11_io_out_control_0_shift) ^ ((fiEnable && (1195 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_11_io_in_control_0_dataflow_b <=( _mesh_7_11_io_out_control_0_dataflow) ^ ((fiEnable && (1196 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_11_io_in_control_0_propagate_b <=( _mesh_7_11_io_out_control_0_propagate) ^ ((fiEnable && (1197 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_11_io_out_valid_0) begin
			b_185_0 <=( _mesh_8_11_io_out_b_0) ^ ((fiEnable && (1198 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_441_0 <=( _mesh_8_11_io_out_c_0) ^ ((fiEnable && (1199 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_11_io_in_control_0_shift_b <=( _mesh_8_11_io_out_control_0_shift) ^ ((fiEnable && (1200 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_11_io_in_control_0_dataflow_b <=( _mesh_8_11_io_out_control_0_dataflow) ^ ((fiEnable && (1201 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_11_io_in_control_0_propagate_b <=( _mesh_8_11_io_out_control_0_propagate) ^ ((fiEnable && (1202 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_11_io_out_valid_0) begin
			b_186_0 <=( _mesh_9_11_io_out_b_0) ^ ((fiEnable && (1203 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_442_0 <=( _mesh_9_11_io_out_c_0) ^ ((fiEnable && (1204 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_11_io_in_control_0_shift_b <=( _mesh_9_11_io_out_control_0_shift) ^ ((fiEnable && (1205 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_11_io_in_control_0_dataflow_b <=( _mesh_9_11_io_out_control_0_dataflow) ^ ((fiEnable && (1206 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_11_io_in_control_0_propagate_b <=( _mesh_9_11_io_out_control_0_propagate) ^ ((fiEnable && (1207 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_11_io_out_valid_0) begin
			b_187_0 <=( _mesh_10_11_io_out_b_0) ^ ((fiEnable && (1208 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_443_0 <=( _mesh_10_11_io_out_c_0) ^ ((fiEnable && (1209 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_11_io_in_control_0_shift_b <=( _mesh_10_11_io_out_control_0_shift) ^ ((fiEnable && (1210 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_11_io_in_control_0_dataflow_b <=( _mesh_10_11_io_out_control_0_dataflow) ^ ((fiEnable && (1211 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_11_io_in_control_0_propagate_b <=( _mesh_10_11_io_out_control_0_propagate) ^ ((fiEnable && (1212 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_11_io_out_valid_0) begin
			b_188_0 <=( _mesh_11_11_io_out_b_0) ^ ((fiEnable && (1213 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_444_0 <=( _mesh_11_11_io_out_c_0) ^ ((fiEnable && (1214 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_11_io_in_control_0_shift_b <=( _mesh_11_11_io_out_control_0_shift) ^ ((fiEnable && (1215 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_11_io_in_control_0_dataflow_b <=( _mesh_11_11_io_out_control_0_dataflow) ^ ((fiEnable && (1216 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_11_io_in_control_0_propagate_b <=( _mesh_11_11_io_out_control_0_propagate) ^ ((fiEnable && (1217 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_11_io_out_valid_0) begin
			b_189_0 <=( _mesh_12_11_io_out_b_0) ^ ((fiEnable && (1218 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_445_0 <=( _mesh_12_11_io_out_c_0) ^ ((fiEnable && (1219 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_11_io_in_control_0_shift_b <=( _mesh_12_11_io_out_control_0_shift) ^ ((fiEnable && (1220 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_11_io_in_control_0_dataflow_b <=( _mesh_12_11_io_out_control_0_dataflow) ^ ((fiEnable && (1221 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_11_io_in_control_0_propagate_b <=( _mesh_12_11_io_out_control_0_propagate) ^ ((fiEnable && (1222 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_11_io_out_valid_0) begin
			b_190_0 <=( _mesh_13_11_io_out_b_0) ^ ((fiEnable && (1223 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_446_0 <=( _mesh_13_11_io_out_c_0) ^ ((fiEnable && (1224 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_11_io_in_control_0_shift_b <=( _mesh_13_11_io_out_control_0_shift) ^ ((fiEnable && (1225 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_11_io_in_control_0_dataflow_b <=( _mesh_13_11_io_out_control_0_dataflow) ^ ((fiEnable && (1226 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_11_io_in_control_0_propagate_b <=( _mesh_13_11_io_out_control_0_propagate) ^ ((fiEnable && (1227 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_11_io_out_valid_0) begin
			b_191_0 <=( _mesh_14_11_io_out_b_0) ^ ((fiEnable && (1228 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_447_0 <=( _mesh_14_11_io_out_c_0) ^ ((fiEnable && (1229 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_11_io_in_control_0_shift_b <=( _mesh_14_11_io_out_control_0_shift) ^ ((fiEnable && (1230 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_11_io_in_control_0_dataflow_b <=( _mesh_14_11_io_out_control_0_dataflow) ^ ((fiEnable && (1231 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_11_io_in_control_0_propagate_b <=( _mesh_14_11_io_out_control_0_propagate) ^ ((fiEnable && (1232 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_12_0) begin
			b_192_0 <=( io_in_b_12_0) ^ ((fiEnable && (1233 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_448_0 <=( io_in_d_12_0) ^ ((fiEnable && (1234 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_12_io_in_control_0_shift_b <=( io_in_control_12_0_shift) ^ ((fiEnable && (1235 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_12_io_in_control_0_dataflow_b <=( io_in_control_12_0_dataflow) ^ ((fiEnable && (1236 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_12_io_in_control_0_propagate_b <=( io_in_control_12_0_propagate) ^ ((fiEnable && (1237 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_12_io_out_valid_0) begin
			b_193_0 <=( _mesh_0_12_io_out_b_0) ^ ((fiEnable && (1238 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_449_0 <=( _mesh_0_12_io_out_c_0) ^ ((fiEnable && (1239 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_12_io_in_control_0_shift_b <=( _mesh_0_12_io_out_control_0_shift) ^ ((fiEnable && (1240 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_12_io_in_control_0_dataflow_b <=( _mesh_0_12_io_out_control_0_dataflow) ^ ((fiEnable && (1241 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_12_io_in_control_0_propagate_b <=( _mesh_0_12_io_out_control_0_propagate) ^ ((fiEnable && (1242 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_12_io_out_valid_0) begin
			b_194_0 <=( _mesh_1_12_io_out_b_0) ^ ((fiEnable && (1243 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_450_0 <=( _mesh_1_12_io_out_c_0) ^ ((fiEnable && (1244 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_12_io_in_control_0_shift_b <=( _mesh_1_12_io_out_control_0_shift) ^ ((fiEnable && (1245 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_12_io_in_control_0_dataflow_b <=( _mesh_1_12_io_out_control_0_dataflow) ^ ((fiEnable && (1246 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_12_io_in_control_0_propagate_b <=( _mesh_1_12_io_out_control_0_propagate) ^ ((fiEnable && (1247 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_12_io_out_valid_0) begin
			b_195_0 <=( _mesh_2_12_io_out_b_0) ^ ((fiEnable && (1248 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_451_0 <=( _mesh_2_12_io_out_c_0) ^ ((fiEnable && (1249 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_12_io_in_control_0_shift_b <=( _mesh_2_12_io_out_control_0_shift) ^ ((fiEnable && (1250 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_12_io_in_control_0_dataflow_b <=( _mesh_2_12_io_out_control_0_dataflow) ^ ((fiEnable && (1251 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_12_io_in_control_0_propagate_b <=( _mesh_2_12_io_out_control_0_propagate) ^ ((fiEnable && (1252 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_12_io_out_valid_0) begin
			b_196_0 <=( _mesh_3_12_io_out_b_0) ^ ((fiEnable && (1253 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_452_0 <=( _mesh_3_12_io_out_c_0) ^ ((fiEnable && (1254 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_12_io_in_control_0_shift_b <=( _mesh_3_12_io_out_control_0_shift) ^ ((fiEnable && (1255 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_12_io_in_control_0_dataflow_b <=( _mesh_3_12_io_out_control_0_dataflow) ^ ((fiEnable && (1256 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_12_io_in_control_0_propagate_b <=( _mesh_3_12_io_out_control_0_propagate) ^ ((fiEnable && (1257 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_12_io_out_valid_0) begin
			b_197_0 <=( _mesh_4_12_io_out_b_0) ^ ((fiEnable && (1258 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_453_0 <=( _mesh_4_12_io_out_c_0) ^ ((fiEnable && (1259 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_12_io_in_control_0_shift_b <=( _mesh_4_12_io_out_control_0_shift) ^ ((fiEnable && (1260 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_12_io_in_control_0_dataflow_b <=( _mesh_4_12_io_out_control_0_dataflow) ^ ((fiEnable && (1261 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_12_io_in_control_0_propagate_b <=( _mesh_4_12_io_out_control_0_propagate) ^ ((fiEnable && (1262 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_12_io_out_valid_0) begin
			b_198_0 <=( _mesh_5_12_io_out_b_0) ^ ((fiEnable && (1263 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_454_0 <=( _mesh_5_12_io_out_c_0) ^ ((fiEnable && (1264 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_12_io_in_control_0_shift_b <=( _mesh_5_12_io_out_control_0_shift) ^ ((fiEnable && (1265 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_12_io_in_control_0_dataflow_b <=( _mesh_5_12_io_out_control_0_dataflow) ^ ((fiEnable && (1266 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_12_io_in_control_0_propagate_b <=( _mesh_5_12_io_out_control_0_propagate) ^ ((fiEnable && (1267 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_12_io_out_valid_0) begin
			b_199_0 <=( _mesh_6_12_io_out_b_0) ^ ((fiEnable && (1268 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_455_0 <=( _mesh_6_12_io_out_c_0) ^ ((fiEnable && (1269 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_12_io_in_control_0_shift_b <=( _mesh_6_12_io_out_control_0_shift) ^ ((fiEnable && (1270 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_12_io_in_control_0_dataflow_b <=( _mesh_6_12_io_out_control_0_dataflow) ^ ((fiEnable && (1271 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_12_io_in_control_0_propagate_b <=( _mesh_6_12_io_out_control_0_propagate) ^ ((fiEnable && (1272 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_12_io_out_valid_0) begin
			b_200_0 <=( _mesh_7_12_io_out_b_0) ^ ((fiEnable && (1273 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_456_0 <=( _mesh_7_12_io_out_c_0) ^ ((fiEnable && (1274 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_12_io_in_control_0_shift_b <=( _mesh_7_12_io_out_control_0_shift) ^ ((fiEnable && (1275 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_12_io_in_control_0_dataflow_b <=( _mesh_7_12_io_out_control_0_dataflow) ^ ((fiEnable && (1276 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_12_io_in_control_0_propagate_b <=( _mesh_7_12_io_out_control_0_propagate) ^ ((fiEnable && (1277 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_12_io_out_valid_0) begin
			b_201_0 <=( _mesh_8_12_io_out_b_0) ^ ((fiEnable && (1278 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_457_0 <=( _mesh_8_12_io_out_c_0) ^ ((fiEnable && (1279 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_12_io_in_control_0_shift_b <=( _mesh_8_12_io_out_control_0_shift) ^ ((fiEnable && (1280 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_12_io_in_control_0_dataflow_b <=( _mesh_8_12_io_out_control_0_dataflow) ^ ((fiEnable && (1281 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_12_io_in_control_0_propagate_b <=( _mesh_8_12_io_out_control_0_propagate) ^ ((fiEnable && (1282 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_12_io_out_valid_0) begin
			b_202_0 <=( _mesh_9_12_io_out_b_0) ^ ((fiEnable && (1283 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_458_0 <=( _mesh_9_12_io_out_c_0) ^ ((fiEnable && (1284 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_12_io_in_control_0_shift_b <=( _mesh_9_12_io_out_control_0_shift) ^ ((fiEnable && (1285 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_12_io_in_control_0_dataflow_b <=( _mesh_9_12_io_out_control_0_dataflow) ^ ((fiEnable && (1286 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_12_io_in_control_0_propagate_b <=( _mesh_9_12_io_out_control_0_propagate) ^ ((fiEnable && (1287 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_12_io_out_valid_0) begin
			b_203_0 <=( _mesh_10_12_io_out_b_0) ^ ((fiEnable && (1288 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_459_0 <=( _mesh_10_12_io_out_c_0) ^ ((fiEnable && (1289 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_12_io_in_control_0_shift_b <=( _mesh_10_12_io_out_control_0_shift) ^ ((fiEnable && (1290 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_12_io_in_control_0_dataflow_b <=( _mesh_10_12_io_out_control_0_dataflow) ^ ((fiEnable && (1291 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_12_io_in_control_0_propagate_b <=( _mesh_10_12_io_out_control_0_propagate) ^ ((fiEnable && (1292 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_12_io_out_valid_0) begin
			b_204_0 <=( _mesh_11_12_io_out_b_0) ^ ((fiEnable && (1293 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_460_0 <=( _mesh_11_12_io_out_c_0) ^ ((fiEnable && (1294 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_12_io_in_control_0_shift_b <=( _mesh_11_12_io_out_control_0_shift) ^ ((fiEnable && (1295 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_12_io_in_control_0_dataflow_b <=( _mesh_11_12_io_out_control_0_dataflow) ^ ((fiEnable && (1296 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_12_io_in_control_0_propagate_b <=( _mesh_11_12_io_out_control_0_propagate) ^ ((fiEnable && (1297 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_12_io_out_valid_0) begin
			b_205_0 <=( _mesh_12_12_io_out_b_0) ^ ((fiEnable && (1298 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_461_0 <=( _mesh_12_12_io_out_c_0) ^ ((fiEnable && (1299 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_12_io_in_control_0_shift_b <=( _mesh_12_12_io_out_control_0_shift) ^ ((fiEnable && (1300 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_12_io_in_control_0_dataflow_b <=( _mesh_12_12_io_out_control_0_dataflow) ^ ((fiEnable && (1301 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_12_io_in_control_0_propagate_b <=( _mesh_12_12_io_out_control_0_propagate) ^ ((fiEnable && (1302 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_12_io_out_valid_0) begin
			b_206_0 <=( _mesh_13_12_io_out_b_0) ^ ((fiEnable && (1303 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_462_0 <=( _mesh_13_12_io_out_c_0) ^ ((fiEnable && (1304 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_12_io_in_control_0_shift_b <=( _mesh_13_12_io_out_control_0_shift) ^ ((fiEnable && (1305 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_12_io_in_control_0_dataflow_b <=( _mesh_13_12_io_out_control_0_dataflow) ^ ((fiEnable && (1306 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_12_io_in_control_0_propagate_b <=( _mesh_13_12_io_out_control_0_propagate) ^ ((fiEnable && (1307 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_12_io_out_valid_0) begin
			b_207_0 <=( _mesh_14_12_io_out_b_0) ^ ((fiEnable && (1308 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_463_0 <=( _mesh_14_12_io_out_c_0) ^ ((fiEnable && (1309 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_12_io_in_control_0_shift_b <=( _mesh_14_12_io_out_control_0_shift) ^ ((fiEnable && (1310 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_12_io_in_control_0_dataflow_b <=( _mesh_14_12_io_out_control_0_dataflow) ^ ((fiEnable && (1311 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_12_io_in_control_0_propagate_b <=( _mesh_14_12_io_out_control_0_propagate) ^ ((fiEnable && (1312 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_13_0) begin
			b_208_0 <=( io_in_b_13_0) ^ ((fiEnable && (1313 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_464_0 <=( io_in_d_13_0) ^ ((fiEnable && (1314 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_13_io_in_control_0_shift_b <=( io_in_control_13_0_shift) ^ ((fiEnable && (1315 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_13_io_in_control_0_dataflow_b <=( io_in_control_13_0_dataflow) ^ ((fiEnable && (1316 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_13_io_in_control_0_propagate_b <=( io_in_control_13_0_propagate) ^ ((fiEnable && (1317 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_13_io_out_valid_0) begin
			b_209_0 <=( _mesh_0_13_io_out_b_0) ^ ((fiEnable && (1318 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_465_0 <=( _mesh_0_13_io_out_c_0) ^ ((fiEnable && (1319 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_13_io_in_control_0_shift_b <=( _mesh_0_13_io_out_control_0_shift) ^ ((fiEnable && (1320 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_13_io_in_control_0_dataflow_b <=( _mesh_0_13_io_out_control_0_dataflow) ^ ((fiEnable && (1321 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_13_io_in_control_0_propagate_b <=( _mesh_0_13_io_out_control_0_propagate) ^ ((fiEnable && (1322 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_13_io_out_valid_0) begin
			b_210_0 <=( _mesh_1_13_io_out_b_0) ^ ((fiEnable && (1323 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_466_0 <=( _mesh_1_13_io_out_c_0) ^ ((fiEnable && (1324 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_13_io_in_control_0_shift_b <=( _mesh_1_13_io_out_control_0_shift) ^ ((fiEnable && (1325 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_13_io_in_control_0_dataflow_b <=( _mesh_1_13_io_out_control_0_dataflow) ^ ((fiEnable && (1326 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_13_io_in_control_0_propagate_b <=( _mesh_1_13_io_out_control_0_propagate) ^ ((fiEnable && (1327 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_13_io_out_valid_0) begin
			b_211_0 <=( _mesh_2_13_io_out_b_0) ^ ((fiEnable && (1328 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_467_0 <=( _mesh_2_13_io_out_c_0) ^ ((fiEnable && (1329 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_13_io_in_control_0_shift_b <=( _mesh_2_13_io_out_control_0_shift) ^ ((fiEnable && (1330 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_13_io_in_control_0_dataflow_b <=( _mesh_2_13_io_out_control_0_dataflow) ^ ((fiEnable && (1331 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_13_io_in_control_0_propagate_b <=( _mesh_2_13_io_out_control_0_propagate) ^ ((fiEnable && (1332 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_13_io_out_valid_0) begin
			b_212_0 <=( _mesh_3_13_io_out_b_0) ^ ((fiEnable && (1333 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_468_0 <=( _mesh_3_13_io_out_c_0) ^ ((fiEnable && (1334 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_13_io_in_control_0_shift_b <=( _mesh_3_13_io_out_control_0_shift) ^ ((fiEnable && (1335 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_13_io_in_control_0_dataflow_b <=( _mesh_3_13_io_out_control_0_dataflow) ^ ((fiEnable && (1336 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_13_io_in_control_0_propagate_b <=( _mesh_3_13_io_out_control_0_propagate) ^ ((fiEnable && (1337 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_13_io_out_valid_0) begin
			b_213_0 <=( _mesh_4_13_io_out_b_0) ^ ((fiEnable && (1338 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_469_0 <=( _mesh_4_13_io_out_c_0) ^ ((fiEnable && (1339 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_13_io_in_control_0_shift_b <=( _mesh_4_13_io_out_control_0_shift) ^ ((fiEnable && (1340 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_13_io_in_control_0_dataflow_b <=( _mesh_4_13_io_out_control_0_dataflow) ^ ((fiEnable && (1341 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_13_io_in_control_0_propagate_b <=( _mesh_4_13_io_out_control_0_propagate) ^ ((fiEnable && (1342 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_13_io_out_valid_0) begin
			b_214_0 <=( _mesh_5_13_io_out_b_0) ^ ((fiEnable && (1343 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_470_0 <=( _mesh_5_13_io_out_c_0) ^ ((fiEnable && (1344 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_13_io_in_control_0_shift_b <=( _mesh_5_13_io_out_control_0_shift) ^ ((fiEnable && (1345 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_13_io_in_control_0_dataflow_b <=( _mesh_5_13_io_out_control_0_dataflow) ^ ((fiEnable && (1346 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_13_io_in_control_0_propagate_b <=( _mesh_5_13_io_out_control_0_propagate) ^ ((fiEnable && (1347 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_13_io_out_valid_0) begin
			b_215_0 <=( _mesh_6_13_io_out_b_0) ^ ((fiEnable && (1348 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_471_0 <=( _mesh_6_13_io_out_c_0) ^ ((fiEnable && (1349 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_13_io_in_control_0_shift_b <=( _mesh_6_13_io_out_control_0_shift) ^ ((fiEnable && (1350 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_13_io_in_control_0_dataflow_b <=( _mesh_6_13_io_out_control_0_dataflow) ^ ((fiEnable && (1351 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_13_io_in_control_0_propagate_b <=( _mesh_6_13_io_out_control_0_propagate) ^ ((fiEnable && (1352 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_13_io_out_valid_0) begin
			b_216_0 <=( _mesh_7_13_io_out_b_0) ^ ((fiEnable && (1353 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_472_0 <=( _mesh_7_13_io_out_c_0) ^ ((fiEnable && (1354 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_13_io_in_control_0_shift_b <=( _mesh_7_13_io_out_control_0_shift) ^ ((fiEnable && (1355 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_13_io_in_control_0_dataflow_b <=( _mesh_7_13_io_out_control_0_dataflow) ^ ((fiEnable && (1356 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_13_io_in_control_0_propagate_b <=( _mesh_7_13_io_out_control_0_propagate) ^ ((fiEnable && (1357 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_13_io_out_valid_0) begin
			b_217_0 <=( _mesh_8_13_io_out_b_0) ^ ((fiEnable && (1358 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_473_0 <=( _mesh_8_13_io_out_c_0) ^ ((fiEnable && (1359 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_13_io_in_control_0_shift_b <=( _mesh_8_13_io_out_control_0_shift) ^ ((fiEnable && (1360 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_13_io_in_control_0_dataflow_b <=( _mesh_8_13_io_out_control_0_dataflow) ^ ((fiEnable && (1361 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_13_io_in_control_0_propagate_b <=( _mesh_8_13_io_out_control_0_propagate) ^ ((fiEnable && (1362 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_13_io_out_valid_0) begin
			b_218_0 <=( _mesh_9_13_io_out_b_0) ^ ((fiEnable && (1363 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_474_0 <=( _mesh_9_13_io_out_c_0) ^ ((fiEnable && (1364 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_13_io_in_control_0_shift_b <=( _mesh_9_13_io_out_control_0_shift) ^ ((fiEnable && (1365 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_13_io_in_control_0_dataflow_b <=( _mesh_9_13_io_out_control_0_dataflow) ^ ((fiEnable && (1366 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_13_io_in_control_0_propagate_b <=( _mesh_9_13_io_out_control_0_propagate) ^ ((fiEnable && (1367 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_13_io_out_valid_0) begin
			b_219_0 <=( _mesh_10_13_io_out_b_0) ^ ((fiEnable && (1368 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_475_0 <=( _mesh_10_13_io_out_c_0) ^ ((fiEnable && (1369 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_13_io_in_control_0_shift_b <=( _mesh_10_13_io_out_control_0_shift) ^ ((fiEnable && (1370 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_13_io_in_control_0_dataflow_b <=( _mesh_10_13_io_out_control_0_dataflow) ^ ((fiEnable && (1371 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_13_io_in_control_0_propagate_b <=( _mesh_10_13_io_out_control_0_propagate) ^ ((fiEnable && (1372 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_13_io_out_valid_0) begin
			b_220_0 <=( _mesh_11_13_io_out_b_0) ^ ((fiEnable && (1373 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_476_0 <=( _mesh_11_13_io_out_c_0) ^ ((fiEnable && (1374 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_13_io_in_control_0_shift_b <=( _mesh_11_13_io_out_control_0_shift) ^ ((fiEnable && (1375 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_13_io_in_control_0_dataflow_b <=( _mesh_11_13_io_out_control_0_dataflow) ^ ((fiEnable && (1376 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_13_io_in_control_0_propagate_b <=( _mesh_11_13_io_out_control_0_propagate) ^ ((fiEnable && (1377 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_13_io_out_valid_0) begin
			b_221_0 <=( _mesh_12_13_io_out_b_0) ^ ((fiEnable && (1378 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_477_0 <=( _mesh_12_13_io_out_c_0) ^ ((fiEnable && (1379 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_13_io_in_control_0_shift_b <=( _mesh_12_13_io_out_control_0_shift) ^ ((fiEnable && (1380 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_13_io_in_control_0_dataflow_b <=( _mesh_12_13_io_out_control_0_dataflow) ^ ((fiEnable && (1381 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_13_io_in_control_0_propagate_b <=( _mesh_12_13_io_out_control_0_propagate) ^ ((fiEnable && (1382 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_13_io_out_valid_0) begin
			b_222_0 <=( _mesh_13_13_io_out_b_0) ^ ((fiEnable && (1383 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_478_0 <=( _mesh_13_13_io_out_c_0) ^ ((fiEnable && (1384 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_13_io_in_control_0_shift_b <=( _mesh_13_13_io_out_control_0_shift) ^ ((fiEnable && (1385 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_13_io_in_control_0_dataflow_b <=( _mesh_13_13_io_out_control_0_dataflow) ^ ((fiEnable && (1386 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_13_io_in_control_0_propagate_b <=( _mesh_13_13_io_out_control_0_propagate) ^ ((fiEnable && (1387 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_13_io_out_valid_0) begin
			b_223_0 <=( _mesh_14_13_io_out_b_0) ^ ((fiEnable && (1388 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_479_0 <=( _mesh_14_13_io_out_c_0) ^ ((fiEnable && (1389 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_13_io_in_control_0_shift_b <=( _mesh_14_13_io_out_control_0_shift) ^ ((fiEnable && (1390 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_13_io_in_control_0_dataflow_b <=( _mesh_14_13_io_out_control_0_dataflow) ^ ((fiEnable && (1391 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_13_io_in_control_0_propagate_b <=( _mesh_14_13_io_out_control_0_propagate) ^ ((fiEnable && (1392 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_14_0) begin
			b_224_0 <=( io_in_b_14_0) ^ ((fiEnable && (1393 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_480_0 <=( io_in_d_14_0) ^ ((fiEnable && (1394 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_14_io_in_control_0_shift_b <=( io_in_control_14_0_shift) ^ ((fiEnable && (1395 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_14_io_in_control_0_dataflow_b <=( io_in_control_14_0_dataflow) ^ ((fiEnable && (1396 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_14_io_in_control_0_propagate_b <=( io_in_control_14_0_propagate) ^ ((fiEnable && (1397 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_14_io_out_valid_0) begin
			b_225_0 <=( _mesh_0_14_io_out_b_0) ^ ((fiEnable && (1398 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_481_0 <=( _mesh_0_14_io_out_c_0) ^ ((fiEnable && (1399 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_14_io_in_control_0_shift_b <=( _mesh_0_14_io_out_control_0_shift) ^ ((fiEnable && (1400 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_14_io_in_control_0_dataflow_b <=( _mesh_0_14_io_out_control_0_dataflow) ^ ((fiEnable && (1401 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_14_io_in_control_0_propagate_b <=( _mesh_0_14_io_out_control_0_propagate) ^ ((fiEnable && (1402 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_14_io_out_valid_0) begin
			b_226_0 <=( _mesh_1_14_io_out_b_0) ^ ((fiEnable && (1403 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_482_0 <=( _mesh_1_14_io_out_c_0) ^ ((fiEnable && (1404 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_14_io_in_control_0_shift_b <=( _mesh_1_14_io_out_control_0_shift) ^ ((fiEnable && (1405 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_14_io_in_control_0_dataflow_b <=( _mesh_1_14_io_out_control_0_dataflow) ^ ((fiEnable && (1406 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_14_io_in_control_0_propagate_b <=( _mesh_1_14_io_out_control_0_propagate) ^ ((fiEnable && (1407 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_14_io_out_valid_0) begin
			b_227_0 <=( _mesh_2_14_io_out_b_0) ^ ((fiEnable && (1408 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_483_0 <=( _mesh_2_14_io_out_c_0) ^ ((fiEnable && (1409 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_14_io_in_control_0_shift_b <=( _mesh_2_14_io_out_control_0_shift) ^ ((fiEnable && (1410 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_14_io_in_control_0_dataflow_b <=( _mesh_2_14_io_out_control_0_dataflow) ^ ((fiEnable && (1411 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_14_io_in_control_0_propagate_b <=( _mesh_2_14_io_out_control_0_propagate) ^ ((fiEnable && (1412 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_14_io_out_valid_0) begin
			b_228_0 <=( _mesh_3_14_io_out_b_0) ^ ((fiEnable && (1413 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_484_0 <=( _mesh_3_14_io_out_c_0) ^ ((fiEnable && (1414 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_14_io_in_control_0_shift_b <=( _mesh_3_14_io_out_control_0_shift) ^ ((fiEnable && (1415 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_14_io_in_control_0_dataflow_b <=( _mesh_3_14_io_out_control_0_dataflow) ^ ((fiEnable && (1416 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_14_io_in_control_0_propagate_b <=( _mesh_3_14_io_out_control_0_propagate) ^ ((fiEnable && (1417 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_14_io_out_valid_0) begin
			b_229_0 <=( _mesh_4_14_io_out_b_0) ^ ((fiEnable && (1418 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_485_0 <=( _mesh_4_14_io_out_c_0) ^ ((fiEnable && (1419 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_14_io_in_control_0_shift_b <=( _mesh_4_14_io_out_control_0_shift) ^ ((fiEnable && (1420 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_14_io_in_control_0_dataflow_b <=( _mesh_4_14_io_out_control_0_dataflow) ^ ((fiEnable && (1421 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_14_io_in_control_0_propagate_b <=( _mesh_4_14_io_out_control_0_propagate) ^ ((fiEnable && (1422 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_14_io_out_valid_0) begin
			b_230_0 <=( _mesh_5_14_io_out_b_0) ^ ((fiEnable && (1423 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_486_0 <=( _mesh_5_14_io_out_c_0) ^ ((fiEnable && (1424 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_14_io_in_control_0_shift_b <=( _mesh_5_14_io_out_control_0_shift) ^ ((fiEnable && (1425 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_14_io_in_control_0_dataflow_b <=( _mesh_5_14_io_out_control_0_dataflow) ^ ((fiEnable && (1426 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_14_io_in_control_0_propagate_b <=( _mesh_5_14_io_out_control_0_propagate) ^ ((fiEnable && (1427 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_14_io_out_valid_0) begin
			b_231_0 <=( _mesh_6_14_io_out_b_0) ^ ((fiEnable && (1428 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_487_0 <=( _mesh_6_14_io_out_c_0) ^ ((fiEnable && (1429 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_14_io_in_control_0_shift_b <=( _mesh_6_14_io_out_control_0_shift) ^ ((fiEnable && (1430 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_14_io_in_control_0_dataflow_b <=( _mesh_6_14_io_out_control_0_dataflow) ^ ((fiEnable && (1431 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_14_io_in_control_0_propagate_b <=( _mesh_6_14_io_out_control_0_propagate) ^ ((fiEnable && (1432 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_14_io_out_valid_0) begin
			b_232_0 <=( _mesh_7_14_io_out_b_0) ^ ((fiEnable && (1433 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_488_0 <=( _mesh_7_14_io_out_c_0) ^ ((fiEnable && (1434 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_14_io_in_control_0_shift_b <=( _mesh_7_14_io_out_control_0_shift) ^ ((fiEnable && (1435 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_14_io_in_control_0_dataflow_b <=( _mesh_7_14_io_out_control_0_dataflow) ^ ((fiEnable && (1436 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_14_io_in_control_0_propagate_b <=( _mesh_7_14_io_out_control_0_propagate) ^ ((fiEnable && (1437 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_14_io_out_valid_0) begin
			b_233_0 <=( _mesh_8_14_io_out_b_0) ^ ((fiEnable && (1438 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_489_0 <=( _mesh_8_14_io_out_c_0) ^ ((fiEnable && (1439 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_14_io_in_control_0_shift_b <=( _mesh_8_14_io_out_control_0_shift) ^ ((fiEnable && (1440 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_14_io_in_control_0_dataflow_b <=( _mesh_8_14_io_out_control_0_dataflow) ^ ((fiEnable && (1441 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_14_io_in_control_0_propagate_b <=( _mesh_8_14_io_out_control_0_propagate) ^ ((fiEnable && (1442 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_14_io_out_valid_0) begin
			b_234_0 <=( _mesh_9_14_io_out_b_0) ^ ((fiEnable && (1443 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_490_0 <=( _mesh_9_14_io_out_c_0) ^ ((fiEnable && (1444 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_14_io_in_control_0_shift_b <=( _mesh_9_14_io_out_control_0_shift) ^ ((fiEnable && (1445 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_14_io_in_control_0_dataflow_b <=( _mesh_9_14_io_out_control_0_dataflow) ^ ((fiEnable && (1446 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_14_io_in_control_0_propagate_b <=( _mesh_9_14_io_out_control_0_propagate) ^ ((fiEnable && (1447 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_14_io_out_valid_0) begin
			b_235_0 <=( _mesh_10_14_io_out_b_0) ^ ((fiEnable && (1448 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_491_0 <=( _mesh_10_14_io_out_c_0) ^ ((fiEnable && (1449 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_14_io_in_control_0_shift_b <=( _mesh_10_14_io_out_control_0_shift) ^ ((fiEnable && (1450 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_14_io_in_control_0_dataflow_b <=( _mesh_10_14_io_out_control_0_dataflow) ^ ((fiEnable && (1451 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_14_io_in_control_0_propagate_b <=( _mesh_10_14_io_out_control_0_propagate) ^ ((fiEnable && (1452 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_14_io_out_valid_0) begin
			b_236_0 <=( _mesh_11_14_io_out_b_0) ^ ((fiEnable && (1453 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_492_0 <=( _mesh_11_14_io_out_c_0) ^ ((fiEnable && (1454 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_14_io_in_control_0_shift_b <=( _mesh_11_14_io_out_control_0_shift) ^ ((fiEnable && (1455 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_14_io_in_control_0_dataflow_b <=( _mesh_11_14_io_out_control_0_dataflow) ^ ((fiEnable && (1456 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_14_io_in_control_0_propagate_b <=( _mesh_11_14_io_out_control_0_propagate) ^ ((fiEnable && (1457 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_14_io_out_valid_0) begin
			b_237_0 <=( _mesh_12_14_io_out_b_0) ^ ((fiEnable && (1458 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_493_0 <=( _mesh_12_14_io_out_c_0) ^ ((fiEnable && (1459 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_14_io_in_control_0_shift_b <=( _mesh_12_14_io_out_control_0_shift) ^ ((fiEnable && (1460 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_14_io_in_control_0_dataflow_b <=( _mesh_12_14_io_out_control_0_dataflow) ^ ((fiEnable && (1461 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_14_io_in_control_0_propagate_b <=( _mesh_12_14_io_out_control_0_propagate) ^ ((fiEnable && (1462 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_14_io_out_valid_0) begin
			b_238_0 <=( _mesh_13_14_io_out_b_0) ^ ((fiEnable && (1463 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_494_0 <=( _mesh_13_14_io_out_c_0) ^ ((fiEnable && (1464 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_14_io_in_control_0_shift_b <=( _mesh_13_14_io_out_control_0_shift) ^ ((fiEnable && (1465 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_14_io_in_control_0_dataflow_b <=( _mesh_13_14_io_out_control_0_dataflow) ^ ((fiEnable && (1466 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_14_io_in_control_0_propagate_b <=( _mesh_13_14_io_out_control_0_propagate) ^ ((fiEnable && (1467 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_14_io_out_valid_0) begin
			b_239_0 <=( _mesh_14_14_io_out_b_0) ^ ((fiEnable && (1468 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_495_0 <=( _mesh_14_14_io_out_c_0) ^ ((fiEnable && (1469 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_14_io_in_control_0_shift_b <=( _mesh_14_14_io_out_control_0_shift) ^ ((fiEnable && (1470 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_14_io_in_control_0_dataflow_b <=( _mesh_14_14_io_out_control_0_dataflow) ^ ((fiEnable && (1471 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_14_io_in_control_0_propagate_b <=( _mesh_14_14_io_out_control_0_propagate) ^ ((fiEnable && (1472 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_15_0) begin
			b_240_0 <=( io_in_b_15_0) ^ ((fiEnable && (1473 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_496_0 <=( io_in_d_15_0) ^ ((fiEnable && (1474 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_15_io_in_control_0_shift_b <=( io_in_control_15_0_shift) ^ ((fiEnable && (1475 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_15_io_in_control_0_dataflow_b <=( io_in_control_15_0_dataflow) ^ ((fiEnable && (1476 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_15_io_in_control_0_propagate_b <=( io_in_control_15_0_propagate) ^ ((fiEnable && (1477 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_15_io_out_valid_0) begin
			b_241_0 <=( _mesh_0_15_io_out_b_0) ^ ((fiEnable && (1478 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_497_0 <=( _mesh_0_15_io_out_c_0) ^ ((fiEnable && (1479 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_15_io_in_control_0_shift_b <=( _mesh_0_15_io_out_control_0_shift) ^ ((fiEnable && (1480 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_15_io_in_control_0_dataflow_b <=( _mesh_0_15_io_out_control_0_dataflow) ^ ((fiEnable && (1481 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_15_io_in_control_0_propagate_b <=( _mesh_0_15_io_out_control_0_propagate) ^ ((fiEnable && (1482 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_15_io_out_valid_0) begin
			b_242_0 <=( _mesh_1_15_io_out_b_0) ^ ((fiEnable && (1483 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_498_0 <=( _mesh_1_15_io_out_c_0) ^ ((fiEnable && (1484 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_15_io_in_control_0_shift_b <=( _mesh_1_15_io_out_control_0_shift) ^ ((fiEnable && (1485 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_15_io_in_control_0_dataflow_b <=( _mesh_1_15_io_out_control_0_dataflow) ^ ((fiEnable && (1486 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_15_io_in_control_0_propagate_b <=( _mesh_1_15_io_out_control_0_propagate) ^ ((fiEnable && (1487 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_15_io_out_valid_0) begin
			b_243_0 <=( _mesh_2_15_io_out_b_0) ^ ((fiEnable && (1488 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_499_0 <=( _mesh_2_15_io_out_c_0) ^ ((fiEnable && (1489 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_15_io_in_control_0_shift_b <=( _mesh_2_15_io_out_control_0_shift) ^ ((fiEnable && (1490 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_15_io_in_control_0_dataflow_b <=( _mesh_2_15_io_out_control_0_dataflow) ^ ((fiEnable && (1491 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_15_io_in_control_0_propagate_b <=( _mesh_2_15_io_out_control_0_propagate) ^ ((fiEnable && (1492 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_15_io_out_valid_0) begin
			b_244_0 <=( _mesh_3_15_io_out_b_0) ^ ((fiEnable && (1493 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_500_0 <=( _mesh_3_15_io_out_c_0) ^ ((fiEnable && (1494 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_15_io_in_control_0_shift_b <=( _mesh_3_15_io_out_control_0_shift) ^ ((fiEnable && (1495 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_15_io_in_control_0_dataflow_b <=( _mesh_3_15_io_out_control_0_dataflow) ^ ((fiEnable && (1496 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_15_io_in_control_0_propagate_b <=( _mesh_3_15_io_out_control_0_propagate) ^ ((fiEnable && (1497 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_15_io_out_valid_0) begin
			b_245_0 <=( _mesh_4_15_io_out_b_0) ^ ((fiEnable && (1498 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_501_0 <=( _mesh_4_15_io_out_c_0) ^ ((fiEnable && (1499 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_15_io_in_control_0_shift_b <=( _mesh_4_15_io_out_control_0_shift) ^ ((fiEnable && (1500 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_15_io_in_control_0_dataflow_b <=( _mesh_4_15_io_out_control_0_dataflow) ^ ((fiEnable && (1501 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_15_io_in_control_0_propagate_b <=( _mesh_4_15_io_out_control_0_propagate) ^ ((fiEnable && (1502 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_15_io_out_valid_0) begin
			b_246_0 <=( _mesh_5_15_io_out_b_0) ^ ((fiEnable && (1503 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_502_0 <=( _mesh_5_15_io_out_c_0) ^ ((fiEnable && (1504 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_15_io_in_control_0_shift_b <=( _mesh_5_15_io_out_control_0_shift) ^ ((fiEnable && (1505 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_15_io_in_control_0_dataflow_b <=( _mesh_5_15_io_out_control_0_dataflow) ^ ((fiEnable && (1506 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_15_io_in_control_0_propagate_b <=( _mesh_5_15_io_out_control_0_propagate) ^ ((fiEnable && (1507 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_15_io_out_valid_0) begin
			b_247_0 <=( _mesh_6_15_io_out_b_0) ^ ((fiEnable && (1508 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_503_0 <=( _mesh_6_15_io_out_c_0) ^ ((fiEnable && (1509 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_15_io_in_control_0_shift_b <=( _mesh_6_15_io_out_control_0_shift) ^ ((fiEnable && (1510 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_15_io_in_control_0_dataflow_b <=( _mesh_6_15_io_out_control_0_dataflow) ^ ((fiEnable && (1511 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_15_io_in_control_0_propagate_b <=( _mesh_6_15_io_out_control_0_propagate) ^ ((fiEnable && (1512 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_15_io_out_valid_0) begin
			b_248_0 <=( _mesh_7_15_io_out_b_0) ^ ((fiEnable && (1513 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_504_0 <=( _mesh_7_15_io_out_c_0) ^ ((fiEnable && (1514 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_15_io_in_control_0_shift_b <=( _mesh_7_15_io_out_control_0_shift) ^ ((fiEnable && (1515 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_15_io_in_control_0_dataflow_b <=( _mesh_7_15_io_out_control_0_dataflow) ^ ((fiEnable && (1516 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_15_io_in_control_0_propagate_b <=( _mesh_7_15_io_out_control_0_propagate) ^ ((fiEnable && (1517 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_15_io_out_valid_0) begin
			b_249_0 <=( _mesh_8_15_io_out_b_0) ^ ((fiEnable && (1518 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_505_0 <=( _mesh_8_15_io_out_c_0) ^ ((fiEnable && (1519 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_15_io_in_control_0_shift_b <=( _mesh_8_15_io_out_control_0_shift) ^ ((fiEnable && (1520 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_15_io_in_control_0_dataflow_b <=( _mesh_8_15_io_out_control_0_dataflow) ^ ((fiEnable && (1521 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_15_io_in_control_0_propagate_b <=( _mesh_8_15_io_out_control_0_propagate) ^ ((fiEnable && (1522 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_15_io_out_valid_0) begin
			b_250_0 <=( _mesh_9_15_io_out_b_0) ^ ((fiEnable && (1523 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_506_0 <=( _mesh_9_15_io_out_c_0) ^ ((fiEnable && (1524 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_15_io_in_control_0_shift_b <=( _mesh_9_15_io_out_control_0_shift) ^ ((fiEnable && (1525 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_15_io_in_control_0_dataflow_b <=( _mesh_9_15_io_out_control_0_dataflow) ^ ((fiEnable && (1526 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_15_io_in_control_0_propagate_b <=( _mesh_9_15_io_out_control_0_propagate) ^ ((fiEnable && (1527 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_15_io_out_valid_0) begin
			b_251_0 <=( _mesh_10_15_io_out_b_0) ^ ((fiEnable && (1528 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_507_0 <=( _mesh_10_15_io_out_c_0) ^ ((fiEnable && (1529 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_15_io_in_control_0_shift_b <=( _mesh_10_15_io_out_control_0_shift) ^ ((fiEnable && (1530 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_15_io_in_control_0_dataflow_b <=( _mesh_10_15_io_out_control_0_dataflow) ^ ((fiEnable && (1531 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_15_io_in_control_0_propagate_b <=( _mesh_10_15_io_out_control_0_propagate) ^ ((fiEnable && (1532 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_15_io_out_valid_0) begin
			b_252_0 <=( _mesh_11_15_io_out_b_0) ^ ((fiEnable && (1533 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_508_0 <=( _mesh_11_15_io_out_c_0) ^ ((fiEnable && (1534 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_15_io_in_control_0_shift_b <=( _mesh_11_15_io_out_control_0_shift) ^ ((fiEnable && (1535 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_15_io_in_control_0_dataflow_b <=( _mesh_11_15_io_out_control_0_dataflow) ^ ((fiEnable && (1536 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_15_io_in_control_0_propagate_b <=( _mesh_11_15_io_out_control_0_propagate) ^ ((fiEnable && (1537 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_15_io_out_valid_0) begin
			b_253_0 <=( _mesh_12_15_io_out_b_0) ^ ((fiEnable && (1538 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_509_0 <=( _mesh_12_15_io_out_c_0) ^ ((fiEnable && (1539 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_15_io_in_control_0_shift_b <=( _mesh_12_15_io_out_control_0_shift) ^ ((fiEnable && (1540 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_15_io_in_control_0_dataflow_b <=( _mesh_12_15_io_out_control_0_dataflow) ^ ((fiEnable && (1541 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_15_io_in_control_0_propagate_b <=( _mesh_12_15_io_out_control_0_propagate) ^ ((fiEnable && (1542 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_15_io_out_valid_0) begin
			b_254_0 <=( _mesh_13_15_io_out_b_0) ^ ((fiEnable && (1543 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_510_0 <=( _mesh_13_15_io_out_c_0) ^ ((fiEnable && (1544 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_15_io_in_control_0_shift_b <=( _mesh_13_15_io_out_control_0_shift) ^ ((fiEnable && (1545 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_15_io_in_control_0_dataflow_b <=( _mesh_13_15_io_out_control_0_dataflow) ^ ((fiEnable && (1546 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_15_io_in_control_0_propagate_b <=( _mesh_13_15_io_out_control_0_propagate) ^ ((fiEnable && (1547 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_15_io_out_valid_0) begin
			b_255_0 <=( _mesh_14_15_io_out_b_0) ^ ((fiEnable && (1548 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_511_0 <=( _mesh_14_15_io_out_c_0) ^ ((fiEnable && (1549 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_15_io_in_control_0_shift_b <=( _mesh_14_15_io_out_control_0_shift) ^ ((fiEnable && (1550 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_15_io_in_control_0_dataflow_b <=( _mesh_14_15_io_out_control_0_dataflow) ^ ((fiEnable && (1551 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_15_io_in_control_0_propagate_b <=( _mesh_14_15_io_out_control_0_propagate) ^ ((fiEnable && (1552 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		r_256_0 <=( io_in_valid_0_0) ^ ((fiEnable && (1553 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_257_0 <=( _mesh_0_0_io_out_valid_0) ^ ((fiEnable && (1554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_258_0 <=( _mesh_1_0_io_out_valid_0) ^ ((fiEnable && (1555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_259_0 <=( _mesh_2_0_io_out_valid_0) ^ ((fiEnable && (1556 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_260_0 <=( _mesh_3_0_io_out_valid_0) ^ ((fiEnable && (1557 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_261_0 <=( _mesh_4_0_io_out_valid_0) ^ ((fiEnable && (1558 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_262_0 <=( _mesh_5_0_io_out_valid_0) ^ ((fiEnable && (1559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_263_0 <=( _mesh_6_0_io_out_valid_0) ^ ((fiEnable && (1560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_264_0 <=( _mesh_7_0_io_out_valid_0) ^ ((fiEnable && (1561 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_265_0 <=( _mesh_8_0_io_out_valid_0) ^ ((fiEnable && (1562 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_266_0 <=( _mesh_9_0_io_out_valid_0) ^ ((fiEnable && (1563 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_267_0 <=( _mesh_10_0_io_out_valid_0) ^ ((fiEnable && (1564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_268_0 <=( _mesh_11_0_io_out_valid_0) ^ ((fiEnable && (1565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_269_0 <=( _mesh_12_0_io_out_valid_0) ^ ((fiEnable && (1566 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_270_0 <=( _mesh_13_0_io_out_valid_0) ^ ((fiEnable && (1567 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_271_0 <=( _mesh_14_0_io_out_valid_0) ^ ((fiEnable && (1568 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_272_0 <=( io_in_valid_1_0) ^ ((fiEnable && (1569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_273_0 <=( _mesh_0_1_io_out_valid_0) ^ ((fiEnable && (1570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_274_0 <=( _mesh_1_1_io_out_valid_0) ^ ((fiEnable && (1571 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_275_0 <=( _mesh_2_1_io_out_valid_0) ^ ((fiEnable && (1572 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_276_0 <=( _mesh_3_1_io_out_valid_0) ^ ((fiEnable && (1573 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_277_0 <=( _mesh_4_1_io_out_valid_0) ^ ((fiEnable && (1574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_278_0 <=( _mesh_5_1_io_out_valid_0) ^ ((fiEnable && (1575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_279_0 <=( _mesh_6_1_io_out_valid_0) ^ ((fiEnable && (1576 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_280_0 <=( _mesh_7_1_io_out_valid_0) ^ ((fiEnable && (1577 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_281_0 <=( _mesh_8_1_io_out_valid_0) ^ ((fiEnable && (1578 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_282_0 <=( _mesh_9_1_io_out_valid_0) ^ ((fiEnable && (1579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_283_0 <=( _mesh_10_1_io_out_valid_0) ^ ((fiEnable && (1580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_284_0 <=( _mesh_11_1_io_out_valid_0) ^ ((fiEnable && (1581 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_285_0 <=( _mesh_12_1_io_out_valid_0) ^ ((fiEnable && (1582 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_286_0 <=( _mesh_13_1_io_out_valid_0) ^ ((fiEnable && (1583 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_287_0 <=( _mesh_14_1_io_out_valid_0) ^ ((fiEnable && (1584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_288_0 <=( io_in_valid_2_0) ^ ((fiEnable && (1585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_289_0 <=( _mesh_0_2_io_out_valid_0) ^ ((fiEnable && (1586 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_290_0 <=( _mesh_1_2_io_out_valid_0) ^ ((fiEnable && (1587 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_291_0 <=( _mesh_2_2_io_out_valid_0) ^ ((fiEnable && (1588 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_292_0 <=( _mesh_3_2_io_out_valid_0) ^ ((fiEnable && (1589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_293_0 <=( _mesh_4_2_io_out_valid_0) ^ ((fiEnable && (1590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_294_0 <=( _mesh_5_2_io_out_valid_0) ^ ((fiEnable && (1591 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_295_0 <=( _mesh_6_2_io_out_valid_0) ^ ((fiEnable && (1592 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_296_0 <=( _mesh_7_2_io_out_valid_0) ^ ((fiEnable && (1593 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_297_0 <=( _mesh_8_2_io_out_valid_0) ^ ((fiEnable && (1594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_298_0 <=( _mesh_9_2_io_out_valid_0) ^ ((fiEnable && (1595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_299_0 <=( _mesh_10_2_io_out_valid_0) ^ ((fiEnable && (1596 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_300_0 <=( _mesh_11_2_io_out_valid_0) ^ ((fiEnable && (1597 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_301_0 <=( _mesh_12_2_io_out_valid_0) ^ ((fiEnable && (1598 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_302_0 <=( _mesh_13_2_io_out_valid_0) ^ ((fiEnable && (1599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_303_0 <=( _mesh_14_2_io_out_valid_0) ^ ((fiEnable && (1600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_304_0 <=( io_in_valid_3_0) ^ ((fiEnable && (1601 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_305_0 <=( _mesh_0_3_io_out_valid_0) ^ ((fiEnable && (1602 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_306_0 <=( _mesh_1_3_io_out_valid_0) ^ ((fiEnable && (1603 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_307_0 <=( _mesh_2_3_io_out_valid_0) ^ ((fiEnable && (1604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_308_0 <=( _mesh_3_3_io_out_valid_0) ^ ((fiEnable && (1605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_309_0 <=( _mesh_4_3_io_out_valid_0) ^ ((fiEnable && (1606 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_310_0 <=( _mesh_5_3_io_out_valid_0) ^ ((fiEnable && (1607 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_311_0 <=( _mesh_6_3_io_out_valid_0) ^ ((fiEnable && (1608 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_312_0 <=( _mesh_7_3_io_out_valid_0) ^ ((fiEnable && (1609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_313_0 <=( _mesh_8_3_io_out_valid_0) ^ ((fiEnable && (1610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_314_0 <=( _mesh_9_3_io_out_valid_0) ^ ((fiEnable && (1611 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_315_0 <=( _mesh_10_3_io_out_valid_0) ^ ((fiEnable && (1612 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_316_0 <=( _mesh_11_3_io_out_valid_0) ^ ((fiEnable && (1613 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_317_0 <=( _mesh_12_3_io_out_valid_0) ^ ((fiEnable && (1614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_318_0 <=( _mesh_13_3_io_out_valid_0) ^ ((fiEnable && (1615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_319_0 <=( _mesh_14_3_io_out_valid_0) ^ ((fiEnable && (1616 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_320_0 <=( io_in_valid_4_0) ^ ((fiEnable && (1617 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_321_0 <=( _mesh_0_4_io_out_valid_0) ^ ((fiEnable && (1618 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_322_0 <=( _mesh_1_4_io_out_valid_0) ^ ((fiEnable && (1619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_323_0 <=( _mesh_2_4_io_out_valid_0) ^ ((fiEnable && (1620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_324_0 <=( _mesh_3_4_io_out_valid_0) ^ ((fiEnable && (1621 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_325_0 <=( _mesh_4_4_io_out_valid_0) ^ ((fiEnable && (1622 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_326_0 <=( _mesh_5_4_io_out_valid_0) ^ ((fiEnable && (1623 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_327_0 <=( _mesh_6_4_io_out_valid_0) ^ ((fiEnable && (1624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_328_0 <=( _mesh_7_4_io_out_valid_0) ^ ((fiEnable && (1625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_329_0 <=( _mesh_8_4_io_out_valid_0) ^ ((fiEnable && (1626 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_330_0 <=( _mesh_9_4_io_out_valid_0) ^ ((fiEnable && (1627 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_331_0 <=( _mesh_10_4_io_out_valid_0) ^ ((fiEnable && (1628 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_332_0 <=( _mesh_11_4_io_out_valid_0) ^ ((fiEnable && (1629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_333_0 <=( _mesh_12_4_io_out_valid_0) ^ ((fiEnable && (1630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_334_0 <=( _mesh_13_4_io_out_valid_0) ^ ((fiEnable && (1631 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_335_0 <=( _mesh_14_4_io_out_valid_0) ^ ((fiEnable && (1632 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_336_0 <=( io_in_valid_5_0) ^ ((fiEnable && (1633 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_337_0 <=( _mesh_0_5_io_out_valid_0) ^ ((fiEnable && (1634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_338_0 <=( _mesh_1_5_io_out_valid_0) ^ ((fiEnable && (1635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_339_0 <=( _mesh_2_5_io_out_valid_0) ^ ((fiEnable && (1636 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_340_0 <=( _mesh_3_5_io_out_valid_0) ^ ((fiEnable && (1637 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_341_0 <=( _mesh_4_5_io_out_valid_0) ^ ((fiEnable && (1638 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_342_0 <=( _mesh_5_5_io_out_valid_0) ^ ((fiEnable && (1639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_343_0 <=( _mesh_6_5_io_out_valid_0) ^ ((fiEnable && (1640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_344_0 <=( _mesh_7_5_io_out_valid_0) ^ ((fiEnable && (1641 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_345_0 <=( _mesh_8_5_io_out_valid_0) ^ ((fiEnable && (1642 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_346_0 <=( _mesh_9_5_io_out_valid_0) ^ ((fiEnable && (1643 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_347_0 <=( _mesh_10_5_io_out_valid_0) ^ ((fiEnable && (1644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_348_0 <=( _mesh_11_5_io_out_valid_0) ^ ((fiEnable && (1645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_349_0 <=( _mesh_12_5_io_out_valid_0) ^ ((fiEnable && (1646 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_350_0 <=( _mesh_13_5_io_out_valid_0) ^ ((fiEnable && (1647 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_351_0 <=( _mesh_14_5_io_out_valid_0) ^ ((fiEnable && (1648 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_352_0 <=( io_in_valid_6_0) ^ ((fiEnable && (1649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_353_0 <=( _mesh_0_6_io_out_valid_0) ^ ((fiEnable && (1650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_354_0 <=( _mesh_1_6_io_out_valid_0) ^ ((fiEnable && (1651 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_355_0 <=( _mesh_2_6_io_out_valid_0) ^ ((fiEnable && (1652 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_356_0 <=( _mesh_3_6_io_out_valid_0) ^ ((fiEnable && (1653 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_357_0 <=( _mesh_4_6_io_out_valid_0) ^ ((fiEnable && (1654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_358_0 <=( _mesh_5_6_io_out_valid_0) ^ ((fiEnable && (1655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_359_0 <=( _mesh_6_6_io_out_valid_0) ^ ((fiEnable && (1656 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_360_0 <=( _mesh_7_6_io_out_valid_0) ^ ((fiEnable && (1657 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_361_0 <=( _mesh_8_6_io_out_valid_0) ^ ((fiEnable && (1658 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_362_0 <=( _mesh_9_6_io_out_valid_0) ^ ((fiEnable && (1659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_363_0 <=( _mesh_10_6_io_out_valid_0) ^ ((fiEnable && (1660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_364_0 <=( _mesh_11_6_io_out_valid_0) ^ ((fiEnable && (1661 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_365_0 <=( _mesh_12_6_io_out_valid_0) ^ ((fiEnable && (1662 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_366_0 <=( _mesh_13_6_io_out_valid_0) ^ ((fiEnable && (1663 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_367_0 <=( _mesh_14_6_io_out_valid_0) ^ ((fiEnable && (1664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_368_0 <=( io_in_valid_7_0) ^ ((fiEnable && (1665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_369_0 <=( _mesh_0_7_io_out_valid_0) ^ ((fiEnable && (1666 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_370_0 <=( _mesh_1_7_io_out_valid_0) ^ ((fiEnable && (1667 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_371_0 <=( _mesh_2_7_io_out_valid_0) ^ ((fiEnable && (1668 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_372_0 <=( _mesh_3_7_io_out_valid_0) ^ ((fiEnable && (1669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_373_0 <=( _mesh_4_7_io_out_valid_0) ^ ((fiEnable && (1670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_374_0 <=( _mesh_5_7_io_out_valid_0) ^ ((fiEnable && (1671 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_375_0 <=( _mesh_6_7_io_out_valid_0) ^ ((fiEnable && (1672 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_376_0 <=( _mesh_7_7_io_out_valid_0) ^ ((fiEnable && (1673 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_377_0 <=( _mesh_8_7_io_out_valid_0) ^ ((fiEnable && (1674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_378_0 <=( _mesh_9_7_io_out_valid_0) ^ ((fiEnable && (1675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_379_0 <=( _mesh_10_7_io_out_valid_0) ^ ((fiEnable && (1676 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_380_0 <=( _mesh_11_7_io_out_valid_0) ^ ((fiEnable && (1677 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_381_0 <=( _mesh_12_7_io_out_valid_0) ^ ((fiEnable && (1678 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_382_0 <=( _mesh_13_7_io_out_valid_0) ^ ((fiEnable && (1679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_383_0 <=( _mesh_14_7_io_out_valid_0) ^ ((fiEnable && (1680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_384_0 <=( io_in_valid_8_0) ^ ((fiEnable && (1681 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_385_0 <=( _mesh_0_8_io_out_valid_0) ^ ((fiEnable && (1682 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_386_0 <=( _mesh_1_8_io_out_valid_0) ^ ((fiEnable && (1683 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_387_0 <=( _mesh_2_8_io_out_valid_0) ^ ((fiEnable && (1684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_388_0 <=( _mesh_3_8_io_out_valid_0) ^ ((fiEnable && (1685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_389_0 <=( _mesh_4_8_io_out_valid_0) ^ ((fiEnable && (1686 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_390_0 <=( _mesh_5_8_io_out_valid_0) ^ ((fiEnable && (1687 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_391_0 <=( _mesh_6_8_io_out_valid_0) ^ ((fiEnable && (1688 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_392_0 <=( _mesh_7_8_io_out_valid_0) ^ ((fiEnable && (1689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_393_0 <=( _mesh_8_8_io_out_valid_0) ^ ((fiEnable && (1690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_394_0 <=( _mesh_9_8_io_out_valid_0) ^ ((fiEnable && (1691 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_395_0 <=( _mesh_10_8_io_out_valid_0) ^ ((fiEnable && (1692 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_396_0 <=( _mesh_11_8_io_out_valid_0) ^ ((fiEnable && (1693 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_397_0 <=( _mesh_12_8_io_out_valid_0) ^ ((fiEnable && (1694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_398_0 <=( _mesh_13_8_io_out_valid_0) ^ ((fiEnable && (1695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_399_0 <=( _mesh_14_8_io_out_valid_0) ^ ((fiEnable && (1696 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_400_0 <=( io_in_valid_9_0) ^ ((fiEnable && (1697 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_401_0 <=( _mesh_0_9_io_out_valid_0) ^ ((fiEnable && (1698 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_402_0 <=( _mesh_1_9_io_out_valid_0) ^ ((fiEnable && (1699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_403_0 <=( _mesh_2_9_io_out_valid_0) ^ ((fiEnable && (1700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_404_0 <=( _mesh_3_9_io_out_valid_0) ^ ((fiEnable && (1701 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_405_0 <=( _mesh_4_9_io_out_valid_0) ^ ((fiEnable && (1702 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_406_0 <=( _mesh_5_9_io_out_valid_0) ^ ((fiEnable && (1703 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_407_0 <=( _mesh_6_9_io_out_valid_0) ^ ((fiEnable && (1704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_408_0 <=( _mesh_7_9_io_out_valid_0) ^ ((fiEnable && (1705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_409_0 <=( _mesh_8_9_io_out_valid_0) ^ ((fiEnable && (1706 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_410_0 <=( _mesh_9_9_io_out_valid_0) ^ ((fiEnable && (1707 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_411_0 <=( _mesh_10_9_io_out_valid_0) ^ ((fiEnable && (1708 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_412_0 <=( _mesh_11_9_io_out_valid_0) ^ ((fiEnable && (1709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_413_0 <=( _mesh_12_9_io_out_valid_0) ^ ((fiEnable && (1710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_414_0 <=( _mesh_13_9_io_out_valid_0) ^ ((fiEnable && (1711 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_415_0 <=( _mesh_14_9_io_out_valid_0) ^ ((fiEnable && (1712 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_416_0 <=( io_in_valid_10_0) ^ ((fiEnable && (1713 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_417_0 <=( _mesh_0_10_io_out_valid_0) ^ ((fiEnable && (1714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_418_0 <=( _mesh_1_10_io_out_valid_0) ^ ((fiEnable && (1715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_419_0 <=( _mesh_2_10_io_out_valid_0) ^ ((fiEnable && (1716 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_420_0 <=( _mesh_3_10_io_out_valid_0) ^ ((fiEnable && (1717 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_421_0 <=( _mesh_4_10_io_out_valid_0) ^ ((fiEnable && (1718 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_422_0 <=( _mesh_5_10_io_out_valid_0) ^ ((fiEnable && (1719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_423_0 <=( _mesh_6_10_io_out_valid_0) ^ ((fiEnable && (1720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_424_0 <=( _mesh_7_10_io_out_valid_0) ^ ((fiEnable && (1721 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_425_0 <=( _mesh_8_10_io_out_valid_0) ^ ((fiEnable && (1722 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_426_0 <=( _mesh_9_10_io_out_valid_0) ^ ((fiEnable && (1723 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_427_0 <=( _mesh_10_10_io_out_valid_0) ^ ((fiEnable && (1724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_428_0 <=( _mesh_11_10_io_out_valid_0) ^ ((fiEnable && (1725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_429_0 <=( _mesh_12_10_io_out_valid_0) ^ ((fiEnable && (1726 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_430_0 <=( _mesh_13_10_io_out_valid_0) ^ ((fiEnable && (1727 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_431_0 <=( _mesh_14_10_io_out_valid_0) ^ ((fiEnable && (1728 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_432_0 <=( io_in_valid_11_0) ^ ((fiEnable && (1729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_433_0 <=( _mesh_0_11_io_out_valid_0) ^ ((fiEnable && (1730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_434_0 <=( _mesh_1_11_io_out_valid_0) ^ ((fiEnable && (1731 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_435_0 <=( _mesh_2_11_io_out_valid_0) ^ ((fiEnable && (1732 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_436_0 <=( _mesh_3_11_io_out_valid_0) ^ ((fiEnable && (1733 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_437_0 <=( _mesh_4_11_io_out_valid_0) ^ ((fiEnable && (1734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_438_0 <=( _mesh_5_11_io_out_valid_0) ^ ((fiEnable && (1735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_439_0 <=( _mesh_6_11_io_out_valid_0) ^ ((fiEnable && (1736 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_440_0 <=( _mesh_7_11_io_out_valid_0) ^ ((fiEnable && (1737 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_441_0 <=( _mesh_8_11_io_out_valid_0) ^ ((fiEnable && (1738 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_442_0 <=( _mesh_9_11_io_out_valid_0) ^ ((fiEnable && (1739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_443_0 <=( _mesh_10_11_io_out_valid_0) ^ ((fiEnable && (1740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_444_0 <=( _mesh_11_11_io_out_valid_0) ^ ((fiEnable && (1741 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_445_0 <=( _mesh_12_11_io_out_valid_0) ^ ((fiEnable && (1742 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_446_0 <=( _mesh_13_11_io_out_valid_0) ^ ((fiEnable && (1743 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_447_0 <=( _mesh_14_11_io_out_valid_0) ^ ((fiEnable && (1744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_448_0 <=( io_in_valid_12_0) ^ ((fiEnable && (1745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_449_0 <=( _mesh_0_12_io_out_valid_0) ^ ((fiEnable && (1746 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_450_0 <=( _mesh_1_12_io_out_valid_0) ^ ((fiEnable && (1747 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_451_0 <=( _mesh_2_12_io_out_valid_0) ^ ((fiEnable && (1748 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_452_0 <=( _mesh_3_12_io_out_valid_0) ^ ((fiEnable && (1749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_453_0 <=( _mesh_4_12_io_out_valid_0) ^ ((fiEnable && (1750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_454_0 <=( _mesh_5_12_io_out_valid_0) ^ ((fiEnable && (1751 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_455_0 <=( _mesh_6_12_io_out_valid_0) ^ ((fiEnable && (1752 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_456_0 <=( _mesh_7_12_io_out_valid_0) ^ ((fiEnable && (1753 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_457_0 <=( _mesh_8_12_io_out_valid_0) ^ ((fiEnable && (1754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_458_0 <=( _mesh_9_12_io_out_valid_0) ^ ((fiEnable && (1755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_459_0 <=( _mesh_10_12_io_out_valid_0) ^ ((fiEnable && (1756 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_460_0 <=( _mesh_11_12_io_out_valid_0) ^ ((fiEnable && (1757 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_461_0 <=( _mesh_12_12_io_out_valid_0) ^ ((fiEnable && (1758 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_462_0 <=( _mesh_13_12_io_out_valid_0) ^ ((fiEnable && (1759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_463_0 <=( _mesh_14_12_io_out_valid_0) ^ ((fiEnable && (1760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_464_0 <=( io_in_valid_13_0) ^ ((fiEnable && (1761 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_465_0 <=( _mesh_0_13_io_out_valid_0) ^ ((fiEnable && (1762 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_466_0 <=( _mesh_1_13_io_out_valid_0) ^ ((fiEnable && (1763 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_467_0 <=( _mesh_2_13_io_out_valid_0) ^ ((fiEnable && (1764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_468_0 <=( _mesh_3_13_io_out_valid_0) ^ ((fiEnable && (1765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_469_0 <=( _mesh_4_13_io_out_valid_0) ^ ((fiEnable && (1766 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_470_0 <=( _mesh_5_13_io_out_valid_0) ^ ((fiEnable && (1767 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_471_0 <=( _mesh_6_13_io_out_valid_0) ^ ((fiEnable && (1768 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_472_0 <=( _mesh_7_13_io_out_valid_0) ^ ((fiEnable && (1769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_473_0 <=( _mesh_8_13_io_out_valid_0) ^ ((fiEnable && (1770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_474_0 <=( _mesh_9_13_io_out_valid_0) ^ ((fiEnable && (1771 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_475_0 <=( _mesh_10_13_io_out_valid_0) ^ ((fiEnable && (1772 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_476_0 <=( _mesh_11_13_io_out_valid_0) ^ ((fiEnable && (1773 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_477_0 <=( _mesh_12_13_io_out_valid_0) ^ ((fiEnable && (1774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_478_0 <=( _mesh_13_13_io_out_valid_0) ^ ((fiEnable && (1775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_479_0 <=( _mesh_14_13_io_out_valid_0) ^ ((fiEnable && (1776 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_480_0 <=( io_in_valid_14_0) ^ ((fiEnable && (1777 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_481_0 <=( _mesh_0_14_io_out_valid_0) ^ ((fiEnable && (1778 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_482_0 <=( _mesh_1_14_io_out_valid_0) ^ ((fiEnable && (1779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_483_0 <=( _mesh_2_14_io_out_valid_0) ^ ((fiEnable && (1780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_484_0 <=( _mesh_3_14_io_out_valid_0) ^ ((fiEnable && (1781 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_485_0 <=( _mesh_4_14_io_out_valid_0) ^ ((fiEnable && (1782 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_486_0 <=( _mesh_5_14_io_out_valid_0) ^ ((fiEnable && (1783 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_487_0 <=( _mesh_6_14_io_out_valid_0) ^ ((fiEnable && (1784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_488_0 <=( _mesh_7_14_io_out_valid_0) ^ ((fiEnable && (1785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_489_0 <=( _mesh_8_14_io_out_valid_0) ^ ((fiEnable && (1786 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_490_0 <=( _mesh_9_14_io_out_valid_0) ^ ((fiEnable && (1787 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_491_0 <=( _mesh_10_14_io_out_valid_0) ^ ((fiEnable && (1788 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_492_0 <=( _mesh_11_14_io_out_valid_0) ^ ((fiEnable && (1789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_493_0 <=( _mesh_12_14_io_out_valid_0) ^ ((fiEnable && (1790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_494_0 <=( _mesh_13_14_io_out_valid_0) ^ ((fiEnable && (1791 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_495_0 <=( _mesh_14_14_io_out_valid_0) ^ ((fiEnable && (1792 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_496_0 <=( io_in_valid_15_0) ^ ((fiEnable && (1793 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_497_0 <=( _mesh_0_15_io_out_valid_0) ^ ((fiEnable && (1794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_498_0 <=( _mesh_1_15_io_out_valid_0) ^ ((fiEnable && (1795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_499_0 <=( _mesh_2_15_io_out_valid_0) ^ ((fiEnable && (1796 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_500_0 <=( _mesh_3_15_io_out_valid_0) ^ ((fiEnable && (1797 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_501_0 <=( _mesh_4_15_io_out_valid_0) ^ ((fiEnable && (1798 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_502_0 <=( _mesh_5_15_io_out_valid_0) ^ ((fiEnable && (1799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_503_0 <=( _mesh_6_15_io_out_valid_0) ^ ((fiEnable && (1800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_504_0 <=( _mesh_7_15_io_out_valid_0) ^ ((fiEnable && (1801 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_505_0 <=( _mesh_8_15_io_out_valid_0) ^ ((fiEnable && (1802 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_506_0 <=( _mesh_9_15_io_out_valid_0) ^ ((fiEnable && (1803 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_507_0 <=( _mesh_10_15_io_out_valid_0) ^ ((fiEnable && (1804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_508_0 <=( _mesh_11_15_io_out_valid_0) ^ ((fiEnable && (1805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_509_0 <=( _mesh_12_15_io_out_valid_0) ^ ((fiEnable && (1806 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_510_0 <=( _mesh_13_15_io_out_valid_0) ^ ((fiEnable && (1807 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_511_0 <=( _mesh_14_15_io_out_valid_0) ^ ((fiEnable && (1808 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_512_0 <=( io_in_id_0_0) ^ ((fiEnable && (1809 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_513_0 <=( _mesh_0_0_io_out_id_0) ^ ((fiEnable && (1810 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_514_0 <=( _mesh_1_0_io_out_id_0) ^ ((fiEnable && (1811 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_515_0 <=( _mesh_2_0_io_out_id_0) ^ ((fiEnable && (1812 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_516_0 <=( _mesh_3_0_io_out_id_0) ^ ((fiEnable && (1813 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_517_0 <=( _mesh_4_0_io_out_id_0) ^ ((fiEnable && (1814 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_518_0 <=( _mesh_5_0_io_out_id_0) ^ ((fiEnable && (1815 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_519_0 <=( _mesh_6_0_io_out_id_0) ^ ((fiEnable && (1816 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_520_0 <=( _mesh_7_0_io_out_id_0) ^ ((fiEnable && (1817 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_521_0 <=( _mesh_8_0_io_out_id_0) ^ ((fiEnable && (1818 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_522_0 <=( _mesh_9_0_io_out_id_0) ^ ((fiEnable && (1819 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_523_0 <=( _mesh_10_0_io_out_id_0) ^ ((fiEnable && (1820 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_524_0 <=( _mesh_11_0_io_out_id_0) ^ ((fiEnable && (1821 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_525_0 <=( _mesh_12_0_io_out_id_0) ^ ((fiEnable && (1822 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_526_0 <=( _mesh_13_0_io_out_id_0) ^ ((fiEnable && (1823 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_527_0 <=( _mesh_14_0_io_out_id_0) ^ ((fiEnable && (1824 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_528_0 <=( io_in_id_1_0) ^ ((fiEnable && (1825 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_529_0 <=( _mesh_0_1_io_out_id_0) ^ ((fiEnable && (1826 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_530_0 <=( _mesh_1_1_io_out_id_0) ^ ((fiEnable && (1827 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_531_0 <=( _mesh_2_1_io_out_id_0) ^ ((fiEnable && (1828 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_532_0 <=( _mesh_3_1_io_out_id_0) ^ ((fiEnable && (1829 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_533_0 <=( _mesh_4_1_io_out_id_0) ^ ((fiEnable && (1830 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_534_0 <=( _mesh_5_1_io_out_id_0) ^ ((fiEnable && (1831 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_535_0 <=( _mesh_6_1_io_out_id_0) ^ ((fiEnable && (1832 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_536_0 <=( _mesh_7_1_io_out_id_0) ^ ((fiEnable && (1833 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_537_0 <=( _mesh_8_1_io_out_id_0) ^ ((fiEnable && (1834 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_538_0 <=( _mesh_9_1_io_out_id_0) ^ ((fiEnable && (1835 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_539_0 <=( _mesh_10_1_io_out_id_0) ^ ((fiEnable && (1836 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_540_0 <=( _mesh_11_1_io_out_id_0) ^ ((fiEnable && (1837 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_541_0 <=( _mesh_12_1_io_out_id_0) ^ ((fiEnable && (1838 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_542_0 <=( _mesh_13_1_io_out_id_0) ^ ((fiEnable && (1839 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_543_0 <=( _mesh_14_1_io_out_id_0) ^ ((fiEnable && (1840 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_544_0 <=( io_in_id_2_0) ^ ((fiEnable && (1841 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_545_0 <=( _mesh_0_2_io_out_id_0) ^ ((fiEnable && (1842 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_546_0 <=( _mesh_1_2_io_out_id_0) ^ ((fiEnable && (1843 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_547_0 <=( _mesh_2_2_io_out_id_0) ^ ((fiEnable && (1844 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_548_0 <=( _mesh_3_2_io_out_id_0) ^ ((fiEnable && (1845 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_549_0 <=( _mesh_4_2_io_out_id_0) ^ ((fiEnable && (1846 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_550_0 <=( _mesh_5_2_io_out_id_0) ^ ((fiEnable && (1847 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_551_0 <=( _mesh_6_2_io_out_id_0) ^ ((fiEnable && (1848 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_552_0 <=( _mesh_7_2_io_out_id_0) ^ ((fiEnable && (1849 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_553_0 <=( _mesh_8_2_io_out_id_0) ^ ((fiEnable && (1850 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_554_0 <=( _mesh_9_2_io_out_id_0) ^ ((fiEnable && (1851 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_555_0 <=( _mesh_10_2_io_out_id_0) ^ ((fiEnable && (1852 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_556_0 <=( _mesh_11_2_io_out_id_0) ^ ((fiEnable && (1853 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_557_0 <=( _mesh_12_2_io_out_id_0) ^ ((fiEnable && (1854 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_558_0 <=( _mesh_13_2_io_out_id_0) ^ ((fiEnable && (1855 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_559_0 <=( _mesh_14_2_io_out_id_0) ^ ((fiEnable && (1856 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_560_0 <=( io_in_id_3_0) ^ ((fiEnable && (1857 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_561_0 <=( _mesh_0_3_io_out_id_0) ^ ((fiEnable && (1858 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_562_0 <=( _mesh_1_3_io_out_id_0) ^ ((fiEnable && (1859 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_563_0 <=( _mesh_2_3_io_out_id_0) ^ ((fiEnable && (1860 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_564_0 <=( _mesh_3_3_io_out_id_0) ^ ((fiEnable && (1861 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_565_0 <=( _mesh_4_3_io_out_id_0) ^ ((fiEnable && (1862 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_566_0 <=( _mesh_5_3_io_out_id_0) ^ ((fiEnable && (1863 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_567_0 <=( _mesh_6_3_io_out_id_0) ^ ((fiEnable && (1864 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_568_0 <=( _mesh_7_3_io_out_id_0) ^ ((fiEnable && (1865 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_569_0 <=( _mesh_8_3_io_out_id_0) ^ ((fiEnable && (1866 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_570_0 <=( _mesh_9_3_io_out_id_0) ^ ((fiEnable && (1867 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_571_0 <=( _mesh_10_3_io_out_id_0) ^ ((fiEnable && (1868 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_572_0 <=( _mesh_11_3_io_out_id_0) ^ ((fiEnable && (1869 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_573_0 <=( _mesh_12_3_io_out_id_0) ^ ((fiEnable && (1870 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_574_0 <=( _mesh_13_3_io_out_id_0) ^ ((fiEnable && (1871 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_575_0 <=( _mesh_14_3_io_out_id_0) ^ ((fiEnable && (1872 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_576_0 <=( io_in_id_4_0) ^ ((fiEnable && (1873 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_577_0 <=( _mesh_0_4_io_out_id_0) ^ ((fiEnable && (1874 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_578_0 <=( _mesh_1_4_io_out_id_0) ^ ((fiEnable && (1875 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_579_0 <=( _mesh_2_4_io_out_id_0) ^ ((fiEnable && (1876 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_580_0 <=( _mesh_3_4_io_out_id_0) ^ ((fiEnable && (1877 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_581_0 <=( _mesh_4_4_io_out_id_0) ^ ((fiEnable && (1878 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_582_0 <=( _mesh_5_4_io_out_id_0) ^ ((fiEnable && (1879 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_583_0 <=( _mesh_6_4_io_out_id_0) ^ ((fiEnable && (1880 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_584_0 <=( _mesh_7_4_io_out_id_0) ^ ((fiEnable && (1881 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_585_0 <=( _mesh_8_4_io_out_id_0) ^ ((fiEnable && (1882 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_586_0 <=( _mesh_9_4_io_out_id_0) ^ ((fiEnable && (1883 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_587_0 <=( _mesh_10_4_io_out_id_0) ^ ((fiEnable && (1884 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_588_0 <=( _mesh_11_4_io_out_id_0) ^ ((fiEnable && (1885 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_589_0 <=( _mesh_12_4_io_out_id_0) ^ ((fiEnable && (1886 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_590_0 <=( _mesh_13_4_io_out_id_0) ^ ((fiEnable && (1887 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_591_0 <=( _mesh_14_4_io_out_id_0) ^ ((fiEnable && (1888 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_592_0 <=( io_in_id_5_0) ^ ((fiEnable && (1889 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_593_0 <=( _mesh_0_5_io_out_id_0) ^ ((fiEnable && (1890 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_594_0 <=( _mesh_1_5_io_out_id_0) ^ ((fiEnable && (1891 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_595_0 <=( _mesh_2_5_io_out_id_0) ^ ((fiEnable && (1892 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_596_0 <=( _mesh_3_5_io_out_id_0) ^ ((fiEnable && (1893 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_597_0 <=( _mesh_4_5_io_out_id_0) ^ ((fiEnable && (1894 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_598_0 <=( _mesh_5_5_io_out_id_0) ^ ((fiEnable && (1895 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_599_0 <=( _mesh_6_5_io_out_id_0) ^ ((fiEnable && (1896 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_600_0 <=( _mesh_7_5_io_out_id_0) ^ ((fiEnable && (1897 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_601_0 <=( _mesh_8_5_io_out_id_0) ^ ((fiEnable && (1898 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_602_0 <=( _mesh_9_5_io_out_id_0) ^ ((fiEnable && (1899 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_603_0 <=( _mesh_10_5_io_out_id_0) ^ ((fiEnable && (1900 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_604_0 <=( _mesh_11_5_io_out_id_0) ^ ((fiEnable && (1901 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_605_0 <=( _mesh_12_5_io_out_id_0) ^ ((fiEnable && (1902 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_606_0 <=( _mesh_13_5_io_out_id_0) ^ ((fiEnable && (1903 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_607_0 <=( _mesh_14_5_io_out_id_0) ^ ((fiEnable && (1904 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_608_0 <=( io_in_id_6_0) ^ ((fiEnable && (1905 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_609_0 <=( _mesh_0_6_io_out_id_0) ^ ((fiEnable && (1906 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_610_0 <=( _mesh_1_6_io_out_id_0) ^ ((fiEnable && (1907 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_611_0 <=( _mesh_2_6_io_out_id_0) ^ ((fiEnable && (1908 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_612_0 <=( _mesh_3_6_io_out_id_0) ^ ((fiEnable && (1909 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_613_0 <=( _mesh_4_6_io_out_id_0) ^ ((fiEnable && (1910 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_614_0 <=( _mesh_5_6_io_out_id_0) ^ ((fiEnable && (1911 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_615_0 <=( _mesh_6_6_io_out_id_0) ^ ((fiEnable && (1912 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_616_0 <=( _mesh_7_6_io_out_id_0) ^ ((fiEnable && (1913 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_617_0 <=( _mesh_8_6_io_out_id_0) ^ ((fiEnable && (1914 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_618_0 <=( _mesh_9_6_io_out_id_0) ^ ((fiEnable && (1915 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_619_0 <=( _mesh_10_6_io_out_id_0) ^ ((fiEnable && (1916 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_620_0 <=( _mesh_11_6_io_out_id_0) ^ ((fiEnable && (1917 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_621_0 <=( _mesh_12_6_io_out_id_0) ^ ((fiEnable && (1918 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_622_0 <=( _mesh_13_6_io_out_id_0) ^ ((fiEnable && (1919 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_623_0 <=( _mesh_14_6_io_out_id_0) ^ ((fiEnable && (1920 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_624_0 <=( io_in_id_7_0) ^ ((fiEnable && (1921 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_625_0 <=( _mesh_0_7_io_out_id_0) ^ ((fiEnable && (1922 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_626_0 <=( _mesh_1_7_io_out_id_0) ^ ((fiEnable && (1923 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_627_0 <=( _mesh_2_7_io_out_id_0) ^ ((fiEnable && (1924 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_628_0 <=( _mesh_3_7_io_out_id_0) ^ ((fiEnable && (1925 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_629_0 <=( _mesh_4_7_io_out_id_0) ^ ((fiEnable && (1926 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_630_0 <=( _mesh_5_7_io_out_id_0) ^ ((fiEnable && (1927 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_631_0 <=( _mesh_6_7_io_out_id_0) ^ ((fiEnable && (1928 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_632_0 <=( _mesh_7_7_io_out_id_0) ^ ((fiEnable && (1929 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_633_0 <=( _mesh_8_7_io_out_id_0) ^ ((fiEnable && (1930 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_634_0 <=( _mesh_9_7_io_out_id_0) ^ ((fiEnable && (1931 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_635_0 <=( _mesh_10_7_io_out_id_0) ^ ((fiEnable && (1932 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_636_0 <=( _mesh_11_7_io_out_id_0) ^ ((fiEnable && (1933 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_637_0 <=( _mesh_12_7_io_out_id_0) ^ ((fiEnable && (1934 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_638_0 <=( _mesh_13_7_io_out_id_0) ^ ((fiEnable && (1935 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_639_0 <=( _mesh_14_7_io_out_id_0) ^ ((fiEnable && (1936 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_640_0 <=( io_in_id_8_0) ^ ((fiEnable && (1937 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_641_0 <=( _mesh_0_8_io_out_id_0) ^ ((fiEnable && (1938 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_642_0 <=( _mesh_1_8_io_out_id_0) ^ ((fiEnable && (1939 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_643_0 <=( _mesh_2_8_io_out_id_0) ^ ((fiEnable && (1940 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_644_0 <=( _mesh_3_8_io_out_id_0) ^ ((fiEnable && (1941 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_645_0 <=( _mesh_4_8_io_out_id_0) ^ ((fiEnable && (1942 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_646_0 <=( _mesh_5_8_io_out_id_0) ^ ((fiEnable && (1943 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_647_0 <=( _mesh_6_8_io_out_id_0) ^ ((fiEnable && (1944 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_648_0 <=( _mesh_7_8_io_out_id_0) ^ ((fiEnable && (1945 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_649_0 <=( _mesh_8_8_io_out_id_0) ^ ((fiEnable && (1946 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_650_0 <=( _mesh_9_8_io_out_id_0) ^ ((fiEnable && (1947 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_651_0 <=( _mesh_10_8_io_out_id_0) ^ ((fiEnable && (1948 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_652_0 <=( _mesh_11_8_io_out_id_0) ^ ((fiEnable && (1949 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_653_0 <=( _mesh_12_8_io_out_id_0) ^ ((fiEnable && (1950 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_654_0 <=( _mesh_13_8_io_out_id_0) ^ ((fiEnable && (1951 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_655_0 <=( _mesh_14_8_io_out_id_0) ^ ((fiEnable && (1952 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_656_0 <=( io_in_id_9_0) ^ ((fiEnable && (1953 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_657_0 <=( _mesh_0_9_io_out_id_0) ^ ((fiEnable && (1954 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_658_0 <=( _mesh_1_9_io_out_id_0) ^ ((fiEnable && (1955 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_659_0 <=( _mesh_2_9_io_out_id_0) ^ ((fiEnable && (1956 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_660_0 <=( _mesh_3_9_io_out_id_0) ^ ((fiEnable && (1957 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_661_0 <=( _mesh_4_9_io_out_id_0) ^ ((fiEnable && (1958 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_662_0 <=( _mesh_5_9_io_out_id_0) ^ ((fiEnable && (1959 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_663_0 <=( _mesh_6_9_io_out_id_0) ^ ((fiEnable && (1960 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_664_0 <=( _mesh_7_9_io_out_id_0) ^ ((fiEnable && (1961 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_665_0 <=( _mesh_8_9_io_out_id_0) ^ ((fiEnable && (1962 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_666_0 <=( _mesh_9_9_io_out_id_0) ^ ((fiEnable && (1963 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_667_0 <=( _mesh_10_9_io_out_id_0) ^ ((fiEnable && (1964 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_668_0 <=( _mesh_11_9_io_out_id_0) ^ ((fiEnable && (1965 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_669_0 <=( _mesh_12_9_io_out_id_0) ^ ((fiEnable && (1966 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_670_0 <=( _mesh_13_9_io_out_id_0) ^ ((fiEnable && (1967 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_671_0 <=( _mesh_14_9_io_out_id_0) ^ ((fiEnable && (1968 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_672_0 <=( io_in_id_10_0) ^ ((fiEnable && (1969 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_673_0 <=( _mesh_0_10_io_out_id_0) ^ ((fiEnable && (1970 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_674_0 <=( _mesh_1_10_io_out_id_0) ^ ((fiEnable && (1971 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_675_0 <=( _mesh_2_10_io_out_id_0) ^ ((fiEnable && (1972 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_676_0 <=( _mesh_3_10_io_out_id_0) ^ ((fiEnable && (1973 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_677_0 <=( _mesh_4_10_io_out_id_0) ^ ((fiEnable && (1974 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_678_0 <=( _mesh_5_10_io_out_id_0) ^ ((fiEnable && (1975 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_679_0 <=( _mesh_6_10_io_out_id_0) ^ ((fiEnable && (1976 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_680_0 <=( _mesh_7_10_io_out_id_0) ^ ((fiEnable && (1977 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_681_0 <=( _mesh_8_10_io_out_id_0) ^ ((fiEnable && (1978 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_682_0 <=( _mesh_9_10_io_out_id_0) ^ ((fiEnable && (1979 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_683_0 <=( _mesh_10_10_io_out_id_0) ^ ((fiEnable && (1980 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_684_0 <=( _mesh_11_10_io_out_id_0) ^ ((fiEnable && (1981 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_685_0 <=( _mesh_12_10_io_out_id_0) ^ ((fiEnable && (1982 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_686_0 <=( _mesh_13_10_io_out_id_0) ^ ((fiEnable && (1983 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_687_0 <=( _mesh_14_10_io_out_id_0) ^ ((fiEnable && (1984 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_688_0 <=( io_in_id_11_0) ^ ((fiEnable && (1985 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_689_0 <=( _mesh_0_11_io_out_id_0) ^ ((fiEnable && (1986 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_690_0 <=( _mesh_1_11_io_out_id_0) ^ ((fiEnable && (1987 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_691_0 <=( _mesh_2_11_io_out_id_0) ^ ((fiEnable && (1988 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_692_0 <=( _mesh_3_11_io_out_id_0) ^ ((fiEnable && (1989 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_693_0 <=( _mesh_4_11_io_out_id_0) ^ ((fiEnable && (1990 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_694_0 <=( _mesh_5_11_io_out_id_0) ^ ((fiEnable && (1991 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_695_0 <=( _mesh_6_11_io_out_id_0) ^ ((fiEnable && (1992 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_696_0 <=( _mesh_7_11_io_out_id_0) ^ ((fiEnable && (1993 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_697_0 <=( _mesh_8_11_io_out_id_0) ^ ((fiEnable && (1994 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_698_0 <=( _mesh_9_11_io_out_id_0) ^ ((fiEnable && (1995 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_699_0 <=( _mesh_10_11_io_out_id_0) ^ ((fiEnable && (1996 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_700_0 <=( _mesh_11_11_io_out_id_0) ^ ((fiEnable && (1997 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_701_0 <=( _mesh_12_11_io_out_id_0) ^ ((fiEnable && (1998 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_702_0 <=( _mesh_13_11_io_out_id_0) ^ ((fiEnable && (1999 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_703_0 <=( _mesh_14_11_io_out_id_0) ^ ((fiEnable && (2000 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_704_0 <=( io_in_id_12_0) ^ ((fiEnable && (2001 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_705_0 <=( _mesh_0_12_io_out_id_0) ^ ((fiEnable && (2002 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_706_0 <=( _mesh_1_12_io_out_id_0) ^ ((fiEnable && (2003 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_707_0 <=( _mesh_2_12_io_out_id_0) ^ ((fiEnable && (2004 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_708_0 <=( _mesh_3_12_io_out_id_0) ^ ((fiEnable && (2005 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_709_0 <=( _mesh_4_12_io_out_id_0) ^ ((fiEnable && (2006 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_710_0 <=( _mesh_5_12_io_out_id_0) ^ ((fiEnable && (2007 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_711_0 <=( _mesh_6_12_io_out_id_0) ^ ((fiEnable && (2008 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_712_0 <=( _mesh_7_12_io_out_id_0) ^ ((fiEnable && (2009 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_713_0 <=( _mesh_8_12_io_out_id_0) ^ ((fiEnable && (2010 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_714_0 <=( _mesh_9_12_io_out_id_0) ^ ((fiEnable && (2011 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_715_0 <=( _mesh_10_12_io_out_id_0) ^ ((fiEnable && (2012 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_716_0 <=( _mesh_11_12_io_out_id_0) ^ ((fiEnable && (2013 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_717_0 <=( _mesh_12_12_io_out_id_0) ^ ((fiEnable && (2014 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_718_0 <=( _mesh_13_12_io_out_id_0) ^ ((fiEnable && (2015 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_719_0 <=( _mesh_14_12_io_out_id_0) ^ ((fiEnable && (2016 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_720_0 <=( io_in_id_13_0) ^ ((fiEnable && (2017 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_721_0 <=( _mesh_0_13_io_out_id_0) ^ ((fiEnable && (2018 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_722_0 <=( _mesh_1_13_io_out_id_0) ^ ((fiEnable && (2019 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_723_0 <=( _mesh_2_13_io_out_id_0) ^ ((fiEnable && (2020 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_724_0 <=( _mesh_3_13_io_out_id_0) ^ ((fiEnable && (2021 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_725_0 <=( _mesh_4_13_io_out_id_0) ^ ((fiEnable && (2022 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_726_0 <=( _mesh_5_13_io_out_id_0) ^ ((fiEnable && (2023 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_727_0 <=( _mesh_6_13_io_out_id_0) ^ ((fiEnable && (2024 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_728_0 <=( _mesh_7_13_io_out_id_0) ^ ((fiEnable && (2025 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_729_0 <=( _mesh_8_13_io_out_id_0) ^ ((fiEnable && (2026 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_730_0 <=( _mesh_9_13_io_out_id_0) ^ ((fiEnable && (2027 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_731_0 <=( _mesh_10_13_io_out_id_0) ^ ((fiEnable && (2028 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_732_0 <=( _mesh_11_13_io_out_id_0) ^ ((fiEnable && (2029 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_733_0 <=( _mesh_12_13_io_out_id_0) ^ ((fiEnable && (2030 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_734_0 <=( _mesh_13_13_io_out_id_0) ^ ((fiEnable && (2031 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_735_0 <=( _mesh_14_13_io_out_id_0) ^ ((fiEnable && (2032 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_736_0 <=( io_in_id_14_0) ^ ((fiEnable && (2033 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_737_0 <=( _mesh_0_14_io_out_id_0) ^ ((fiEnable && (2034 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_738_0 <=( _mesh_1_14_io_out_id_0) ^ ((fiEnable && (2035 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_739_0 <=( _mesh_2_14_io_out_id_0) ^ ((fiEnable && (2036 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_740_0 <=( _mesh_3_14_io_out_id_0) ^ ((fiEnable && (2037 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_741_0 <=( _mesh_4_14_io_out_id_0) ^ ((fiEnable && (2038 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_742_0 <=( _mesh_5_14_io_out_id_0) ^ ((fiEnable && (2039 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_743_0 <=( _mesh_6_14_io_out_id_0) ^ ((fiEnable && (2040 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_744_0 <=( _mesh_7_14_io_out_id_0) ^ ((fiEnable && (2041 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_745_0 <=( _mesh_8_14_io_out_id_0) ^ ((fiEnable && (2042 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_746_0 <=( _mesh_9_14_io_out_id_0) ^ ((fiEnable && (2043 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_747_0 <=( _mesh_10_14_io_out_id_0) ^ ((fiEnable && (2044 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_748_0 <=( _mesh_11_14_io_out_id_0) ^ ((fiEnable && (2045 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_749_0 <=( _mesh_12_14_io_out_id_0) ^ ((fiEnable && (2046 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_750_0 <=( _mesh_13_14_io_out_id_0) ^ ((fiEnable && (2047 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_751_0 <=( _mesh_14_14_io_out_id_0) ^ ((fiEnable && (2048 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_752_0 <=( io_in_id_15_0) ^ ((fiEnable && (2049 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_753_0 <=( _mesh_0_15_io_out_id_0) ^ ((fiEnable && (2050 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_754_0 <=( _mesh_1_15_io_out_id_0) ^ ((fiEnable && (2051 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_755_0 <=( _mesh_2_15_io_out_id_0) ^ ((fiEnable && (2052 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_756_0 <=( _mesh_3_15_io_out_id_0) ^ ((fiEnable && (2053 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_757_0 <=( _mesh_4_15_io_out_id_0) ^ ((fiEnable && (2054 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_758_0 <=( _mesh_5_15_io_out_id_0) ^ ((fiEnable && (2055 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_759_0 <=( _mesh_6_15_io_out_id_0) ^ ((fiEnable && (2056 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_760_0 <=( _mesh_7_15_io_out_id_0) ^ ((fiEnable && (2057 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_761_0 <=( _mesh_8_15_io_out_id_0) ^ ((fiEnable && (2058 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_762_0 <=( _mesh_9_15_io_out_id_0) ^ ((fiEnable && (2059 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_763_0 <=( _mesh_10_15_io_out_id_0) ^ ((fiEnable && (2060 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_764_0 <=( _mesh_11_15_io_out_id_0) ^ ((fiEnable && (2061 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_765_0 <=( _mesh_12_15_io_out_id_0) ^ ((fiEnable && (2062 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_766_0 <=( _mesh_13_15_io_out_id_0) ^ ((fiEnable && (2063 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_767_0 <=( _mesh_14_15_io_out_id_0) ^ ((fiEnable && (2064 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_768_0 <=( io_in_last_0_0) ^ ((fiEnable && (2065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_769_0 <=( _mesh_0_0_io_out_last_0) ^ ((fiEnable && (2066 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_770_0 <=( _mesh_1_0_io_out_last_0) ^ ((fiEnable && (2067 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_771_0 <=( _mesh_2_0_io_out_last_0) ^ ((fiEnable && (2068 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_772_0 <=( _mesh_3_0_io_out_last_0) ^ ((fiEnable && (2069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_773_0 <=( _mesh_4_0_io_out_last_0) ^ ((fiEnable && (2070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_774_0 <=( _mesh_5_0_io_out_last_0) ^ ((fiEnable && (2071 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_775_0 <=( _mesh_6_0_io_out_last_0) ^ ((fiEnable && (2072 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_776_0 <=( _mesh_7_0_io_out_last_0) ^ ((fiEnable && (2073 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_777_0 <=( _mesh_8_0_io_out_last_0) ^ ((fiEnable && (2074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_778_0 <=( _mesh_9_0_io_out_last_0) ^ ((fiEnable && (2075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_779_0 <=( _mesh_10_0_io_out_last_0) ^ ((fiEnable && (2076 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_780_0 <=( _mesh_11_0_io_out_last_0) ^ ((fiEnable && (2077 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_781_0 <=( _mesh_12_0_io_out_last_0) ^ ((fiEnable && (2078 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_782_0 <=( _mesh_13_0_io_out_last_0) ^ ((fiEnable && (2079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_783_0 <=( _mesh_14_0_io_out_last_0) ^ ((fiEnable && (2080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_784_0 <=( io_in_last_1_0) ^ ((fiEnable && (2081 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_785_0 <=( _mesh_0_1_io_out_last_0) ^ ((fiEnable && (2082 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_786_0 <=( _mesh_1_1_io_out_last_0) ^ ((fiEnable && (2083 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_787_0 <=( _mesh_2_1_io_out_last_0) ^ ((fiEnable && (2084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_788_0 <=( _mesh_3_1_io_out_last_0) ^ ((fiEnable && (2085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_789_0 <=( _mesh_4_1_io_out_last_0) ^ ((fiEnable && (2086 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_790_0 <=( _mesh_5_1_io_out_last_0) ^ ((fiEnable && (2087 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_791_0 <=( _mesh_6_1_io_out_last_0) ^ ((fiEnable && (2088 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_792_0 <=( _mesh_7_1_io_out_last_0) ^ ((fiEnable && (2089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_793_0 <=( _mesh_8_1_io_out_last_0) ^ ((fiEnable && (2090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_794_0 <=( _mesh_9_1_io_out_last_0) ^ ((fiEnable && (2091 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_795_0 <=( _mesh_10_1_io_out_last_0) ^ ((fiEnable && (2092 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_796_0 <=( _mesh_11_1_io_out_last_0) ^ ((fiEnable && (2093 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_797_0 <=( _mesh_12_1_io_out_last_0) ^ ((fiEnable && (2094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_798_0 <=( _mesh_13_1_io_out_last_0) ^ ((fiEnable && (2095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_799_0 <=( _mesh_14_1_io_out_last_0) ^ ((fiEnable && (2096 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_800_0 <=( io_in_last_2_0) ^ ((fiEnable && (2097 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_801_0 <=( _mesh_0_2_io_out_last_0) ^ ((fiEnable && (2098 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_802_0 <=( _mesh_1_2_io_out_last_0) ^ ((fiEnable && (2099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_803_0 <=( _mesh_2_2_io_out_last_0) ^ ((fiEnable && (2100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_804_0 <=( _mesh_3_2_io_out_last_0) ^ ((fiEnable && (2101 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_805_0 <=( _mesh_4_2_io_out_last_0) ^ ((fiEnable && (2102 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_806_0 <=( _mesh_5_2_io_out_last_0) ^ ((fiEnable && (2103 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_807_0 <=( _mesh_6_2_io_out_last_0) ^ ((fiEnable && (2104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_808_0 <=( _mesh_7_2_io_out_last_0) ^ ((fiEnable && (2105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_809_0 <=( _mesh_8_2_io_out_last_0) ^ ((fiEnable && (2106 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_810_0 <=( _mesh_9_2_io_out_last_0) ^ ((fiEnable && (2107 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_811_0 <=( _mesh_10_2_io_out_last_0) ^ ((fiEnable && (2108 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_812_0 <=( _mesh_11_2_io_out_last_0) ^ ((fiEnable && (2109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_813_0 <=( _mesh_12_2_io_out_last_0) ^ ((fiEnable && (2110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_814_0 <=( _mesh_13_2_io_out_last_0) ^ ((fiEnable && (2111 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_815_0 <=( _mesh_14_2_io_out_last_0) ^ ((fiEnable && (2112 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_816_0 <=( io_in_last_3_0) ^ ((fiEnable && (2113 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_817_0 <=( _mesh_0_3_io_out_last_0) ^ ((fiEnable && (2114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_818_0 <=( _mesh_1_3_io_out_last_0) ^ ((fiEnable && (2115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_819_0 <=( _mesh_2_3_io_out_last_0) ^ ((fiEnable && (2116 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_820_0 <=( _mesh_3_3_io_out_last_0) ^ ((fiEnable && (2117 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_821_0 <=( _mesh_4_3_io_out_last_0) ^ ((fiEnable && (2118 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_822_0 <=( _mesh_5_3_io_out_last_0) ^ ((fiEnable && (2119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_823_0 <=( _mesh_6_3_io_out_last_0) ^ ((fiEnable && (2120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_824_0 <=( _mesh_7_3_io_out_last_0) ^ ((fiEnable && (2121 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_825_0 <=( _mesh_8_3_io_out_last_0) ^ ((fiEnable && (2122 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_826_0 <=( _mesh_9_3_io_out_last_0) ^ ((fiEnable && (2123 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_827_0 <=( _mesh_10_3_io_out_last_0) ^ ((fiEnable && (2124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_828_0 <=( _mesh_11_3_io_out_last_0) ^ ((fiEnable && (2125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_829_0 <=( _mesh_12_3_io_out_last_0) ^ ((fiEnable && (2126 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_830_0 <=( _mesh_13_3_io_out_last_0) ^ ((fiEnable && (2127 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_831_0 <=( _mesh_14_3_io_out_last_0) ^ ((fiEnable && (2128 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_832_0 <=( io_in_last_4_0) ^ ((fiEnable && (2129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_833_0 <=( _mesh_0_4_io_out_last_0) ^ ((fiEnable && (2130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_834_0 <=( _mesh_1_4_io_out_last_0) ^ ((fiEnable && (2131 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_835_0 <=( _mesh_2_4_io_out_last_0) ^ ((fiEnable && (2132 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_836_0 <=( _mesh_3_4_io_out_last_0) ^ ((fiEnable && (2133 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_837_0 <=( _mesh_4_4_io_out_last_0) ^ ((fiEnable && (2134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_838_0 <=( _mesh_5_4_io_out_last_0) ^ ((fiEnable && (2135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_839_0 <=( _mesh_6_4_io_out_last_0) ^ ((fiEnable && (2136 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_840_0 <=( _mesh_7_4_io_out_last_0) ^ ((fiEnable && (2137 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_841_0 <=( _mesh_8_4_io_out_last_0) ^ ((fiEnable && (2138 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_842_0 <=( _mesh_9_4_io_out_last_0) ^ ((fiEnable && (2139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_843_0 <=( _mesh_10_4_io_out_last_0) ^ ((fiEnable && (2140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_844_0 <=( _mesh_11_4_io_out_last_0) ^ ((fiEnable && (2141 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_845_0 <=( _mesh_12_4_io_out_last_0) ^ ((fiEnable && (2142 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_846_0 <=( _mesh_13_4_io_out_last_0) ^ ((fiEnable && (2143 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_847_0 <=( _mesh_14_4_io_out_last_0) ^ ((fiEnable && (2144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_848_0 <=( io_in_last_5_0) ^ ((fiEnable && (2145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_849_0 <=( _mesh_0_5_io_out_last_0) ^ ((fiEnable && (2146 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_850_0 <=( _mesh_1_5_io_out_last_0) ^ ((fiEnable && (2147 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_851_0 <=( _mesh_2_5_io_out_last_0) ^ ((fiEnable && (2148 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_852_0 <=( _mesh_3_5_io_out_last_0) ^ ((fiEnable && (2149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_853_0 <=( _mesh_4_5_io_out_last_0) ^ ((fiEnable && (2150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_854_0 <=( _mesh_5_5_io_out_last_0) ^ ((fiEnable && (2151 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_855_0 <=( _mesh_6_5_io_out_last_0) ^ ((fiEnable && (2152 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_856_0 <=( _mesh_7_5_io_out_last_0) ^ ((fiEnable && (2153 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_857_0 <=( _mesh_8_5_io_out_last_0) ^ ((fiEnable && (2154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_858_0 <=( _mesh_9_5_io_out_last_0) ^ ((fiEnable && (2155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_859_0 <=( _mesh_10_5_io_out_last_0) ^ ((fiEnable && (2156 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_860_0 <=( _mesh_11_5_io_out_last_0) ^ ((fiEnable && (2157 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_861_0 <=( _mesh_12_5_io_out_last_0) ^ ((fiEnable && (2158 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_862_0 <=( _mesh_13_5_io_out_last_0) ^ ((fiEnable && (2159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_863_0 <=( _mesh_14_5_io_out_last_0) ^ ((fiEnable && (2160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_864_0 <=( io_in_last_6_0) ^ ((fiEnable && (2161 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_865_0 <=( _mesh_0_6_io_out_last_0) ^ ((fiEnable && (2162 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_866_0 <=( _mesh_1_6_io_out_last_0) ^ ((fiEnable && (2163 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_867_0 <=( _mesh_2_6_io_out_last_0) ^ ((fiEnable && (2164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_868_0 <=( _mesh_3_6_io_out_last_0) ^ ((fiEnable && (2165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_869_0 <=( _mesh_4_6_io_out_last_0) ^ ((fiEnable && (2166 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_870_0 <=( _mesh_5_6_io_out_last_0) ^ ((fiEnable && (2167 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_871_0 <=( _mesh_6_6_io_out_last_0) ^ ((fiEnable && (2168 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_872_0 <=( _mesh_7_6_io_out_last_0) ^ ((fiEnable && (2169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_873_0 <=( _mesh_8_6_io_out_last_0) ^ ((fiEnable && (2170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_874_0 <=( _mesh_9_6_io_out_last_0) ^ ((fiEnable && (2171 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_875_0 <=( _mesh_10_6_io_out_last_0) ^ ((fiEnable && (2172 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_876_0 <=( _mesh_11_6_io_out_last_0) ^ ((fiEnable && (2173 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_877_0 <=( _mesh_12_6_io_out_last_0) ^ ((fiEnable && (2174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_878_0 <=( _mesh_13_6_io_out_last_0) ^ ((fiEnable && (2175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_879_0 <=( _mesh_14_6_io_out_last_0) ^ ((fiEnable && (2176 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_880_0 <=( io_in_last_7_0) ^ ((fiEnable && (2177 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_881_0 <=( _mesh_0_7_io_out_last_0) ^ ((fiEnable && (2178 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_882_0 <=( _mesh_1_7_io_out_last_0) ^ ((fiEnable && (2179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_883_0 <=( _mesh_2_7_io_out_last_0) ^ ((fiEnable && (2180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_884_0 <=( _mesh_3_7_io_out_last_0) ^ ((fiEnable && (2181 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_885_0 <=( _mesh_4_7_io_out_last_0) ^ ((fiEnable && (2182 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_886_0 <=( _mesh_5_7_io_out_last_0) ^ ((fiEnable && (2183 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_887_0 <=( _mesh_6_7_io_out_last_0) ^ ((fiEnable && (2184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_888_0 <=( _mesh_7_7_io_out_last_0) ^ ((fiEnable && (2185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_889_0 <=( _mesh_8_7_io_out_last_0) ^ ((fiEnable && (2186 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_890_0 <=( _mesh_9_7_io_out_last_0) ^ ((fiEnable && (2187 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_891_0 <=( _mesh_10_7_io_out_last_0) ^ ((fiEnable && (2188 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_892_0 <=( _mesh_11_7_io_out_last_0) ^ ((fiEnable && (2189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_893_0 <=( _mesh_12_7_io_out_last_0) ^ ((fiEnable && (2190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_894_0 <=( _mesh_13_7_io_out_last_0) ^ ((fiEnable && (2191 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_895_0 <=( _mesh_14_7_io_out_last_0) ^ ((fiEnable && (2192 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_896_0 <=( io_in_last_8_0) ^ ((fiEnable && (2193 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_897_0 <=( _mesh_0_8_io_out_last_0) ^ ((fiEnable && (2194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_898_0 <=( _mesh_1_8_io_out_last_0) ^ ((fiEnable && (2195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_899_0 <=( _mesh_2_8_io_out_last_0) ^ ((fiEnable && (2196 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_900_0 <=( _mesh_3_8_io_out_last_0) ^ ((fiEnable && (2197 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_901_0 <=( _mesh_4_8_io_out_last_0) ^ ((fiEnable && (2198 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_902_0 <=( _mesh_5_8_io_out_last_0) ^ ((fiEnable && (2199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_903_0 <=( _mesh_6_8_io_out_last_0) ^ ((fiEnable && (2200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_904_0 <=( _mesh_7_8_io_out_last_0) ^ ((fiEnable && (2201 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_905_0 <=( _mesh_8_8_io_out_last_0) ^ ((fiEnable && (2202 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_906_0 <=( _mesh_9_8_io_out_last_0) ^ ((fiEnable && (2203 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_907_0 <=( _mesh_10_8_io_out_last_0) ^ ((fiEnable && (2204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_908_0 <=( _mesh_11_8_io_out_last_0) ^ ((fiEnable && (2205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_909_0 <=( _mesh_12_8_io_out_last_0) ^ ((fiEnable && (2206 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_910_0 <=( _mesh_13_8_io_out_last_0) ^ ((fiEnable && (2207 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_911_0 <=( _mesh_14_8_io_out_last_0) ^ ((fiEnable && (2208 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_912_0 <=( io_in_last_9_0) ^ ((fiEnable && (2209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_913_0 <=( _mesh_0_9_io_out_last_0) ^ ((fiEnable && (2210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_914_0 <=( _mesh_1_9_io_out_last_0) ^ ((fiEnable && (2211 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_915_0 <=( _mesh_2_9_io_out_last_0) ^ ((fiEnable && (2212 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_916_0 <=( _mesh_3_9_io_out_last_0) ^ ((fiEnable && (2213 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_917_0 <=( _mesh_4_9_io_out_last_0) ^ ((fiEnable && (2214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_918_0 <=( _mesh_5_9_io_out_last_0) ^ ((fiEnable && (2215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_919_0 <=( _mesh_6_9_io_out_last_0) ^ ((fiEnable && (2216 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_920_0 <=( _mesh_7_9_io_out_last_0) ^ ((fiEnable && (2217 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_921_0 <=( _mesh_8_9_io_out_last_0) ^ ((fiEnable && (2218 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_922_0 <=( _mesh_9_9_io_out_last_0) ^ ((fiEnable && (2219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_923_0 <=( _mesh_10_9_io_out_last_0) ^ ((fiEnable && (2220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_924_0 <=( _mesh_11_9_io_out_last_0) ^ ((fiEnable && (2221 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_925_0 <=( _mesh_12_9_io_out_last_0) ^ ((fiEnable && (2222 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_926_0 <=( _mesh_13_9_io_out_last_0) ^ ((fiEnable && (2223 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_927_0 <=( _mesh_14_9_io_out_last_0) ^ ((fiEnable && (2224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_928_0 <=( io_in_last_10_0) ^ ((fiEnable && (2225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_929_0 <=( _mesh_0_10_io_out_last_0) ^ ((fiEnable && (2226 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_930_0 <=( _mesh_1_10_io_out_last_0) ^ ((fiEnable && (2227 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_931_0 <=( _mesh_2_10_io_out_last_0) ^ ((fiEnable && (2228 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_932_0 <=( _mesh_3_10_io_out_last_0) ^ ((fiEnable && (2229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_933_0 <=( _mesh_4_10_io_out_last_0) ^ ((fiEnable && (2230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_934_0 <=( _mesh_5_10_io_out_last_0) ^ ((fiEnable && (2231 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_935_0 <=( _mesh_6_10_io_out_last_0) ^ ((fiEnable && (2232 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_936_0 <=( _mesh_7_10_io_out_last_0) ^ ((fiEnable && (2233 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_937_0 <=( _mesh_8_10_io_out_last_0) ^ ((fiEnable && (2234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_938_0 <=( _mesh_9_10_io_out_last_0) ^ ((fiEnable && (2235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_939_0 <=( _mesh_10_10_io_out_last_0) ^ ((fiEnable && (2236 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_940_0 <=( _mesh_11_10_io_out_last_0) ^ ((fiEnable && (2237 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_941_0 <=( _mesh_12_10_io_out_last_0) ^ ((fiEnable && (2238 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_942_0 <=( _mesh_13_10_io_out_last_0) ^ ((fiEnable && (2239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_943_0 <=( _mesh_14_10_io_out_last_0) ^ ((fiEnable && (2240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_944_0 <=( io_in_last_11_0) ^ ((fiEnable && (2241 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_945_0 <=( _mesh_0_11_io_out_last_0) ^ ((fiEnable && (2242 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_946_0 <=( _mesh_1_11_io_out_last_0) ^ ((fiEnable && (2243 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_947_0 <=( _mesh_2_11_io_out_last_0) ^ ((fiEnable && (2244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_948_0 <=( _mesh_3_11_io_out_last_0) ^ ((fiEnable && (2245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_949_0 <=( _mesh_4_11_io_out_last_0) ^ ((fiEnable && (2246 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_950_0 <=( _mesh_5_11_io_out_last_0) ^ ((fiEnable && (2247 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_951_0 <=( _mesh_6_11_io_out_last_0) ^ ((fiEnable && (2248 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_952_0 <=( _mesh_7_11_io_out_last_0) ^ ((fiEnable && (2249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_953_0 <=( _mesh_8_11_io_out_last_0) ^ ((fiEnable && (2250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_954_0 <=( _mesh_9_11_io_out_last_0) ^ ((fiEnable && (2251 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_955_0 <=( _mesh_10_11_io_out_last_0) ^ ((fiEnable && (2252 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_956_0 <=( _mesh_11_11_io_out_last_0) ^ ((fiEnable && (2253 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_957_0 <=( _mesh_12_11_io_out_last_0) ^ ((fiEnable && (2254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_958_0 <=( _mesh_13_11_io_out_last_0) ^ ((fiEnable && (2255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_959_0 <=( _mesh_14_11_io_out_last_0) ^ ((fiEnable && (2256 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_960_0 <=( io_in_last_12_0) ^ ((fiEnable && (2257 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_961_0 <=( _mesh_0_12_io_out_last_0) ^ ((fiEnable && (2258 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_962_0 <=( _mesh_1_12_io_out_last_0) ^ ((fiEnable && (2259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_963_0 <=( _mesh_2_12_io_out_last_0) ^ ((fiEnable && (2260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_964_0 <=( _mesh_3_12_io_out_last_0) ^ ((fiEnable && (2261 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_965_0 <=( _mesh_4_12_io_out_last_0) ^ ((fiEnable && (2262 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_966_0 <=( _mesh_5_12_io_out_last_0) ^ ((fiEnable && (2263 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_967_0 <=( _mesh_6_12_io_out_last_0) ^ ((fiEnable && (2264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_968_0 <=( _mesh_7_12_io_out_last_0) ^ ((fiEnable && (2265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_969_0 <=( _mesh_8_12_io_out_last_0) ^ ((fiEnable && (2266 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_970_0 <=( _mesh_9_12_io_out_last_0) ^ ((fiEnable && (2267 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_971_0 <=( _mesh_10_12_io_out_last_0) ^ ((fiEnable && (2268 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_972_0 <=( _mesh_11_12_io_out_last_0) ^ ((fiEnable && (2269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_973_0 <=( _mesh_12_12_io_out_last_0) ^ ((fiEnable && (2270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_974_0 <=( _mesh_13_12_io_out_last_0) ^ ((fiEnable && (2271 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_975_0 <=( _mesh_14_12_io_out_last_0) ^ ((fiEnable && (2272 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_976_0 <=( io_in_last_13_0) ^ ((fiEnable && (2273 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_977_0 <=( _mesh_0_13_io_out_last_0) ^ ((fiEnable && (2274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_978_0 <=( _mesh_1_13_io_out_last_0) ^ ((fiEnable && (2275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_979_0 <=( _mesh_2_13_io_out_last_0) ^ ((fiEnable && (2276 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_980_0 <=( _mesh_3_13_io_out_last_0) ^ ((fiEnable && (2277 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_981_0 <=( _mesh_4_13_io_out_last_0) ^ ((fiEnable && (2278 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_982_0 <=( _mesh_5_13_io_out_last_0) ^ ((fiEnable && (2279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_983_0 <=( _mesh_6_13_io_out_last_0) ^ ((fiEnable && (2280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_984_0 <=( _mesh_7_13_io_out_last_0) ^ ((fiEnable && (2281 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_985_0 <=( _mesh_8_13_io_out_last_0) ^ ((fiEnable && (2282 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_986_0 <=( _mesh_9_13_io_out_last_0) ^ ((fiEnable && (2283 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_987_0 <=( _mesh_10_13_io_out_last_0) ^ ((fiEnable && (2284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_988_0 <=( _mesh_11_13_io_out_last_0) ^ ((fiEnable && (2285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_989_0 <=( _mesh_12_13_io_out_last_0) ^ ((fiEnable && (2286 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_990_0 <=( _mesh_13_13_io_out_last_0) ^ ((fiEnable && (2287 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_991_0 <=( _mesh_14_13_io_out_last_0) ^ ((fiEnable && (2288 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_992_0 <=( io_in_last_14_0) ^ ((fiEnable && (2289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_993_0 <=( _mesh_0_14_io_out_last_0) ^ ((fiEnable && (2290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_994_0 <=( _mesh_1_14_io_out_last_0) ^ ((fiEnable && (2291 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_995_0 <=( _mesh_2_14_io_out_last_0) ^ ((fiEnable && (2292 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_996_0 <=( _mesh_3_14_io_out_last_0) ^ ((fiEnable && (2293 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_997_0 <=( _mesh_4_14_io_out_last_0) ^ ((fiEnable && (2294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_998_0 <=( _mesh_5_14_io_out_last_0) ^ ((fiEnable && (2295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_999_0 <=( _mesh_6_14_io_out_last_0) ^ ((fiEnable && (2296 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1000_0 <=( _mesh_7_14_io_out_last_0) ^ ((fiEnable && (2297 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1001_0 <=( _mesh_8_14_io_out_last_0) ^ ((fiEnable && (2298 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1002_0 <=( _mesh_9_14_io_out_last_0) ^ ((fiEnable && (2299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1003_0 <=( _mesh_10_14_io_out_last_0) ^ ((fiEnable && (2300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1004_0 <=( _mesh_11_14_io_out_last_0) ^ ((fiEnable && (2301 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1005_0 <=( _mesh_12_14_io_out_last_0) ^ ((fiEnable && (2302 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1006_0 <=( _mesh_13_14_io_out_last_0) ^ ((fiEnable && (2303 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1007_0 <=( _mesh_14_14_io_out_last_0) ^ ((fiEnable && (2304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1008_0 <=( io_in_last_15_0) ^ ((fiEnable && (2305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1009_0 <=( _mesh_0_15_io_out_last_0) ^ ((fiEnable && (2306 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1010_0 <=( _mesh_1_15_io_out_last_0) ^ ((fiEnable && (2307 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1011_0 <=( _mesh_2_15_io_out_last_0) ^ ((fiEnable && (2308 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1012_0 <=( _mesh_3_15_io_out_last_0) ^ ((fiEnable && (2309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1013_0 <=( _mesh_4_15_io_out_last_0) ^ ((fiEnable && (2310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1014_0 <=( _mesh_5_15_io_out_last_0) ^ ((fiEnable && (2311 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1015_0 <=( _mesh_6_15_io_out_last_0) ^ ((fiEnable && (2312 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1016_0 <=( _mesh_7_15_io_out_last_0) ^ ((fiEnable && (2313 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1017_0 <=( _mesh_8_15_io_out_last_0) ^ ((fiEnable && (2314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1018_0 <=( _mesh_9_15_io_out_last_0) ^ ((fiEnable && (2315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1019_0 <=( _mesh_10_15_io_out_last_0) ^ ((fiEnable && (2316 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1020_0 <=( _mesh_11_15_io_out_last_0) ^ ((fiEnable && (2317 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1021_0 <=( _mesh_12_15_io_out_last_0) ^ ((fiEnable && (2318 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1022_0 <=( _mesh_13_15_io_out_last_0) ^ ((fiEnable && (2319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1023_0 <=( _mesh_14_15_io_out_last_0) ^ ((fiEnable && (2320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1024_0 <=( _mesh_15_0_io_out_b_0) ^ ((fiEnable && (2321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1025_0 <=( _mesh_15_0_io_out_c_0) ^ ((fiEnable && (2322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1026_0 <=( _mesh_15_0_io_out_valid_0) ^ ((fiEnable && (2323 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1027_0_dataflow <=( _mesh_15_0_io_out_control_0_dataflow) ^ ((fiEnable && (2324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1028_0 <=( _mesh_15_0_io_out_id_0) ^ ((fiEnable && (2325 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_1029_0 <=( _mesh_15_0_io_out_last_0) ^ ((fiEnable && (2326 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1030_0 <=( _mesh_15_1_io_out_b_0) ^ ((fiEnable && (2327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1031_0 <=( _mesh_15_1_io_out_c_0) ^ ((fiEnable && (2328 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1036_0 <=( _mesh_15_2_io_out_b_0) ^ ((fiEnable && (2329 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1037_0 <=( _mesh_15_2_io_out_c_0) ^ ((fiEnable && (2330 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1042_0 <=( _mesh_15_3_io_out_b_0) ^ ((fiEnable && (2331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1043_0 <=( _mesh_15_3_io_out_c_0) ^ ((fiEnable && (2332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1048_0 <=( _mesh_15_4_io_out_b_0) ^ ((fiEnable && (2333 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1049_0 <=( _mesh_15_4_io_out_c_0) ^ ((fiEnable && (2334 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1054_0 <=( _mesh_15_5_io_out_b_0) ^ ((fiEnable && (2335 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1055_0 <=( _mesh_15_5_io_out_c_0) ^ ((fiEnable && (2336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1060_0 <=( _mesh_15_6_io_out_b_0) ^ ((fiEnable && (2337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1061_0 <=( _mesh_15_6_io_out_c_0) ^ ((fiEnable && (2338 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1066_0 <=( _mesh_15_7_io_out_b_0) ^ ((fiEnable && (2339 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1067_0 <=( _mesh_15_7_io_out_c_0) ^ ((fiEnable && (2340 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1072_0 <=( _mesh_15_8_io_out_b_0) ^ ((fiEnable && (2341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1073_0 <=( _mesh_15_8_io_out_c_0) ^ ((fiEnable && (2342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1078_0 <=( _mesh_15_9_io_out_b_0) ^ ((fiEnable && (2343 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1079_0 <=( _mesh_15_9_io_out_c_0) ^ ((fiEnable && (2344 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1084_0 <=( _mesh_15_10_io_out_b_0) ^ ((fiEnable && (2345 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1085_0 <=( _mesh_15_10_io_out_c_0) ^ ((fiEnable && (2346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1090_0 <=( _mesh_15_11_io_out_b_0) ^ ((fiEnable && (2347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1091_0 <=( _mesh_15_11_io_out_c_0) ^ ((fiEnable && (2348 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1096_0 <=( _mesh_15_12_io_out_b_0) ^ ((fiEnable && (2349 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1097_0 <=( _mesh_15_12_io_out_c_0) ^ ((fiEnable && (2350 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1102_0 <=( _mesh_15_13_io_out_b_0) ^ ((fiEnable && (2351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1103_0 <=( _mesh_15_13_io_out_c_0) ^ ((fiEnable && (2352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1108_0 <=( _mesh_15_14_io_out_b_0) ^ ((fiEnable && (2353 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1109_0 <=( _mesh_15_14_io_out_c_0) ^ ((fiEnable && (2354 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1114_0 <=( _mesh_15_15_io_out_b_0) ^ ((fiEnable && (2355 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1115_0 <=( _mesh_15_15_io_out_c_0) ^ ((fiEnable && (2356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	logic [31:0] _RANDOM_3;
	logic [31:0] _RANDOM_4;
	logic [31:0] _RANDOM_5;
	logic [31:0] _RANDOM_6;
	logic [31:0] _RANDOM_7;
	logic [31:0] _RANDOM_8;
	logic [31:0] _RANDOM_9;
	logic [31:0] _RANDOM_10;
	logic [31:0] _RANDOM_11;
	logic [31:0] _RANDOM_12;
	logic [31:0] _RANDOM_13;
	logic [31:0] _RANDOM_14;
	logic [31:0] _RANDOM_15;
	logic [31:0] _RANDOM_16;
	logic [31:0] _RANDOM_17;
	logic [31:0] _RANDOM_18;
	logic [31:0] _RANDOM_19;
	logic [31:0] _RANDOM_20;
	logic [31:0] _RANDOM_21;
	logic [31:0] _RANDOM_22;
	logic [31:0] _RANDOM_23;
	logic [31:0] _RANDOM_24;
	logic [31:0] _RANDOM_25;
	logic [31:0] _RANDOM_26;
	logic [31:0] _RANDOM_27;
	logic [31:0] _RANDOM_28;
	logic [31:0] _RANDOM_29;
	logic [31:0] _RANDOM_30;
	logic [31:0] _RANDOM_31;
	logic [31:0] _RANDOM_32;
	logic [31:0] _RANDOM_33;
	logic [31:0] _RANDOM_34;
	logic [31:0] _RANDOM_35;
	logic [31:0] _RANDOM_36;
	logic [31:0] _RANDOM_37;
	logic [31:0] _RANDOM_38;
	logic [31:0] _RANDOM_39;
	logic [31:0] _RANDOM_40;
	logic [31:0] _RANDOM_41;
	logic [31:0] _RANDOM_42;
	logic [31:0] _RANDOM_43;
	logic [31:0] _RANDOM_44;
	logic [31:0] _RANDOM_45;
	logic [31:0] _RANDOM_46;
	logic [31:0] _RANDOM_47;
	logic [31:0] _RANDOM_48;
	logic [31:0] _RANDOM_49;
	logic [31:0] _RANDOM_50;
	logic [31:0] _RANDOM_51;
	logic [31:0] _RANDOM_52;
	logic [31:0] _RANDOM_53;
	logic [31:0] _RANDOM_54;
	logic [31:0] _RANDOM_55;
	logic [31:0] _RANDOM_56;
	logic [31:0] _RANDOM_57;
	logic [31:0] _RANDOM_58;
	logic [31:0] _RANDOM_59;
	logic [31:0] _RANDOM_60;
	logic [31:0] _RANDOM_61;
	logic [31:0] _RANDOM_62;
	logic [31:0] _RANDOM_63;
	logic [31:0] _RANDOM_64;
	logic [31:0] _RANDOM_65;
	logic [31:0] _RANDOM_66;
	logic [31:0] _RANDOM_67;
	logic [31:0] _RANDOM_68;
	logic [31:0] _RANDOM_69;
	logic [31:0] _RANDOM_70;
	logic [31:0] _RANDOM_71;
	logic [31:0] _RANDOM_72;
	logic [31:0] _RANDOM_73;
	logic [31:0] _RANDOM_74;
	logic [31:0] _RANDOM_75;
	logic [31:0] _RANDOM_76;
	logic [31:0] _RANDOM_77;
	logic [31:0] _RANDOM_78;
	logic [31:0] _RANDOM_79;
	logic [31:0] _RANDOM_80;
	logic [31:0] _RANDOM_81;
	logic [31:0] _RANDOM_82;
	logic [31:0] _RANDOM_83;
	logic [31:0] _RANDOM_84;
	logic [31:0] _RANDOM_85;
	logic [31:0] _RANDOM_86;
	logic [31:0] _RANDOM_87;
	logic [31:0] _RANDOM_88;
	logic [31:0] _RANDOM_89;
	logic [31:0] _RANDOM_90;
	logic [31:0] _RANDOM_91;
	logic [31:0] _RANDOM_92;
	logic [31:0] _RANDOM_93;
	logic [31:0] _RANDOM_94;
	logic [31:0] _RANDOM_95;
	logic [31:0] _RANDOM_96;
	logic [31:0] _RANDOM_97;
	logic [31:0] _RANDOM_98;
	logic [31:0] _RANDOM_99;
	logic [31:0] _RANDOM_100;
	logic [31:0] _RANDOM_101;
	logic [31:0] _RANDOM_102;
	logic [31:0] _RANDOM_103;
	logic [31:0] _RANDOM_104;
	logic [31:0] _RANDOM_105;
	logic [31:0] _RANDOM_106;
	logic [31:0] _RANDOM_107;
	logic [31:0] _RANDOM_108;
	logic [31:0] _RANDOM_109;
	logic [31:0] _RANDOM_110;
	logic [31:0] _RANDOM_111;
	logic [31:0] _RANDOM_112;
	logic [31:0] _RANDOM_113;
	logic [31:0] _RANDOM_114;
	logic [31:0] _RANDOM_115;
	logic [31:0] _RANDOM_116;
	logic [31:0] _RANDOM_117;
	logic [31:0] _RANDOM_118;
	logic [31:0] _RANDOM_119;
	logic [31:0] _RANDOM_120;
	logic [31:0] _RANDOM_121;
	logic [31:0] _RANDOM_122;
	logic [31:0] _RANDOM_123;
	logic [31:0] _RANDOM_124;
	logic [31:0] _RANDOM_125;
	logic [31:0] _RANDOM_126;
	logic [31:0] _RANDOM_127;
	logic [31:0] _RANDOM_128;
	logic [31:0] _RANDOM_129;
	logic [31:0] _RANDOM_130;
	logic [31:0] _RANDOM_131;
	logic [31:0] _RANDOM_132;
	logic [31:0] _RANDOM_133;
	logic [31:0] _RANDOM_134;
	logic [31:0] _RANDOM_135;
	logic [31:0] _RANDOM_136;
	logic [31:0] _RANDOM_137;
	logic [31:0] _RANDOM_138;
	logic [31:0] _RANDOM_139;
	logic [31:0] _RANDOM_140;
	logic [31:0] _RANDOM_141;
	logic [31:0] _RANDOM_142;
	logic [31:0] _RANDOM_143;
	logic [31:0] _RANDOM_144;
	logic [31:0] _RANDOM_145;
	logic [31:0] _RANDOM_146;
	logic [31:0] _RANDOM_147;
	logic [31:0] _RANDOM_148;
	logic [31:0] _RANDOM_149;
	logic [31:0] _RANDOM_150;
	logic [31:0] _RANDOM_151;
	logic [31:0] _RANDOM_152;
	logic [31:0] _RANDOM_153;
	logic [31:0] _RANDOM_154;
	logic [31:0] _RANDOM_155;
	logic [31:0] _RANDOM_156;
	logic [31:0] _RANDOM_157;
	logic [31:0] _RANDOM_158;
	logic [31:0] _RANDOM_159;
	logic [31:0] _RANDOM_160;
	logic [31:0] _RANDOM_161;
	logic [31:0] _RANDOM_162;
	logic [31:0] _RANDOM_163;
	logic [31:0] _RANDOM_164;
	logic [31:0] _RANDOM_165;
	logic [31:0] _RANDOM_166;
	logic [31:0] _RANDOM_167;
	logic [31:0] _RANDOM_168;
	logic [31:0] _RANDOM_169;
	logic [31:0] _RANDOM_170;
	logic [31:0] _RANDOM_171;
	logic [31:0] _RANDOM_172;
	logic [31:0] _RANDOM_173;
	logic [31:0] _RANDOM_174;
	logic [31:0] _RANDOM_175;
	logic [31:0] _RANDOM_176;
	logic [31:0] _RANDOM_177;
	logic [31:0] _RANDOM_178;
	logic [31:0] _RANDOM_179;
	logic [31:0] _RANDOM_180;
	logic [31:0] _RANDOM_181;
	logic [31:0] _RANDOM_182;
	logic [31:0] _RANDOM_183;
	logic [31:0] _RANDOM_184;
	logic [31:0] _RANDOM_185;
	logic [31:0] _RANDOM_186;
	logic [31:0] _RANDOM_187;
	logic [31:0] _RANDOM_188;
	logic [31:0] _RANDOM_189;
	logic [31:0] _RANDOM_190;
	logic [31:0] _RANDOM_191;
	logic [31:0] _RANDOM_192;
	logic [31:0] _RANDOM_193;
	logic [31:0] _RANDOM_194;
	logic [31:0] _RANDOM_195;
	logic [31:0] _RANDOM_196;
	logic [31:0] _RANDOM_197;
	logic [31:0] _RANDOM_198;
	logic [31:0] _RANDOM_199;
	logic [31:0] _RANDOM_200;
	logic [31:0] _RANDOM_201;
	logic [31:0] _RANDOM_202;
	logic [31:0] _RANDOM_203;
	logic [31:0] _RANDOM_204;
	logic [31:0] _RANDOM_205;
	logic [31:0] _RANDOM_206;
	logic [31:0] _RANDOM_207;
	logic [31:0] _RANDOM_208;
	logic [31:0] _RANDOM_209;
	logic [31:0] _RANDOM_210;
	logic [31:0] _RANDOM_211;
	logic [31:0] _RANDOM_212;
	logic [31:0] _RANDOM_213;
	logic [31:0] _RANDOM_214;
	logic [31:0] _RANDOM_215;
	logic [31:0] _RANDOM_216;
	logic [31:0] _RANDOM_217;
	logic [31:0] _RANDOM_218;
	logic [31:0] _RANDOM_219;
	logic [31:0] _RANDOM_220;
	logic [31:0] _RANDOM_221;
	logic [31:0] _RANDOM_222;
	logic [31:0] _RANDOM_223;
	logic [31:0] _RANDOM_224;
	logic [31:0] _RANDOM_225;
	logic [31:0] _RANDOM_226;
	logic [31:0] _RANDOM_227;
	logic [31:0] _RANDOM_228;
	logic [31:0] _RANDOM_229;
	logic [31:0] _RANDOM_230;
	logic [31:0] _RANDOM_231;
	logic [31:0] _RANDOM_232;
	logic [31:0] _RANDOM_233;
	logic [31:0] _RANDOM_234;
	logic [31:0] _RANDOM_235;
	logic [31:0] _RANDOM_236;
	logic [31:0] _RANDOM_237;
	logic [31:0] _RANDOM_238;
	logic [31:0] _RANDOM_239;
	logic [31:0] _RANDOM_240;
	logic [31:0] _RANDOM_241;
	logic [31:0] _RANDOM_242;
	logic [31:0] _RANDOM_243;
	logic [31:0] _RANDOM_244;
	logic [31:0] _RANDOM_245;
	logic [31:0] _RANDOM_246;
	logic [31:0] _RANDOM_247;
	logic [31:0] _RANDOM_248;
	logic [31:0] _RANDOM_249;
	logic [31:0] _RANDOM_250;
	logic [31:0] _RANDOM_251;
	logic [31:0] _RANDOM_252;
	logic [31:0] _RANDOM_253;
	logic [31:0] _RANDOM_254;
	logic [31:0] _RANDOM_255;
	logic [31:0] _RANDOM_256;
	logic [31:0] _RANDOM_257;
	logic [31:0] _RANDOM_258;
	logic [31:0] _RANDOM_259;
	logic [31:0] _RANDOM_260;
	logic [31:0] _RANDOM_261;
	logic [31:0] _RANDOM_262;
	logic [31:0] _RANDOM_263;
	logic [31:0] _RANDOM_264;
	logic [31:0] _RANDOM_265;
	logic [31:0] _RANDOM_266;
	logic [31:0] _RANDOM_267;
	logic [31:0] _RANDOM_268;
	logic [31:0] _RANDOM_269;
	logic [31:0] _RANDOM_270;
	logic [31:0] _RANDOM_271;
	logic [31:0] _RANDOM_272;
	logic [31:0] _RANDOM_273;
	logic [31:0] _RANDOM_274;
	logic [31:0] _RANDOM_275;
	logic [31:0] _RANDOM_276;
	logic [31:0] _RANDOM_277;
	logic [31:0] _RANDOM_278;
	logic [31:0] _RANDOM_279;
	logic [31:0] _RANDOM_280;
	logic [31:0] _RANDOM_281;
	logic [31:0] _RANDOM_282;
	logic [31:0] _RANDOM_283;
	logic [31:0] _RANDOM_284;
	logic [31:0] _RANDOM_285;
	logic [31:0] _RANDOM_286;
	logic [31:0] _RANDOM_287;
	logic [31:0] _RANDOM_288;
	logic [31:0] _RANDOM_289;
	logic [31:0] _RANDOM_290;
	logic [31:0] _RANDOM_291;
	logic [31:0] _RANDOM_292;
	logic [31:0] _RANDOM_293;
	logic [31:0] _RANDOM_294;
	logic [31:0] _RANDOM_295;
	logic [31:0] _RANDOM_296;
	logic [31:0] _RANDOM_297;
	logic [31:0] _RANDOM_298;
	logic [31:0] _RANDOM_299;
	logic [31:0] _RANDOM_300;
	logic [31:0] _RANDOM_301;
	logic [31:0] _RANDOM_302;
	logic [31:0] _RANDOM_303;
	logic [31:0] _RANDOM_304;
	logic [31:0] _RANDOM_305;
	logic [31:0] _RANDOM_306;
	logic [31:0] _RANDOM_307;
	logic [31:0] _RANDOM_308;
	logic [31:0] _RANDOM_309;
	logic [31:0] _RANDOM_310;
	logic [31:0] _RANDOM_311;
	logic [31:0] _RANDOM_312;
	logic [31:0] _RANDOM_313;
	logic [31:0] _RANDOM_314;
	logic [31:0] _RANDOM_315;
	logic [31:0] _RANDOM_316;
	logic [31:0] _RANDOM_317;
	logic [31:0] _RANDOM_318;
	logic [31:0] _RANDOM_319;
	logic [31:0] _RANDOM_320;
	logic [31:0] _RANDOM_321;
	logic [31:0] _RANDOM_322;
	logic [31:0] _RANDOM_323;
	logic [31:0] _RANDOM_324;
	logic [31:0] _RANDOM_325;
	logic [31:0] _RANDOM_326;
	logic [31:0] _RANDOM_327;
	logic [31:0] _RANDOM_328;
	logic [31:0] _RANDOM_329;
	logic [31:0] _RANDOM_330;
	logic [31:0] _RANDOM_331;
	logic [31:0] _RANDOM_332;
	logic [31:0] _RANDOM_333;
	logic [31:0] _RANDOM_334;
	logic [31:0] _RANDOM_335;
	logic [31:0] _RANDOM_336;
	logic [31:0] _RANDOM_337;
	logic [31:0] _RANDOM_338;
	logic [31:0] _RANDOM_339;
	logic [31:0] _RANDOM_340;
	logic [31:0] _RANDOM_341;
	logic [31:0] _RANDOM_342;
	logic [31:0] _RANDOM_343;
	logic [31:0] _RANDOM_344;
	logic [31:0] _RANDOM_345;
	logic [31:0] _RANDOM_346;
	logic [31:0] _RANDOM_347;
	logic [31:0] _RANDOM_348;
	logic [31:0] _RANDOM_349;
	logic [31:0] _RANDOM_350;
	logic [31:0] _RANDOM_351;
	logic [31:0] _RANDOM_352;
	logic [31:0] _RANDOM_353;
	logic [31:0] _RANDOM_354;
	logic [31:0] _RANDOM_355;
	logic [31:0] _RANDOM_356;
	logic [31:0] _RANDOM_357;
	logic [31:0] _RANDOM_358;
	logic [31:0] _RANDOM_359;
	logic [31:0] _RANDOM_360;
	logic [31:0] _RANDOM_361;
	logic [31:0] _RANDOM_362;
	logic [31:0] _RANDOM_363;
	logic [31:0] _RANDOM_364;
	logic [31:0] _RANDOM_365;
	logic [31:0] _RANDOM_366;
	logic [31:0] _RANDOM_367;
	logic [31:0] _RANDOM_368;
	logic [31:0] _RANDOM_369;
	logic [31:0] _RANDOM_370;
	logic [31:0] _RANDOM_371;
	logic [31:0] _RANDOM_372;
	logic [31:0] _RANDOM_373;
	logic [31:0] _RANDOM_374;
	logic [31:0] _RANDOM_375;
	logic [31:0] _RANDOM_376;
	logic [31:0] _RANDOM_377;
	logic [31:0] _RANDOM_378;
	logic [31:0] _RANDOM_379;
	logic [31:0] _RANDOM_380;
	logic [31:0] _RANDOM_381;
	logic [31:0] _RANDOM_382;
	logic [31:0] _RANDOM_383;
	logic [31:0] _RANDOM_384;
	logic [31:0] _RANDOM_385;
	logic [31:0] _RANDOM_386;
	logic [31:0] _RANDOM_387;
	logic [31:0] _RANDOM_388;
	logic [31:0] _RANDOM_389;
	logic [31:0] _RANDOM_390;
	logic [31:0] _RANDOM_391;
	logic [31:0] _RANDOM_392;
	logic [31:0] _RANDOM_393;
	logic [31:0] _RANDOM_394;
	logic [31:0] _RANDOM_395;
	logic [31:0] _RANDOM_396;
	logic [31:0] _RANDOM_397;
	logic [31:0] _RANDOM_398;
	logic [31:0] _RANDOM_399;
	logic [31:0] _RANDOM_400;
	logic [31:0] _RANDOM_401;
	logic [31:0] _RANDOM_402;
	logic [31:0] _RANDOM_403;
	logic [31:0] _RANDOM_404;
	logic [31:0] _RANDOM_405;
	logic [31:0] _RANDOM_406;
	logic [31:0] _RANDOM_407;
	logic [31:0] _RANDOM_408;
	logic [31:0] _RANDOM_409;
	logic [31:0] _RANDOM_410;
	logic [31:0] _RANDOM_411;
	logic [31:0] _RANDOM_412;
	logic [31:0] _RANDOM_413;
	logic [31:0] _RANDOM_414;
	logic [31:0] _RANDOM_415;
	logic [31:0] _RANDOM_416;
	logic [31:0] _RANDOM_417;
	logic [31:0] _RANDOM_418;
	logic [31:0] _RANDOM_419;
	logic [31:0] _RANDOM_420;
	logic [31:0] _RANDOM_421;
	logic [31:0] _RANDOM_422;
	logic [31:0] _RANDOM_423;
	logic [31:0] _RANDOM_424;
	logic [31:0] _RANDOM_425;
	logic [31:0] _RANDOM_426;
	logic [31:0] _RANDOM_427;
	logic [31:0] _RANDOM_428;
	logic [31:0] _RANDOM_429;
	logic [31:0] _RANDOM_430;
	logic [31:0] _RANDOM_431;
	logic [31:0] _RANDOM_432;
	logic [31:0] _RANDOM_433;
	logic [31:0] _RANDOM_434;
	logic [31:0] _RANDOM_435;
	logic [31:0] _RANDOM_436;
	logic [31:0] _RANDOM_437;
	logic [31:0] _RANDOM_438;
	logic [31:0] _RANDOM_439;
	logic [31:0] _RANDOM_440;
	logic [31:0] _RANDOM_441;
	logic [31:0] _RANDOM_442;
	logic [31:0] _RANDOM_443;
	logic [31:0] _RANDOM_444;
	logic [31:0] _RANDOM_445;
	logic [31:0] _RANDOM_446;
	logic [31:0] _RANDOM_447;
	logic [31:0] _RANDOM_448;
	logic [31:0] _RANDOM_449;
	logic [31:0] _RANDOM_450;
	logic [31:0] _RANDOM_451;
	logic [31:0] _RANDOM_452;
	logic [31:0] _RANDOM_453;
	logic [31:0] _RANDOM_454;
	logic [31:0] _RANDOM_455;
	logic [31:0] _RANDOM_456;
	logic [31:0] _RANDOM_457;
	logic [31:0] _RANDOM_458;
	logic [31:0] _RANDOM_459;
	logic [31:0] _RANDOM_460;
	logic [31:0] _RANDOM_461;
	logic [31:0] _RANDOM_462;
	logic [31:0] _RANDOM_463;
	logic [31:0] _RANDOM_464;
	logic [31:0] _RANDOM_465;
	logic [31:0] _RANDOM_466;
	logic [31:0] _RANDOM_467;
	logic [31:0] _RANDOM_468;
	logic [31:0] _RANDOM_469;
	logic [31:0] _RANDOM_470;
	logic [31:0] _RANDOM_471;
	logic [31:0] _RANDOM_472;
	logic [31:0] _RANDOM_473;
	logic [31:0] _RANDOM_474;
	logic [31:0] _RANDOM_475;
	logic [31:0] _RANDOM_476;
	logic [31:0] _RANDOM_477;
	logic [31:0] _RANDOM_478;
	logic [31:0] _RANDOM_479;
	logic [31:0] _RANDOM_480;
	logic [31:0] _RANDOM_481;
	logic [31:0] _RANDOM_482;
	logic [31:0] _RANDOM_483;
	logic [31:0] _RANDOM_484;
	logic [31:0] _RANDOM_485;
	logic [31:0] _RANDOM_486;
	logic [31:0] _RANDOM_487;
	logic [31:0] _RANDOM_488;
	logic [31:0] _RANDOM_489;
	logic [31:0] _RANDOM_490;
	logic [31:0] _RANDOM_491;
	logic [31:0] _RANDOM_492;
	logic [31:0] _RANDOM_493;
	logic [31:0] _RANDOM_494;
	logic [31:0] _RANDOM_495;
	logic [31:0] _RANDOM_496;
	logic [31:0] _RANDOM_497;
	logic [31:0] _RANDOM_498;
	logic [31:0] _RANDOM_499;
	logic [31:0] _RANDOM_500;
	logic [31:0] _RANDOM_501;
	logic [31:0] _RANDOM_502;
	logic [31:0] _RANDOM_503;
	logic [31:0] _RANDOM_504;
	logic [31:0] _RANDOM_505;
	logic [31:0] _RANDOM_506;
	logic [31:0] _RANDOM_507;
	logic [31:0] _RANDOM_508;
	logic [31:0] _RANDOM_509;
	logic [31:0] _RANDOM_510;
	logic [31:0] _RANDOM_511;
	logic [31:0] _RANDOM_512;
	logic [31:0] _RANDOM_513;
	logic [31:0] _RANDOM_514;
	logic [31:0] _RANDOM_515;
	logic [31:0] _RANDOM_516;
	logic [31:0] _RANDOM_517;
	logic [31:0] _RANDOM_518;
	logic [31:0] _RANDOM_519;
	logic [31:0] _RANDOM_520;
	logic [31:0] _RANDOM_521;
	logic [31:0] _RANDOM_522;
	logic [31:0] _RANDOM_523;
	logic [31:0] _RANDOM_524;
	logic [31:0] _RANDOM_525;
	logic [31:0] _RANDOM_526;
	logic [31:0] _RANDOM_527;
	logic [31:0] _RANDOM_528;
	logic [31:0] _RANDOM_529;
	logic [31:0] _RANDOM_530;
	logic [31:0] _RANDOM_531;
	logic [31:0] _RANDOM_532;
	logic [31:0] _RANDOM_533;
	logic [31:0] _RANDOM_534;
	logic [31:0] _RANDOM_535;
	logic [31:0] _RANDOM_536;
	logic [31:0] _RANDOM_537;
	logic [31:0] _RANDOM_538;
	logic [31:0] _RANDOM_539;
	logic [31:0] _RANDOM_540;
	logic [31:0] _RANDOM_541;
	logic [31:0] _RANDOM_542;
	logic [31:0] _RANDOM_543;
	logic [31:0] _RANDOM_544;
	logic [31:0] _RANDOM_545;
	logic [31:0] _RANDOM_546;
	logic [31:0] _RANDOM_547;
	logic [31:0] _RANDOM_548;
	logic [31:0] _RANDOM_549;
	logic [31:0] _RANDOM_550;
	logic [31:0] _RANDOM_551;
	logic [31:0] _RANDOM_552;
	logic [31:0] _RANDOM_553;
	logic [31:0] _RANDOM_554;
	logic [31:0] _RANDOM_555;
	logic [31:0] _RANDOM_556;
	logic [31:0] _RANDOM_557;
	logic [31:0] _RANDOM_558;
	logic [31:0] _RANDOM_559;
	logic [31:0] _RANDOM_560;
	logic [31:0] _RANDOM_561;
	logic [31:0] _RANDOM_562;
	logic [31:0] _RANDOM_563;
	logic [31:0] _RANDOM_564;
	logic [31:0] _RANDOM_565;
	logic [31:0] _RANDOM_566;
	logic [31:0] _RANDOM_567;
	logic [31:0] _RANDOM_568;
	logic [31:0] _RANDOM_569;
	logic [31:0] _RANDOM_570;
	logic [31:0] _RANDOM_571;
	logic [31:0] _RANDOM_572;
	logic [31:0] _RANDOM_573;
	logic [31:0] _RANDOM_574;
	logic [31:0] _RANDOM_575;
	logic [31:0] _RANDOM_576;
	logic [31:0] _RANDOM_577;
	logic [31:0] _RANDOM_578;
	logic [31:0] _RANDOM_579;
	logic [31:0] _RANDOM_580;
	logic [31:0] _RANDOM_581;
	logic [31:0] _RANDOM_582;
	logic [31:0] _RANDOM_583;
	logic [31:0] _RANDOM_584;
	logic [31:0] _RANDOM_585;
	logic [31:0] _RANDOM_586;
	logic [31:0] _RANDOM_587;
	logic [31:0] _RANDOM_588;
	logic [31:0] _RANDOM_589;
	logic [31:0] _RANDOM_590;
	logic [31:0] _RANDOM_591;
	logic [31:0] _RANDOM_592;
	logic [31:0] _RANDOM_593;
	logic [31:0] _RANDOM_594;
	logic [31:0] _RANDOM_595;
	logic [31:0] _RANDOM_596;
	logic [31:0] _RANDOM_597;
	logic [31:0] _RANDOM_598;
	logic [31:0] _RANDOM_599;
	logic [31:0] _RANDOM_600;
	logic [31:0] _RANDOM_601;
	logic [31:0] _RANDOM_602;
	logic [31:0] _RANDOM_603;
	logic [31:0] _RANDOM_604;
	logic [31:0] _RANDOM_605;
	logic [31:0] _RANDOM_606;
	logic [31:0] _RANDOM_607;
	logic [31:0] _RANDOM_608;
	logic [31:0] _RANDOM_609;
	logic [31:0] _RANDOM_610;
	logic [31:0] _RANDOM_611;
	logic [31:0] _RANDOM_612;
	logic [31:0] _RANDOM_613;
	logic [31:0] _RANDOM_614;
	logic [31:0] _RANDOM_615;
	logic [31:0] _RANDOM_616;
	logic [31:0] _RANDOM_617;
	logic [31:0] _RANDOM_618;
	logic [31:0] _RANDOM_619;
	logic [31:0] _RANDOM_620;
	logic [31:0] _RANDOM_621;
	logic [31:0] _RANDOM_622;
	logic [31:0] _RANDOM_623;
	logic [31:0] _RANDOM_624;
	logic [31:0] _RANDOM_625;
	logic [31:0] _RANDOM_626;
	logic [31:0] _RANDOM_627;
	logic [31:0] _RANDOM_628;
	logic [31:0] _RANDOM_629;
	logic [31:0] _RANDOM_630;
	logic [31:0] _RANDOM_631;
	logic [31:0] _RANDOM_632;
	logic [31:0] _RANDOM_633;
	logic [31:0] _RANDOM_634;
	logic [31:0] _RANDOM_635;
	logic [31:0] _RANDOM_636;
	logic [31:0] _RANDOM_637;
	logic [31:0] _RANDOM_638;
	logic [31:0] _RANDOM_639;
	logic [31:0] _RANDOM_640;
	logic [31:0] _RANDOM_641;
	logic [31:0] _RANDOM_642;
	logic [31:0] _RANDOM_643;
	logic [31:0] _RANDOM_644;
	logic [31:0] _RANDOM_645;
	logic [31:0] _RANDOM_646;
	logic [31:0] _RANDOM_647;
	logic [31:0] _RANDOM_648;
	logic [31:0] _RANDOM_649;
	logic [31:0] _RANDOM_650;
	logic [31:0] _RANDOM_651;
	logic [31:0] _RANDOM_652;
	logic [31:0] _RANDOM_653;
	logic [31:0] _RANDOM_654;
	logic [31:0] _RANDOM_655;
	logic [31:0] _RANDOM_656;
	logic [31:0] _RANDOM_657;
	logic [31:0] _RANDOM_658;
	logic [31:0] _RANDOM_659;
	logic [31:0] _RANDOM_660;
	logic [31:0] _RANDOM_661;
	logic [31:0] _RANDOM_662;
	logic [31:0] _RANDOM_663;
	logic [31:0] _RANDOM_664;
	logic [31:0] _RANDOM_665;
	logic [31:0] _RANDOM_666;
	logic [31:0] _RANDOM_667;
	logic [31:0] _RANDOM_668;
	logic [31:0] _RANDOM_669;
	logic [31:0] _RANDOM_670;
	logic [31:0] _RANDOM_671;
	logic [31:0] _RANDOM_672;
	logic [31:0] _RANDOM_673;
	logic [31:0] _RANDOM_674;
	logic [31:0] _RANDOM_675;
	logic [31:0] _RANDOM_676;
	logic [31:0] _RANDOM_677;
	logic [31:0] _RANDOM_678;
	logic [31:0] _RANDOM_679;
	logic [31:0] _RANDOM_680;
	logic [31:0] _RANDOM_681;
	logic [31:0] _RANDOM_682;
	logic [31:0] _RANDOM_683;
	logic [31:0] _RANDOM_684;
	logic [31:0] _RANDOM_685;
	logic [31:0] _RANDOM_686;
	logic [31:0] _RANDOM_687;
	logic [31:0] _RANDOM_688;
	logic [31:0] _RANDOM_689;
	logic [31:0] _RANDOM_690;
	logic [31:0] _RANDOM_691;
	logic [31:0] _RANDOM_692;
	logic [31:0] _RANDOM_693;
	logic [31:0] _RANDOM_694;
	logic [31:0] _RANDOM_695;
	logic [31:0] _RANDOM_696;
	logic [31:0] _RANDOM_697;
	logic [31:0] _RANDOM_698;
	logic [31:0] _RANDOM_699;
	logic [31:0] _RANDOM_700;
	logic [31:0] _RANDOM_701;
	logic [31:0] _RANDOM_702;
	logic [31:0] _RANDOM_703;
	logic [31:0] _RANDOM_704;
	logic [31:0] _RANDOM_705;
	logic [31:0] _RANDOM_706;
	logic [31:0] _RANDOM_707;
	logic [31:0] _RANDOM_708;
	logic [31:0] _RANDOM_709;
	logic [31:0] _RANDOM_710;
	logic [31:0] _RANDOM_711;
	logic [31:0] _RANDOM_712;
	logic [31:0] _RANDOM_713;
	logic [31:0] _RANDOM_714;
	logic [31:0] _RANDOM_715;
	logic [31:0] _RANDOM_716;
	logic [31:0] _RANDOM_717;
	logic [31:0] _RANDOM_718;
	logic [31:0] _RANDOM_719;
	logic [31:0] _RANDOM_720;
	logic [31:0] _RANDOM_721;
	logic [31:0] _RANDOM_722;
	logic [31:0] _RANDOM_723;
	logic [31:0] _RANDOM_724;
	logic [31:0] _RANDOM_725;
	logic [31:0] _RANDOM_726;
	logic [31:0] _RANDOM_727;
	logic [31:0] _RANDOM_728;
	logic [31:0] _RANDOM_729;
	logic [31:0] _RANDOM_730;
	logic [31:0] _RANDOM_731;
	logic [31:0] _RANDOM_732;
	logic [31:0] _RANDOM_733;
	logic [31:0] _RANDOM_734;
	logic [31:0] _RANDOM_735;
	logic [31:0] _RANDOM_736;
	logic [31:0] _RANDOM_737;
	logic [31:0] _RANDOM_738;
	logic [31:0] _RANDOM_739;
	logic [31:0] _RANDOM_740;
	logic [31:0] _RANDOM_741;
	logic [31:0] _RANDOM_742;
	logic [31:0] _RANDOM_743;
	logic [31:0] _RANDOM_744;
	logic [31:0] _RANDOM_745;
	logic [31:0] _RANDOM_746;
	logic [31:0] _RANDOM_747;
	logic [31:0] _RANDOM_748;
	logic [31:0] _RANDOM_749;
	logic [31:0] _RANDOM_750;
	logic [31:0] _RANDOM_751;
	logic [31:0] _RANDOM_752;
	logic [31:0] _RANDOM_753;
	logic [31:0] _RANDOM_754;
	logic [31:0] _RANDOM_755;
	logic [31:0] _RANDOM_756;
	logic [31:0] _RANDOM_757;
	logic [31:0] _RANDOM_758;
	logic [31:0] _RANDOM_759;
	logic [31:0] _RANDOM_760;
	logic [31:0] _RANDOM_761;
	logic [31:0] _RANDOM_762;
	logic [31:0] _RANDOM_763;
	logic [31:0] _RANDOM_764;
	logic [31:0] _RANDOM_765;
	logic [31:0] _RANDOM_766;
	logic [31:0] _RANDOM_767;
	logic [31:0] _RANDOM_768;
	logic [31:0] _RANDOM_769;
	logic [31:0] _RANDOM_770;
	logic [31:0] _RANDOM_771;
	logic [31:0] _RANDOM_772;
	logic [31:0] _RANDOM_773;
	logic [31:0] _RANDOM_774;
	logic [31:0] _RANDOM_775;
	logic [31:0] _RANDOM_776;
	logic [31:0] _RANDOM_777;
	logic [31:0] _RANDOM_778;
	logic [31:0] _RANDOM_779;
	logic [31:0] _RANDOM_780;
	logic [31:0] _RANDOM_781;
	logic [31:0] _RANDOM_782;
	logic [31:0] _RANDOM_783;
	logic [31:0] _RANDOM_784;
	logic [31:0] _RANDOM_785;
	logic [31:0] _RANDOM_786;
	logic [31:0] _RANDOM_787;
	logic [31:0] _RANDOM_788;
	logic [31:0] _RANDOM_789;
	logic [31:0] _RANDOM_790;
	logic [31:0] _RANDOM_791;
	logic [31:0] _RANDOM_792;
	logic [31:0] _RANDOM_793;
	logic [31:0] _RANDOM_794;
	logic [31:0] _RANDOM_795;
	logic [31:0] _RANDOM_796;
	logic [31:0] _RANDOM_797;
	logic [31:0] _RANDOM_798;
	logic [31:0] _RANDOM_799;
	logic [31:0] _RANDOM_800;
	logic [31:0] _RANDOM_801;
	logic [31:0] _RANDOM_802;
	logic [31:0] _RANDOM_803;
	logic [31:0] _RANDOM_804;
	logic [31:0] _RANDOM_805;
	logic [31:0] _RANDOM_806;
	logic [31:0] _RANDOM_807;
	logic [31:0] _RANDOM_808;
	logic [31:0] _RANDOM_809;
	logic [31:0] _RANDOM_810;
	logic [31:0] _RANDOM_811;
	logic [31:0] _RANDOM_812;
	logic [31:0] _RANDOM_813;
	logic [31:0] _RANDOM_814;
	logic [31:0] _RANDOM_815;
	logic [31:0] _RANDOM_816;
	logic [31:0] _RANDOM_817;
	logic [31:0] _RANDOM_818;
	logic [31:0] _RANDOM_819;
	logic [31:0] _RANDOM_820;
	logic [31:0] _RANDOM_821;
	logic [31:0] _RANDOM_822;
	logic [31:0] _RANDOM_823;
	logic [31:0] _RANDOM_824;
	logic [31:0] _RANDOM_825;
	logic [31:0] _RANDOM_826;
	logic [31:0] _RANDOM_827;
	logic [31:0] _RANDOM_828;
	logic [31:0] _RANDOM_829;
	logic [31:0] _RANDOM_830;
	logic [31:0] _RANDOM_831;
	logic [31:0] _RANDOM_832;
	logic [31:0] _RANDOM_833;
	logic [31:0] _RANDOM_834;
	logic [31:0] _RANDOM_835;
	logic [31:0] _RANDOM_836;
	logic [31:0] _RANDOM_837;
	logic [31:0] _RANDOM_838;
	logic [31:0] _RANDOM_839;
	logic [31:0] _RANDOM_840;
	logic [31:0] _RANDOM_841;
	logic [31:0] _RANDOM_842;
	logic [31:0] _RANDOM_843;
	logic [31:0] _RANDOM_844;
	logic [31:0] _RANDOM_845;
	logic [31:0] _RANDOM_846;
	logic [31:0] _RANDOM_847;
	logic [31:0] _RANDOM_848;
	logic [31:0] _RANDOM_849;
	logic [31:0] _RANDOM_850;
	logic [31:0] _RANDOM_851;
	logic [31:0] _RANDOM_852;
	logic [31:0] _RANDOM_853;
	logic [31:0] _RANDOM_854;
	logic [31:0] _RANDOM_855;
	logic [31:0] _RANDOM_856;
	logic [31:0] _RANDOM_857;
	logic [31:0] _RANDOM_858;
	logic [31:0] _RANDOM_859;
	logic [31:0] _RANDOM_860;
	logic [31:0] _RANDOM_861;
	logic [31:0] _RANDOM_862;
	logic [31:0] _RANDOM_863;
	logic [31:0] _RANDOM_864;
	logic [31:0] _RANDOM_865;
	logic [31:0] _RANDOM_866;
	logic [31:0] _RANDOM_867;
	logic [31:0] _RANDOM_868;
	logic [31:0] _RANDOM_869;
	logic [31:0] _RANDOM_870;
	logic [31:0] _RANDOM_871;
	logic [31:0] _RANDOM_872;
	logic [31:0] _RANDOM_873;
	logic [31:0] _RANDOM_874;
	logic [31:0] _RANDOM_875;
	logic [31:0] _RANDOM_876;
	logic [31:0] _RANDOM_877;
	logic [31:0] _RANDOM_878;
	logic [31:0] _RANDOM_879;
	logic [31:0] _RANDOM_880;
	logic [31:0] _RANDOM_881;
	logic [31:0] _RANDOM_882;
	logic [31:0] _RANDOM_883;
	logic [31:0] _RANDOM_884;
	logic [31:0] _RANDOM_885;
	logic [31:0] _RANDOM_886;
	logic [31:0] _RANDOM_887;
	logic [31:0] _RANDOM_888;
	logic [31:0] _RANDOM_889;
	logic [31:0] _RANDOM_890;
	logic [31:0] _RANDOM_891;
	logic [31:0] _RANDOM_892;
	logic [31:0] _RANDOM_893;
	logic [31:0] _RANDOM_894;
	logic [31:0] _RANDOM_895;
	logic [31:0] _RANDOM_896;
	logic [31:0] _RANDOM_897;
	logic [31:0] _RANDOM_898;
	logic [31:0] _RANDOM_899;
	logic [31:0] _RANDOM_900;
	logic [31:0] _RANDOM_901;
	logic [31:0] _RANDOM_902;
	logic [31:0] _RANDOM_903;
	logic [31:0] _RANDOM_904;
	logic [31:0] _RANDOM_905;
	logic [31:0] _RANDOM_906;
	logic [31:0] _RANDOM_907;
	logic [31:0] _RANDOM_908;
	logic [31:0] _RANDOM_909;
	logic [31:0] _RANDOM_910;
	logic [31:0] _RANDOM_911;
	logic [31:0] _RANDOM_912;
	logic [31:0] _RANDOM_913;
	logic [31:0] _RANDOM_914;
	logic [31:0] _RANDOM_915;
	logic [31:0] _RANDOM_916;
	logic [31:0] _RANDOM_917;
	logic [31:0] _RANDOM_918;
	logic [31:0] _RANDOM_919;
	logic [31:0] _RANDOM_920;
	logic [31:0] _RANDOM_921;
	logic [31:0] _RANDOM_922;
	logic [31:0] _RANDOM_923;
	logic [31:0] _RANDOM_924;
	logic [31:0] _RANDOM_925;
	logic [31:0] _RANDOM_926;
	logic [31:0] _RANDOM_927;
	logic [31:0] _RANDOM_928;
	logic [31:0] _RANDOM_929;
	logic [31:0] _RANDOM_930;
	logic [31:0] _RANDOM_931;
	logic [31:0] _RANDOM_932;
	logic [31:0] _RANDOM_933;
	logic [31:0] _RANDOM_934;
	logic [31:0] _RANDOM_935;
	logic [31:0] _RANDOM_936;
	logic [31:0] _RANDOM_937;
	logic [31:0] _RANDOM_938;
	logic [31:0] _RANDOM_939;
	logic [31:0] _RANDOM_940;
	logic [31:0] _RANDOM_941;
	Tile mesh_0_0(
		.clock(clock),
		.io_in_a_0(r_0),
		.io_in_b_0(b_0),
		.io_in_d_0(b_256_0),
		.io_in_control_0_dataflow(mesh_0_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_0_io_in_control_0_shift_b),
		.io_in_id_0(r_512_0),
		.io_in_last_0(r_768_0),
		.io_in_valid_0(r_256_0),
		.io_out_a_0(_mesh_0_0_io_out_a_0),
		.io_out_c_0(_mesh_0_0_io_out_c_0),
		.io_out_b_0(_mesh_0_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_0_io_out_id_0),
		.io_out_last_0(_mesh_0_0_io_out_last_0),
		.io_out_valid_0(_mesh_0_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2395 == GlobalFiModInstNr[0]) || (2395 == GlobalFiModInstNr[1]) || (2395 == GlobalFiModInstNr[2]) || (2395 == GlobalFiModInstNr[3]))));
	Tile mesh_0_1(
		.clock(clock),
		.io_in_a_0(r_1_0),
		.io_in_b_0(b_16_0),
		.io_in_d_0(b_272_0),
		.io_in_control_0_dataflow(mesh_0_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_1_io_in_control_0_shift_b),
		.io_in_id_0(r_528_0),
		.io_in_last_0(r_784_0),
		.io_in_valid_0(r_272_0),
		.io_out_a_0(_mesh_0_1_io_out_a_0),
		.io_out_c_0(_mesh_0_1_io_out_c_0),
		.io_out_b_0(_mesh_0_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_1_io_out_id_0),
		.io_out_last_0(_mesh_0_1_io_out_last_0),
		.io_out_valid_0(_mesh_0_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2396 == GlobalFiModInstNr[0]) || (2396 == GlobalFiModInstNr[1]) || (2396 == GlobalFiModInstNr[2]) || (2396 == GlobalFiModInstNr[3]))));
	Tile mesh_0_2(
		.clock(clock),
		.io_in_a_0(r_2_0),
		.io_in_b_0(b_32_0),
		.io_in_d_0(b_288_0),
		.io_in_control_0_dataflow(mesh_0_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_2_io_in_control_0_shift_b),
		.io_in_id_0(r_544_0),
		.io_in_last_0(r_800_0),
		.io_in_valid_0(r_288_0),
		.io_out_a_0(_mesh_0_2_io_out_a_0),
		.io_out_c_0(_mesh_0_2_io_out_c_0),
		.io_out_b_0(_mesh_0_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_2_io_out_id_0),
		.io_out_last_0(_mesh_0_2_io_out_last_0),
		.io_out_valid_0(_mesh_0_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2397 == GlobalFiModInstNr[0]) || (2397 == GlobalFiModInstNr[1]) || (2397 == GlobalFiModInstNr[2]) || (2397 == GlobalFiModInstNr[3]))));
	Tile mesh_0_3(
		.clock(clock),
		.io_in_a_0(r_3_0),
		.io_in_b_0(b_48_0),
		.io_in_d_0(b_304_0),
		.io_in_control_0_dataflow(mesh_0_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_3_io_in_control_0_shift_b),
		.io_in_id_0(r_560_0),
		.io_in_last_0(r_816_0),
		.io_in_valid_0(r_304_0),
		.io_out_a_0(_mesh_0_3_io_out_a_0),
		.io_out_c_0(_mesh_0_3_io_out_c_0),
		.io_out_b_0(_mesh_0_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_3_io_out_id_0),
		.io_out_last_0(_mesh_0_3_io_out_last_0),
		.io_out_valid_0(_mesh_0_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2398 == GlobalFiModInstNr[0]) || (2398 == GlobalFiModInstNr[1]) || (2398 == GlobalFiModInstNr[2]) || (2398 == GlobalFiModInstNr[3]))));
	Tile mesh_0_4(
		.clock(clock),
		.io_in_a_0(r_4_0),
		.io_in_b_0(b_64_0),
		.io_in_d_0(b_320_0),
		.io_in_control_0_dataflow(mesh_0_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_4_io_in_control_0_shift_b),
		.io_in_id_0(r_576_0),
		.io_in_last_0(r_832_0),
		.io_in_valid_0(r_320_0),
		.io_out_a_0(_mesh_0_4_io_out_a_0),
		.io_out_c_0(_mesh_0_4_io_out_c_0),
		.io_out_b_0(_mesh_0_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_4_io_out_id_0),
		.io_out_last_0(_mesh_0_4_io_out_last_0),
		.io_out_valid_0(_mesh_0_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2399 == GlobalFiModInstNr[0]) || (2399 == GlobalFiModInstNr[1]) || (2399 == GlobalFiModInstNr[2]) || (2399 == GlobalFiModInstNr[3]))));
	Tile mesh_0_5(
		.clock(clock),
		.io_in_a_0(r_5_0),
		.io_in_b_0(b_80_0),
		.io_in_d_0(b_336_0),
		.io_in_control_0_dataflow(mesh_0_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_5_io_in_control_0_shift_b),
		.io_in_id_0(r_592_0),
		.io_in_last_0(r_848_0),
		.io_in_valid_0(r_336_0),
		.io_out_a_0(_mesh_0_5_io_out_a_0),
		.io_out_c_0(_mesh_0_5_io_out_c_0),
		.io_out_b_0(_mesh_0_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_5_io_out_id_0),
		.io_out_last_0(_mesh_0_5_io_out_last_0),
		.io_out_valid_0(_mesh_0_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2400 == GlobalFiModInstNr[0]) || (2400 == GlobalFiModInstNr[1]) || (2400 == GlobalFiModInstNr[2]) || (2400 == GlobalFiModInstNr[3]))));
	Tile mesh_0_6(
		.clock(clock),
		.io_in_a_0(r_6_0),
		.io_in_b_0(b_96_0),
		.io_in_d_0(b_352_0),
		.io_in_control_0_dataflow(mesh_0_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_6_io_in_control_0_shift_b),
		.io_in_id_0(r_608_0),
		.io_in_last_0(r_864_0),
		.io_in_valid_0(r_352_0),
		.io_out_a_0(_mesh_0_6_io_out_a_0),
		.io_out_c_0(_mesh_0_6_io_out_c_0),
		.io_out_b_0(_mesh_0_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_6_io_out_id_0),
		.io_out_last_0(_mesh_0_6_io_out_last_0),
		.io_out_valid_0(_mesh_0_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2401 == GlobalFiModInstNr[0]) || (2401 == GlobalFiModInstNr[1]) || (2401 == GlobalFiModInstNr[2]) || (2401 == GlobalFiModInstNr[3]))));
	Tile mesh_0_7(
		.clock(clock),
		.io_in_a_0(r_7_0),
		.io_in_b_0(b_112_0),
		.io_in_d_0(b_368_0),
		.io_in_control_0_dataflow(mesh_0_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_7_io_in_control_0_shift_b),
		.io_in_id_0(r_624_0),
		.io_in_last_0(r_880_0),
		.io_in_valid_0(r_368_0),
		.io_out_a_0(_mesh_0_7_io_out_a_0),
		.io_out_c_0(_mesh_0_7_io_out_c_0),
		.io_out_b_0(_mesh_0_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_7_io_out_id_0),
		.io_out_last_0(_mesh_0_7_io_out_last_0),
		.io_out_valid_0(_mesh_0_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2402 == GlobalFiModInstNr[0]) || (2402 == GlobalFiModInstNr[1]) || (2402 == GlobalFiModInstNr[2]) || (2402 == GlobalFiModInstNr[3]))));
	Tile mesh_0_8(
		.clock(clock),
		.io_in_a_0(r_8_0),
		.io_in_b_0(b_128_0),
		.io_in_d_0(b_384_0),
		.io_in_control_0_dataflow(mesh_0_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_8_io_in_control_0_shift_b),
		.io_in_id_0(r_640_0),
		.io_in_last_0(r_896_0),
		.io_in_valid_0(r_384_0),
		.io_out_a_0(_mesh_0_8_io_out_a_0),
		.io_out_c_0(_mesh_0_8_io_out_c_0),
		.io_out_b_0(_mesh_0_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_8_io_out_id_0),
		.io_out_last_0(_mesh_0_8_io_out_last_0),
		.io_out_valid_0(_mesh_0_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2403 == GlobalFiModInstNr[0]) || (2403 == GlobalFiModInstNr[1]) || (2403 == GlobalFiModInstNr[2]) || (2403 == GlobalFiModInstNr[3]))));
	Tile mesh_0_9(
		.clock(clock),
		.io_in_a_0(r_9_0),
		.io_in_b_0(b_144_0),
		.io_in_d_0(b_400_0),
		.io_in_control_0_dataflow(mesh_0_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_9_io_in_control_0_shift_b),
		.io_in_id_0(r_656_0),
		.io_in_last_0(r_912_0),
		.io_in_valid_0(r_400_0),
		.io_out_a_0(_mesh_0_9_io_out_a_0),
		.io_out_c_0(_mesh_0_9_io_out_c_0),
		.io_out_b_0(_mesh_0_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_9_io_out_id_0),
		.io_out_last_0(_mesh_0_9_io_out_last_0),
		.io_out_valid_0(_mesh_0_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2404 == GlobalFiModInstNr[0]) || (2404 == GlobalFiModInstNr[1]) || (2404 == GlobalFiModInstNr[2]) || (2404 == GlobalFiModInstNr[3]))));
	Tile mesh_0_10(
		.clock(clock),
		.io_in_a_0(r_10_0),
		.io_in_b_0(b_160_0),
		.io_in_d_0(b_416_0),
		.io_in_control_0_dataflow(mesh_0_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_10_io_in_control_0_shift_b),
		.io_in_id_0(r_672_0),
		.io_in_last_0(r_928_0),
		.io_in_valid_0(r_416_0),
		.io_out_a_0(_mesh_0_10_io_out_a_0),
		.io_out_c_0(_mesh_0_10_io_out_c_0),
		.io_out_b_0(_mesh_0_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_10_io_out_id_0),
		.io_out_last_0(_mesh_0_10_io_out_last_0),
		.io_out_valid_0(_mesh_0_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2405 == GlobalFiModInstNr[0]) || (2405 == GlobalFiModInstNr[1]) || (2405 == GlobalFiModInstNr[2]) || (2405 == GlobalFiModInstNr[3]))));
	Tile mesh_0_11(
		.clock(clock),
		.io_in_a_0(r_11_0),
		.io_in_b_0(b_176_0),
		.io_in_d_0(b_432_0),
		.io_in_control_0_dataflow(mesh_0_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_11_io_in_control_0_shift_b),
		.io_in_id_0(r_688_0),
		.io_in_last_0(r_944_0),
		.io_in_valid_0(r_432_0),
		.io_out_a_0(_mesh_0_11_io_out_a_0),
		.io_out_c_0(_mesh_0_11_io_out_c_0),
		.io_out_b_0(_mesh_0_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_11_io_out_id_0),
		.io_out_last_0(_mesh_0_11_io_out_last_0),
		.io_out_valid_0(_mesh_0_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2406 == GlobalFiModInstNr[0]) || (2406 == GlobalFiModInstNr[1]) || (2406 == GlobalFiModInstNr[2]) || (2406 == GlobalFiModInstNr[3]))));
	Tile mesh_0_12(
		.clock(clock),
		.io_in_a_0(r_12_0),
		.io_in_b_0(b_192_0),
		.io_in_d_0(b_448_0),
		.io_in_control_0_dataflow(mesh_0_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_12_io_in_control_0_shift_b),
		.io_in_id_0(r_704_0),
		.io_in_last_0(r_960_0),
		.io_in_valid_0(r_448_0),
		.io_out_a_0(_mesh_0_12_io_out_a_0),
		.io_out_c_0(_mesh_0_12_io_out_c_0),
		.io_out_b_0(_mesh_0_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_12_io_out_id_0),
		.io_out_last_0(_mesh_0_12_io_out_last_0),
		.io_out_valid_0(_mesh_0_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2407 == GlobalFiModInstNr[0]) || (2407 == GlobalFiModInstNr[1]) || (2407 == GlobalFiModInstNr[2]) || (2407 == GlobalFiModInstNr[3]))));
	Tile mesh_0_13(
		.clock(clock),
		.io_in_a_0(r_13_0),
		.io_in_b_0(b_208_0),
		.io_in_d_0(b_464_0),
		.io_in_control_0_dataflow(mesh_0_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_13_io_in_control_0_shift_b),
		.io_in_id_0(r_720_0),
		.io_in_last_0(r_976_0),
		.io_in_valid_0(r_464_0),
		.io_out_a_0(_mesh_0_13_io_out_a_0),
		.io_out_c_0(_mesh_0_13_io_out_c_0),
		.io_out_b_0(_mesh_0_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_13_io_out_id_0),
		.io_out_last_0(_mesh_0_13_io_out_last_0),
		.io_out_valid_0(_mesh_0_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2408 == GlobalFiModInstNr[0]) || (2408 == GlobalFiModInstNr[1]) || (2408 == GlobalFiModInstNr[2]) || (2408 == GlobalFiModInstNr[3]))));
	Tile mesh_0_14(
		.clock(clock),
		.io_in_a_0(r_14_0),
		.io_in_b_0(b_224_0),
		.io_in_d_0(b_480_0),
		.io_in_control_0_dataflow(mesh_0_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_14_io_in_control_0_shift_b),
		.io_in_id_0(r_736_0),
		.io_in_last_0(r_992_0),
		.io_in_valid_0(r_480_0),
		.io_out_a_0(_mesh_0_14_io_out_a_0),
		.io_out_c_0(_mesh_0_14_io_out_c_0),
		.io_out_b_0(_mesh_0_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_14_io_out_id_0),
		.io_out_last_0(_mesh_0_14_io_out_last_0),
		.io_out_valid_0(_mesh_0_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2409 == GlobalFiModInstNr[0]) || (2409 == GlobalFiModInstNr[1]) || (2409 == GlobalFiModInstNr[2]) || (2409 == GlobalFiModInstNr[3]))));
	Tile mesh_0_15(
		.clock(clock),
		.io_in_a_0(r_15_0),
		.io_in_b_0(b_240_0),
		.io_in_d_0(b_496_0),
		.io_in_control_0_dataflow(mesh_0_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_15_io_in_control_0_shift_b),
		.io_in_id_0(r_752_0),
		.io_in_last_0(r_1008_0),
		.io_in_valid_0(r_496_0),
		.io_out_a_0(_mesh_0_15_io_out_a_0),
		.io_out_c_0(_mesh_0_15_io_out_c_0),
		.io_out_b_0(_mesh_0_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_15_io_out_id_0),
		.io_out_last_0(_mesh_0_15_io_out_last_0),
		.io_out_valid_0(_mesh_0_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2410 == GlobalFiModInstNr[0]) || (2410 == GlobalFiModInstNr[1]) || (2410 == GlobalFiModInstNr[2]) || (2410 == GlobalFiModInstNr[3]))));
	Tile mesh_1_0(
		.clock(clock),
		.io_in_a_0(r_16_0),
		.io_in_b_0(b_1_0),
		.io_in_d_0(b_257_0),
		.io_in_control_0_dataflow(mesh_1_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_0_io_in_control_0_shift_b),
		.io_in_id_0(r_513_0),
		.io_in_last_0(r_769_0),
		.io_in_valid_0(r_257_0),
		.io_out_a_0(_mesh_1_0_io_out_a_0),
		.io_out_c_0(_mesh_1_0_io_out_c_0),
		.io_out_b_0(_mesh_1_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_0_io_out_id_0),
		.io_out_last_0(_mesh_1_0_io_out_last_0),
		.io_out_valid_0(_mesh_1_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2411 == GlobalFiModInstNr[0]) || (2411 == GlobalFiModInstNr[1]) || (2411 == GlobalFiModInstNr[2]) || (2411 == GlobalFiModInstNr[3]))));
	Tile mesh_1_1(
		.clock(clock),
		.io_in_a_0(r_17_0),
		.io_in_b_0(b_17_0),
		.io_in_d_0(b_273_0),
		.io_in_control_0_dataflow(mesh_1_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_1_io_in_control_0_shift_b),
		.io_in_id_0(r_529_0),
		.io_in_last_0(r_785_0),
		.io_in_valid_0(r_273_0),
		.io_out_a_0(_mesh_1_1_io_out_a_0),
		.io_out_c_0(_mesh_1_1_io_out_c_0),
		.io_out_b_0(_mesh_1_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_1_io_out_id_0),
		.io_out_last_0(_mesh_1_1_io_out_last_0),
		.io_out_valid_0(_mesh_1_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2412 == GlobalFiModInstNr[0]) || (2412 == GlobalFiModInstNr[1]) || (2412 == GlobalFiModInstNr[2]) || (2412 == GlobalFiModInstNr[3]))));
	Tile mesh_1_2(
		.clock(clock),
		.io_in_a_0(r_18_0),
		.io_in_b_0(b_33_0),
		.io_in_d_0(b_289_0),
		.io_in_control_0_dataflow(mesh_1_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_2_io_in_control_0_shift_b),
		.io_in_id_0(r_545_0),
		.io_in_last_0(r_801_0),
		.io_in_valid_0(r_289_0),
		.io_out_a_0(_mesh_1_2_io_out_a_0),
		.io_out_c_0(_mesh_1_2_io_out_c_0),
		.io_out_b_0(_mesh_1_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_2_io_out_id_0),
		.io_out_last_0(_mesh_1_2_io_out_last_0),
		.io_out_valid_0(_mesh_1_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2413 == GlobalFiModInstNr[0]) || (2413 == GlobalFiModInstNr[1]) || (2413 == GlobalFiModInstNr[2]) || (2413 == GlobalFiModInstNr[3]))));
	Tile mesh_1_3(
		.clock(clock),
		.io_in_a_0(r_19_0),
		.io_in_b_0(b_49_0),
		.io_in_d_0(b_305_0),
		.io_in_control_0_dataflow(mesh_1_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_3_io_in_control_0_shift_b),
		.io_in_id_0(r_561_0),
		.io_in_last_0(r_817_0),
		.io_in_valid_0(r_305_0),
		.io_out_a_0(_mesh_1_3_io_out_a_0),
		.io_out_c_0(_mesh_1_3_io_out_c_0),
		.io_out_b_0(_mesh_1_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_3_io_out_id_0),
		.io_out_last_0(_mesh_1_3_io_out_last_0),
		.io_out_valid_0(_mesh_1_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2414 == GlobalFiModInstNr[0]) || (2414 == GlobalFiModInstNr[1]) || (2414 == GlobalFiModInstNr[2]) || (2414 == GlobalFiModInstNr[3]))));
	Tile mesh_1_4(
		.clock(clock),
		.io_in_a_0(r_20_0),
		.io_in_b_0(b_65_0),
		.io_in_d_0(b_321_0),
		.io_in_control_0_dataflow(mesh_1_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_4_io_in_control_0_shift_b),
		.io_in_id_0(r_577_0),
		.io_in_last_0(r_833_0),
		.io_in_valid_0(r_321_0),
		.io_out_a_0(_mesh_1_4_io_out_a_0),
		.io_out_c_0(_mesh_1_4_io_out_c_0),
		.io_out_b_0(_mesh_1_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_4_io_out_id_0),
		.io_out_last_0(_mesh_1_4_io_out_last_0),
		.io_out_valid_0(_mesh_1_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2415 == GlobalFiModInstNr[0]) || (2415 == GlobalFiModInstNr[1]) || (2415 == GlobalFiModInstNr[2]) || (2415 == GlobalFiModInstNr[3]))));
	Tile mesh_1_5(
		.clock(clock),
		.io_in_a_0(r_21_0),
		.io_in_b_0(b_81_0),
		.io_in_d_0(b_337_0),
		.io_in_control_0_dataflow(mesh_1_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_5_io_in_control_0_shift_b),
		.io_in_id_0(r_593_0),
		.io_in_last_0(r_849_0),
		.io_in_valid_0(r_337_0),
		.io_out_a_0(_mesh_1_5_io_out_a_0),
		.io_out_c_0(_mesh_1_5_io_out_c_0),
		.io_out_b_0(_mesh_1_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_5_io_out_id_0),
		.io_out_last_0(_mesh_1_5_io_out_last_0),
		.io_out_valid_0(_mesh_1_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2416 == GlobalFiModInstNr[0]) || (2416 == GlobalFiModInstNr[1]) || (2416 == GlobalFiModInstNr[2]) || (2416 == GlobalFiModInstNr[3]))));
	Tile mesh_1_6(
		.clock(clock),
		.io_in_a_0(r_22_0),
		.io_in_b_0(b_97_0),
		.io_in_d_0(b_353_0),
		.io_in_control_0_dataflow(mesh_1_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_6_io_in_control_0_shift_b),
		.io_in_id_0(r_609_0),
		.io_in_last_0(r_865_0),
		.io_in_valid_0(r_353_0),
		.io_out_a_0(_mesh_1_6_io_out_a_0),
		.io_out_c_0(_mesh_1_6_io_out_c_0),
		.io_out_b_0(_mesh_1_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_6_io_out_id_0),
		.io_out_last_0(_mesh_1_6_io_out_last_0),
		.io_out_valid_0(_mesh_1_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2417 == GlobalFiModInstNr[0]) || (2417 == GlobalFiModInstNr[1]) || (2417 == GlobalFiModInstNr[2]) || (2417 == GlobalFiModInstNr[3]))));
	Tile mesh_1_7(
		.clock(clock),
		.io_in_a_0(r_23_0),
		.io_in_b_0(b_113_0),
		.io_in_d_0(b_369_0),
		.io_in_control_0_dataflow(mesh_1_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_7_io_in_control_0_shift_b),
		.io_in_id_0(r_625_0),
		.io_in_last_0(r_881_0),
		.io_in_valid_0(r_369_0),
		.io_out_a_0(_mesh_1_7_io_out_a_0),
		.io_out_c_0(_mesh_1_7_io_out_c_0),
		.io_out_b_0(_mesh_1_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_7_io_out_id_0),
		.io_out_last_0(_mesh_1_7_io_out_last_0),
		.io_out_valid_0(_mesh_1_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2418 == GlobalFiModInstNr[0]) || (2418 == GlobalFiModInstNr[1]) || (2418 == GlobalFiModInstNr[2]) || (2418 == GlobalFiModInstNr[3]))));
	Tile mesh_1_8(
		.clock(clock),
		.io_in_a_0(r_24_0),
		.io_in_b_0(b_129_0),
		.io_in_d_0(b_385_0),
		.io_in_control_0_dataflow(mesh_1_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_8_io_in_control_0_shift_b),
		.io_in_id_0(r_641_0),
		.io_in_last_0(r_897_0),
		.io_in_valid_0(r_385_0),
		.io_out_a_0(_mesh_1_8_io_out_a_0),
		.io_out_c_0(_mesh_1_8_io_out_c_0),
		.io_out_b_0(_mesh_1_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_8_io_out_id_0),
		.io_out_last_0(_mesh_1_8_io_out_last_0),
		.io_out_valid_0(_mesh_1_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2419 == GlobalFiModInstNr[0]) || (2419 == GlobalFiModInstNr[1]) || (2419 == GlobalFiModInstNr[2]) || (2419 == GlobalFiModInstNr[3]))));
	Tile mesh_1_9(
		.clock(clock),
		.io_in_a_0(r_25_0),
		.io_in_b_0(b_145_0),
		.io_in_d_0(b_401_0),
		.io_in_control_0_dataflow(mesh_1_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_9_io_in_control_0_shift_b),
		.io_in_id_0(r_657_0),
		.io_in_last_0(r_913_0),
		.io_in_valid_0(r_401_0),
		.io_out_a_0(_mesh_1_9_io_out_a_0),
		.io_out_c_0(_mesh_1_9_io_out_c_0),
		.io_out_b_0(_mesh_1_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_9_io_out_id_0),
		.io_out_last_0(_mesh_1_9_io_out_last_0),
		.io_out_valid_0(_mesh_1_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2420 == GlobalFiModInstNr[0]) || (2420 == GlobalFiModInstNr[1]) || (2420 == GlobalFiModInstNr[2]) || (2420 == GlobalFiModInstNr[3]))));
	Tile mesh_1_10(
		.clock(clock),
		.io_in_a_0(r_26_0),
		.io_in_b_0(b_161_0),
		.io_in_d_0(b_417_0),
		.io_in_control_0_dataflow(mesh_1_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_10_io_in_control_0_shift_b),
		.io_in_id_0(r_673_0),
		.io_in_last_0(r_929_0),
		.io_in_valid_0(r_417_0),
		.io_out_a_0(_mesh_1_10_io_out_a_0),
		.io_out_c_0(_mesh_1_10_io_out_c_0),
		.io_out_b_0(_mesh_1_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_10_io_out_id_0),
		.io_out_last_0(_mesh_1_10_io_out_last_0),
		.io_out_valid_0(_mesh_1_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2421 == GlobalFiModInstNr[0]) || (2421 == GlobalFiModInstNr[1]) || (2421 == GlobalFiModInstNr[2]) || (2421 == GlobalFiModInstNr[3]))));
	Tile mesh_1_11(
		.clock(clock),
		.io_in_a_0(r_27_0),
		.io_in_b_0(b_177_0),
		.io_in_d_0(b_433_0),
		.io_in_control_0_dataflow(mesh_1_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_11_io_in_control_0_shift_b),
		.io_in_id_0(r_689_0),
		.io_in_last_0(r_945_0),
		.io_in_valid_0(r_433_0),
		.io_out_a_0(_mesh_1_11_io_out_a_0),
		.io_out_c_0(_mesh_1_11_io_out_c_0),
		.io_out_b_0(_mesh_1_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_11_io_out_id_0),
		.io_out_last_0(_mesh_1_11_io_out_last_0),
		.io_out_valid_0(_mesh_1_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2422 == GlobalFiModInstNr[0]) || (2422 == GlobalFiModInstNr[1]) || (2422 == GlobalFiModInstNr[2]) || (2422 == GlobalFiModInstNr[3]))));
	Tile mesh_1_12(
		.clock(clock),
		.io_in_a_0(r_28_0),
		.io_in_b_0(b_193_0),
		.io_in_d_0(b_449_0),
		.io_in_control_0_dataflow(mesh_1_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_12_io_in_control_0_shift_b),
		.io_in_id_0(r_705_0),
		.io_in_last_0(r_961_0),
		.io_in_valid_0(r_449_0),
		.io_out_a_0(_mesh_1_12_io_out_a_0),
		.io_out_c_0(_mesh_1_12_io_out_c_0),
		.io_out_b_0(_mesh_1_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_12_io_out_id_0),
		.io_out_last_0(_mesh_1_12_io_out_last_0),
		.io_out_valid_0(_mesh_1_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2423 == GlobalFiModInstNr[0]) || (2423 == GlobalFiModInstNr[1]) || (2423 == GlobalFiModInstNr[2]) || (2423 == GlobalFiModInstNr[3]))));
	Tile mesh_1_13(
		.clock(clock),
		.io_in_a_0(r_29_0),
		.io_in_b_0(b_209_0),
		.io_in_d_0(b_465_0),
		.io_in_control_0_dataflow(mesh_1_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_13_io_in_control_0_shift_b),
		.io_in_id_0(r_721_0),
		.io_in_last_0(r_977_0),
		.io_in_valid_0(r_465_0),
		.io_out_a_0(_mesh_1_13_io_out_a_0),
		.io_out_c_0(_mesh_1_13_io_out_c_0),
		.io_out_b_0(_mesh_1_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_13_io_out_id_0),
		.io_out_last_0(_mesh_1_13_io_out_last_0),
		.io_out_valid_0(_mesh_1_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2424 == GlobalFiModInstNr[0]) || (2424 == GlobalFiModInstNr[1]) || (2424 == GlobalFiModInstNr[2]) || (2424 == GlobalFiModInstNr[3]))));
	Tile mesh_1_14(
		.clock(clock),
		.io_in_a_0(r_30_0),
		.io_in_b_0(b_225_0),
		.io_in_d_0(b_481_0),
		.io_in_control_0_dataflow(mesh_1_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_14_io_in_control_0_shift_b),
		.io_in_id_0(r_737_0),
		.io_in_last_0(r_993_0),
		.io_in_valid_0(r_481_0),
		.io_out_a_0(_mesh_1_14_io_out_a_0),
		.io_out_c_0(_mesh_1_14_io_out_c_0),
		.io_out_b_0(_mesh_1_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_14_io_out_id_0),
		.io_out_last_0(_mesh_1_14_io_out_last_0),
		.io_out_valid_0(_mesh_1_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2425 == GlobalFiModInstNr[0]) || (2425 == GlobalFiModInstNr[1]) || (2425 == GlobalFiModInstNr[2]) || (2425 == GlobalFiModInstNr[3]))));
	Tile mesh_1_15(
		.clock(clock),
		.io_in_a_0(r_31_0),
		.io_in_b_0(b_241_0),
		.io_in_d_0(b_497_0),
		.io_in_control_0_dataflow(mesh_1_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_15_io_in_control_0_shift_b),
		.io_in_id_0(r_753_0),
		.io_in_last_0(r_1009_0),
		.io_in_valid_0(r_497_0),
		.io_out_a_0(_mesh_1_15_io_out_a_0),
		.io_out_c_0(_mesh_1_15_io_out_c_0),
		.io_out_b_0(_mesh_1_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_15_io_out_id_0),
		.io_out_last_0(_mesh_1_15_io_out_last_0),
		.io_out_valid_0(_mesh_1_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2426 == GlobalFiModInstNr[0]) || (2426 == GlobalFiModInstNr[1]) || (2426 == GlobalFiModInstNr[2]) || (2426 == GlobalFiModInstNr[3]))));
	Tile mesh_2_0(
		.clock(clock),
		.io_in_a_0(r_32_0),
		.io_in_b_0(b_2_0),
		.io_in_d_0(b_258_0),
		.io_in_control_0_dataflow(mesh_2_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_0_io_in_control_0_shift_b),
		.io_in_id_0(r_514_0),
		.io_in_last_0(r_770_0),
		.io_in_valid_0(r_258_0),
		.io_out_a_0(_mesh_2_0_io_out_a_0),
		.io_out_c_0(_mesh_2_0_io_out_c_0),
		.io_out_b_0(_mesh_2_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_0_io_out_id_0),
		.io_out_last_0(_mesh_2_0_io_out_last_0),
		.io_out_valid_0(_mesh_2_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2427 == GlobalFiModInstNr[0]) || (2427 == GlobalFiModInstNr[1]) || (2427 == GlobalFiModInstNr[2]) || (2427 == GlobalFiModInstNr[3]))));
	Tile mesh_2_1(
		.clock(clock),
		.io_in_a_0(r_33_0),
		.io_in_b_0(b_18_0),
		.io_in_d_0(b_274_0),
		.io_in_control_0_dataflow(mesh_2_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_1_io_in_control_0_shift_b),
		.io_in_id_0(r_530_0),
		.io_in_last_0(r_786_0),
		.io_in_valid_0(r_274_0),
		.io_out_a_0(_mesh_2_1_io_out_a_0),
		.io_out_c_0(_mesh_2_1_io_out_c_0),
		.io_out_b_0(_mesh_2_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_1_io_out_id_0),
		.io_out_last_0(_mesh_2_1_io_out_last_0),
		.io_out_valid_0(_mesh_2_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2428 == GlobalFiModInstNr[0]) || (2428 == GlobalFiModInstNr[1]) || (2428 == GlobalFiModInstNr[2]) || (2428 == GlobalFiModInstNr[3]))));
	Tile mesh_2_2(
		.clock(clock),
		.io_in_a_0(r_34_0),
		.io_in_b_0(b_34_0),
		.io_in_d_0(b_290_0),
		.io_in_control_0_dataflow(mesh_2_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_2_io_in_control_0_shift_b),
		.io_in_id_0(r_546_0),
		.io_in_last_0(r_802_0),
		.io_in_valid_0(r_290_0),
		.io_out_a_0(_mesh_2_2_io_out_a_0),
		.io_out_c_0(_mesh_2_2_io_out_c_0),
		.io_out_b_0(_mesh_2_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_2_io_out_id_0),
		.io_out_last_0(_mesh_2_2_io_out_last_0),
		.io_out_valid_0(_mesh_2_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2429 == GlobalFiModInstNr[0]) || (2429 == GlobalFiModInstNr[1]) || (2429 == GlobalFiModInstNr[2]) || (2429 == GlobalFiModInstNr[3]))));
	Tile mesh_2_3(
		.clock(clock),
		.io_in_a_0(r_35_0),
		.io_in_b_0(b_50_0),
		.io_in_d_0(b_306_0),
		.io_in_control_0_dataflow(mesh_2_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_3_io_in_control_0_shift_b),
		.io_in_id_0(r_562_0),
		.io_in_last_0(r_818_0),
		.io_in_valid_0(r_306_0),
		.io_out_a_0(_mesh_2_3_io_out_a_0),
		.io_out_c_0(_mesh_2_3_io_out_c_0),
		.io_out_b_0(_mesh_2_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_3_io_out_id_0),
		.io_out_last_0(_mesh_2_3_io_out_last_0),
		.io_out_valid_0(_mesh_2_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2430 == GlobalFiModInstNr[0]) || (2430 == GlobalFiModInstNr[1]) || (2430 == GlobalFiModInstNr[2]) || (2430 == GlobalFiModInstNr[3]))));
	Tile mesh_2_4(
		.clock(clock),
		.io_in_a_0(r_36_0),
		.io_in_b_0(b_66_0),
		.io_in_d_0(b_322_0),
		.io_in_control_0_dataflow(mesh_2_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_4_io_in_control_0_shift_b),
		.io_in_id_0(r_578_0),
		.io_in_last_0(r_834_0),
		.io_in_valid_0(r_322_0),
		.io_out_a_0(_mesh_2_4_io_out_a_0),
		.io_out_c_0(_mesh_2_4_io_out_c_0),
		.io_out_b_0(_mesh_2_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_4_io_out_id_0),
		.io_out_last_0(_mesh_2_4_io_out_last_0),
		.io_out_valid_0(_mesh_2_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2431 == GlobalFiModInstNr[0]) || (2431 == GlobalFiModInstNr[1]) || (2431 == GlobalFiModInstNr[2]) || (2431 == GlobalFiModInstNr[3]))));
	Tile mesh_2_5(
		.clock(clock),
		.io_in_a_0(r_37_0),
		.io_in_b_0(b_82_0),
		.io_in_d_0(b_338_0),
		.io_in_control_0_dataflow(mesh_2_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_5_io_in_control_0_shift_b),
		.io_in_id_0(r_594_0),
		.io_in_last_0(r_850_0),
		.io_in_valid_0(r_338_0),
		.io_out_a_0(_mesh_2_5_io_out_a_0),
		.io_out_c_0(_mesh_2_5_io_out_c_0),
		.io_out_b_0(_mesh_2_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_5_io_out_id_0),
		.io_out_last_0(_mesh_2_5_io_out_last_0),
		.io_out_valid_0(_mesh_2_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2432 == GlobalFiModInstNr[0]) || (2432 == GlobalFiModInstNr[1]) || (2432 == GlobalFiModInstNr[2]) || (2432 == GlobalFiModInstNr[3]))));
	Tile mesh_2_6(
		.clock(clock),
		.io_in_a_0(r_38_0),
		.io_in_b_0(b_98_0),
		.io_in_d_0(b_354_0),
		.io_in_control_0_dataflow(mesh_2_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_6_io_in_control_0_shift_b),
		.io_in_id_0(r_610_0),
		.io_in_last_0(r_866_0),
		.io_in_valid_0(r_354_0),
		.io_out_a_0(_mesh_2_6_io_out_a_0),
		.io_out_c_0(_mesh_2_6_io_out_c_0),
		.io_out_b_0(_mesh_2_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_6_io_out_id_0),
		.io_out_last_0(_mesh_2_6_io_out_last_0),
		.io_out_valid_0(_mesh_2_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2433 == GlobalFiModInstNr[0]) || (2433 == GlobalFiModInstNr[1]) || (2433 == GlobalFiModInstNr[2]) || (2433 == GlobalFiModInstNr[3]))));
	Tile mesh_2_7(
		.clock(clock),
		.io_in_a_0(r_39_0),
		.io_in_b_0(b_114_0),
		.io_in_d_0(b_370_0),
		.io_in_control_0_dataflow(mesh_2_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_7_io_in_control_0_shift_b),
		.io_in_id_0(r_626_0),
		.io_in_last_0(r_882_0),
		.io_in_valid_0(r_370_0),
		.io_out_a_0(_mesh_2_7_io_out_a_0),
		.io_out_c_0(_mesh_2_7_io_out_c_0),
		.io_out_b_0(_mesh_2_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_7_io_out_id_0),
		.io_out_last_0(_mesh_2_7_io_out_last_0),
		.io_out_valid_0(_mesh_2_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2434 == GlobalFiModInstNr[0]) || (2434 == GlobalFiModInstNr[1]) || (2434 == GlobalFiModInstNr[2]) || (2434 == GlobalFiModInstNr[3]))));
	Tile mesh_2_8(
		.clock(clock),
		.io_in_a_0(r_40_0),
		.io_in_b_0(b_130_0),
		.io_in_d_0(b_386_0),
		.io_in_control_0_dataflow(mesh_2_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_8_io_in_control_0_shift_b),
		.io_in_id_0(r_642_0),
		.io_in_last_0(r_898_0),
		.io_in_valid_0(r_386_0),
		.io_out_a_0(_mesh_2_8_io_out_a_0),
		.io_out_c_0(_mesh_2_8_io_out_c_0),
		.io_out_b_0(_mesh_2_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_8_io_out_id_0),
		.io_out_last_0(_mesh_2_8_io_out_last_0),
		.io_out_valid_0(_mesh_2_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2435 == GlobalFiModInstNr[0]) || (2435 == GlobalFiModInstNr[1]) || (2435 == GlobalFiModInstNr[2]) || (2435 == GlobalFiModInstNr[3]))));
	Tile mesh_2_9(
		.clock(clock),
		.io_in_a_0(r_41_0),
		.io_in_b_0(b_146_0),
		.io_in_d_0(b_402_0),
		.io_in_control_0_dataflow(mesh_2_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_9_io_in_control_0_shift_b),
		.io_in_id_0(r_658_0),
		.io_in_last_0(r_914_0),
		.io_in_valid_0(r_402_0),
		.io_out_a_0(_mesh_2_9_io_out_a_0),
		.io_out_c_0(_mesh_2_9_io_out_c_0),
		.io_out_b_0(_mesh_2_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_9_io_out_id_0),
		.io_out_last_0(_mesh_2_9_io_out_last_0),
		.io_out_valid_0(_mesh_2_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2436 == GlobalFiModInstNr[0]) || (2436 == GlobalFiModInstNr[1]) || (2436 == GlobalFiModInstNr[2]) || (2436 == GlobalFiModInstNr[3]))));
	Tile mesh_2_10(
		.clock(clock),
		.io_in_a_0(r_42_0),
		.io_in_b_0(b_162_0),
		.io_in_d_0(b_418_0),
		.io_in_control_0_dataflow(mesh_2_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_10_io_in_control_0_shift_b),
		.io_in_id_0(r_674_0),
		.io_in_last_0(r_930_0),
		.io_in_valid_0(r_418_0),
		.io_out_a_0(_mesh_2_10_io_out_a_0),
		.io_out_c_0(_mesh_2_10_io_out_c_0),
		.io_out_b_0(_mesh_2_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_10_io_out_id_0),
		.io_out_last_0(_mesh_2_10_io_out_last_0),
		.io_out_valid_0(_mesh_2_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2437 == GlobalFiModInstNr[0]) || (2437 == GlobalFiModInstNr[1]) || (2437 == GlobalFiModInstNr[2]) || (2437 == GlobalFiModInstNr[3]))));
	Tile mesh_2_11(
		.clock(clock),
		.io_in_a_0(r_43_0),
		.io_in_b_0(b_178_0),
		.io_in_d_0(b_434_0),
		.io_in_control_0_dataflow(mesh_2_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_11_io_in_control_0_shift_b),
		.io_in_id_0(r_690_0),
		.io_in_last_0(r_946_0),
		.io_in_valid_0(r_434_0),
		.io_out_a_0(_mesh_2_11_io_out_a_0),
		.io_out_c_0(_mesh_2_11_io_out_c_0),
		.io_out_b_0(_mesh_2_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_11_io_out_id_0),
		.io_out_last_0(_mesh_2_11_io_out_last_0),
		.io_out_valid_0(_mesh_2_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2438 == GlobalFiModInstNr[0]) || (2438 == GlobalFiModInstNr[1]) || (2438 == GlobalFiModInstNr[2]) || (2438 == GlobalFiModInstNr[3]))));
	Tile mesh_2_12(
		.clock(clock),
		.io_in_a_0(r_44_0),
		.io_in_b_0(b_194_0),
		.io_in_d_0(b_450_0),
		.io_in_control_0_dataflow(mesh_2_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_12_io_in_control_0_shift_b),
		.io_in_id_0(r_706_0),
		.io_in_last_0(r_962_0),
		.io_in_valid_0(r_450_0),
		.io_out_a_0(_mesh_2_12_io_out_a_0),
		.io_out_c_0(_mesh_2_12_io_out_c_0),
		.io_out_b_0(_mesh_2_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_12_io_out_id_0),
		.io_out_last_0(_mesh_2_12_io_out_last_0),
		.io_out_valid_0(_mesh_2_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2439 == GlobalFiModInstNr[0]) || (2439 == GlobalFiModInstNr[1]) || (2439 == GlobalFiModInstNr[2]) || (2439 == GlobalFiModInstNr[3]))));
	Tile mesh_2_13(
		.clock(clock),
		.io_in_a_0(r_45_0),
		.io_in_b_0(b_210_0),
		.io_in_d_0(b_466_0),
		.io_in_control_0_dataflow(mesh_2_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_13_io_in_control_0_shift_b),
		.io_in_id_0(r_722_0),
		.io_in_last_0(r_978_0),
		.io_in_valid_0(r_466_0),
		.io_out_a_0(_mesh_2_13_io_out_a_0),
		.io_out_c_0(_mesh_2_13_io_out_c_0),
		.io_out_b_0(_mesh_2_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_13_io_out_id_0),
		.io_out_last_0(_mesh_2_13_io_out_last_0),
		.io_out_valid_0(_mesh_2_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2440 == GlobalFiModInstNr[0]) || (2440 == GlobalFiModInstNr[1]) || (2440 == GlobalFiModInstNr[2]) || (2440 == GlobalFiModInstNr[3]))));
	Tile mesh_2_14(
		.clock(clock),
		.io_in_a_0(r_46_0),
		.io_in_b_0(b_226_0),
		.io_in_d_0(b_482_0),
		.io_in_control_0_dataflow(mesh_2_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_14_io_in_control_0_shift_b),
		.io_in_id_0(r_738_0),
		.io_in_last_0(r_994_0),
		.io_in_valid_0(r_482_0),
		.io_out_a_0(_mesh_2_14_io_out_a_0),
		.io_out_c_0(_mesh_2_14_io_out_c_0),
		.io_out_b_0(_mesh_2_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_14_io_out_id_0),
		.io_out_last_0(_mesh_2_14_io_out_last_0),
		.io_out_valid_0(_mesh_2_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2441 == GlobalFiModInstNr[0]) || (2441 == GlobalFiModInstNr[1]) || (2441 == GlobalFiModInstNr[2]) || (2441 == GlobalFiModInstNr[3]))));
	Tile mesh_2_15(
		.clock(clock),
		.io_in_a_0(r_47_0),
		.io_in_b_0(b_242_0),
		.io_in_d_0(b_498_0),
		.io_in_control_0_dataflow(mesh_2_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_15_io_in_control_0_shift_b),
		.io_in_id_0(r_754_0),
		.io_in_last_0(r_1010_0),
		.io_in_valid_0(r_498_0),
		.io_out_a_0(_mesh_2_15_io_out_a_0),
		.io_out_c_0(_mesh_2_15_io_out_c_0),
		.io_out_b_0(_mesh_2_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_15_io_out_id_0),
		.io_out_last_0(_mesh_2_15_io_out_last_0),
		.io_out_valid_0(_mesh_2_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2442 == GlobalFiModInstNr[0]) || (2442 == GlobalFiModInstNr[1]) || (2442 == GlobalFiModInstNr[2]) || (2442 == GlobalFiModInstNr[3]))));
	Tile mesh_3_0(
		.clock(clock),
		.io_in_a_0(r_48_0),
		.io_in_b_0(b_3_0),
		.io_in_d_0(b_259_0),
		.io_in_control_0_dataflow(mesh_3_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_0_io_in_control_0_shift_b),
		.io_in_id_0(r_515_0),
		.io_in_last_0(r_771_0),
		.io_in_valid_0(r_259_0),
		.io_out_a_0(_mesh_3_0_io_out_a_0),
		.io_out_c_0(_mesh_3_0_io_out_c_0),
		.io_out_b_0(_mesh_3_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_0_io_out_id_0),
		.io_out_last_0(_mesh_3_0_io_out_last_0),
		.io_out_valid_0(_mesh_3_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2443 == GlobalFiModInstNr[0]) || (2443 == GlobalFiModInstNr[1]) || (2443 == GlobalFiModInstNr[2]) || (2443 == GlobalFiModInstNr[3]))));
	Tile mesh_3_1(
		.clock(clock),
		.io_in_a_0(r_49_0),
		.io_in_b_0(b_19_0),
		.io_in_d_0(b_275_0),
		.io_in_control_0_dataflow(mesh_3_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_1_io_in_control_0_shift_b),
		.io_in_id_0(r_531_0),
		.io_in_last_0(r_787_0),
		.io_in_valid_0(r_275_0),
		.io_out_a_0(_mesh_3_1_io_out_a_0),
		.io_out_c_0(_mesh_3_1_io_out_c_0),
		.io_out_b_0(_mesh_3_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_1_io_out_id_0),
		.io_out_last_0(_mesh_3_1_io_out_last_0),
		.io_out_valid_0(_mesh_3_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2444 == GlobalFiModInstNr[0]) || (2444 == GlobalFiModInstNr[1]) || (2444 == GlobalFiModInstNr[2]) || (2444 == GlobalFiModInstNr[3]))));
	Tile mesh_3_2(
		.clock(clock),
		.io_in_a_0(r_50_0),
		.io_in_b_0(b_35_0),
		.io_in_d_0(b_291_0),
		.io_in_control_0_dataflow(mesh_3_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_2_io_in_control_0_shift_b),
		.io_in_id_0(r_547_0),
		.io_in_last_0(r_803_0),
		.io_in_valid_0(r_291_0),
		.io_out_a_0(_mesh_3_2_io_out_a_0),
		.io_out_c_0(_mesh_3_2_io_out_c_0),
		.io_out_b_0(_mesh_3_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_2_io_out_id_0),
		.io_out_last_0(_mesh_3_2_io_out_last_0),
		.io_out_valid_0(_mesh_3_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2445 == GlobalFiModInstNr[0]) || (2445 == GlobalFiModInstNr[1]) || (2445 == GlobalFiModInstNr[2]) || (2445 == GlobalFiModInstNr[3]))));
	Tile mesh_3_3(
		.clock(clock),
		.io_in_a_0(r_51_0),
		.io_in_b_0(b_51_0),
		.io_in_d_0(b_307_0),
		.io_in_control_0_dataflow(mesh_3_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_3_io_in_control_0_shift_b),
		.io_in_id_0(r_563_0),
		.io_in_last_0(r_819_0),
		.io_in_valid_0(r_307_0),
		.io_out_a_0(_mesh_3_3_io_out_a_0),
		.io_out_c_0(_mesh_3_3_io_out_c_0),
		.io_out_b_0(_mesh_3_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_3_io_out_id_0),
		.io_out_last_0(_mesh_3_3_io_out_last_0),
		.io_out_valid_0(_mesh_3_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2446 == GlobalFiModInstNr[0]) || (2446 == GlobalFiModInstNr[1]) || (2446 == GlobalFiModInstNr[2]) || (2446 == GlobalFiModInstNr[3]))));
	Tile mesh_3_4(
		.clock(clock),
		.io_in_a_0(r_52_0),
		.io_in_b_0(b_67_0),
		.io_in_d_0(b_323_0),
		.io_in_control_0_dataflow(mesh_3_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_4_io_in_control_0_shift_b),
		.io_in_id_0(r_579_0),
		.io_in_last_0(r_835_0),
		.io_in_valid_0(r_323_0),
		.io_out_a_0(_mesh_3_4_io_out_a_0),
		.io_out_c_0(_mesh_3_4_io_out_c_0),
		.io_out_b_0(_mesh_3_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_4_io_out_id_0),
		.io_out_last_0(_mesh_3_4_io_out_last_0),
		.io_out_valid_0(_mesh_3_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2447 == GlobalFiModInstNr[0]) || (2447 == GlobalFiModInstNr[1]) || (2447 == GlobalFiModInstNr[2]) || (2447 == GlobalFiModInstNr[3]))));
	Tile mesh_3_5(
		.clock(clock),
		.io_in_a_0(r_53_0),
		.io_in_b_0(b_83_0),
		.io_in_d_0(b_339_0),
		.io_in_control_0_dataflow(mesh_3_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_5_io_in_control_0_shift_b),
		.io_in_id_0(r_595_0),
		.io_in_last_0(r_851_0),
		.io_in_valid_0(r_339_0),
		.io_out_a_0(_mesh_3_5_io_out_a_0),
		.io_out_c_0(_mesh_3_5_io_out_c_0),
		.io_out_b_0(_mesh_3_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_5_io_out_id_0),
		.io_out_last_0(_mesh_3_5_io_out_last_0),
		.io_out_valid_0(_mesh_3_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2448 == GlobalFiModInstNr[0]) || (2448 == GlobalFiModInstNr[1]) || (2448 == GlobalFiModInstNr[2]) || (2448 == GlobalFiModInstNr[3]))));
	Tile mesh_3_6(
		.clock(clock),
		.io_in_a_0(r_54_0),
		.io_in_b_0(b_99_0),
		.io_in_d_0(b_355_0),
		.io_in_control_0_dataflow(mesh_3_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_6_io_in_control_0_shift_b),
		.io_in_id_0(r_611_0),
		.io_in_last_0(r_867_0),
		.io_in_valid_0(r_355_0),
		.io_out_a_0(_mesh_3_6_io_out_a_0),
		.io_out_c_0(_mesh_3_6_io_out_c_0),
		.io_out_b_0(_mesh_3_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_6_io_out_id_0),
		.io_out_last_0(_mesh_3_6_io_out_last_0),
		.io_out_valid_0(_mesh_3_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2449 == GlobalFiModInstNr[0]) || (2449 == GlobalFiModInstNr[1]) || (2449 == GlobalFiModInstNr[2]) || (2449 == GlobalFiModInstNr[3]))));
	Tile mesh_3_7(
		.clock(clock),
		.io_in_a_0(r_55_0),
		.io_in_b_0(b_115_0),
		.io_in_d_0(b_371_0),
		.io_in_control_0_dataflow(mesh_3_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_7_io_in_control_0_shift_b),
		.io_in_id_0(r_627_0),
		.io_in_last_0(r_883_0),
		.io_in_valid_0(r_371_0),
		.io_out_a_0(_mesh_3_7_io_out_a_0),
		.io_out_c_0(_mesh_3_7_io_out_c_0),
		.io_out_b_0(_mesh_3_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_7_io_out_id_0),
		.io_out_last_0(_mesh_3_7_io_out_last_0),
		.io_out_valid_0(_mesh_3_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2450 == GlobalFiModInstNr[0]) || (2450 == GlobalFiModInstNr[1]) || (2450 == GlobalFiModInstNr[2]) || (2450 == GlobalFiModInstNr[3]))));
	Tile mesh_3_8(
		.clock(clock),
		.io_in_a_0(r_56_0),
		.io_in_b_0(b_131_0),
		.io_in_d_0(b_387_0),
		.io_in_control_0_dataflow(mesh_3_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_8_io_in_control_0_shift_b),
		.io_in_id_0(r_643_0),
		.io_in_last_0(r_899_0),
		.io_in_valid_0(r_387_0),
		.io_out_a_0(_mesh_3_8_io_out_a_0),
		.io_out_c_0(_mesh_3_8_io_out_c_0),
		.io_out_b_0(_mesh_3_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_8_io_out_id_0),
		.io_out_last_0(_mesh_3_8_io_out_last_0),
		.io_out_valid_0(_mesh_3_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2451 == GlobalFiModInstNr[0]) || (2451 == GlobalFiModInstNr[1]) || (2451 == GlobalFiModInstNr[2]) || (2451 == GlobalFiModInstNr[3]))));
	Tile mesh_3_9(
		.clock(clock),
		.io_in_a_0(r_57_0),
		.io_in_b_0(b_147_0),
		.io_in_d_0(b_403_0),
		.io_in_control_0_dataflow(mesh_3_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_9_io_in_control_0_shift_b),
		.io_in_id_0(r_659_0),
		.io_in_last_0(r_915_0),
		.io_in_valid_0(r_403_0),
		.io_out_a_0(_mesh_3_9_io_out_a_0),
		.io_out_c_0(_mesh_3_9_io_out_c_0),
		.io_out_b_0(_mesh_3_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_9_io_out_id_0),
		.io_out_last_0(_mesh_3_9_io_out_last_0),
		.io_out_valid_0(_mesh_3_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2452 == GlobalFiModInstNr[0]) || (2452 == GlobalFiModInstNr[1]) || (2452 == GlobalFiModInstNr[2]) || (2452 == GlobalFiModInstNr[3]))));
	Tile mesh_3_10(
		.clock(clock),
		.io_in_a_0(r_58_0),
		.io_in_b_0(b_163_0),
		.io_in_d_0(b_419_0),
		.io_in_control_0_dataflow(mesh_3_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_10_io_in_control_0_shift_b),
		.io_in_id_0(r_675_0),
		.io_in_last_0(r_931_0),
		.io_in_valid_0(r_419_0),
		.io_out_a_0(_mesh_3_10_io_out_a_0),
		.io_out_c_0(_mesh_3_10_io_out_c_0),
		.io_out_b_0(_mesh_3_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_10_io_out_id_0),
		.io_out_last_0(_mesh_3_10_io_out_last_0),
		.io_out_valid_0(_mesh_3_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2453 == GlobalFiModInstNr[0]) || (2453 == GlobalFiModInstNr[1]) || (2453 == GlobalFiModInstNr[2]) || (2453 == GlobalFiModInstNr[3]))));
	Tile mesh_3_11(
		.clock(clock),
		.io_in_a_0(r_59_0),
		.io_in_b_0(b_179_0),
		.io_in_d_0(b_435_0),
		.io_in_control_0_dataflow(mesh_3_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_11_io_in_control_0_shift_b),
		.io_in_id_0(r_691_0),
		.io_in_last_0(r_947_0),
		.io_in_valid_0(r_435_0),
		.io_out_a_0(_mesh_3_11_io_out_a_0),
		.io_out_c_0(_mesh_3_11_io_out_c_0),
		.io_out_b_0(_mesh_3_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_11_io_out_id_0),
		.io_out_last_0(_mesh_3_11_io_out_last_0),
		.io_out_valid_0(_mesh_3_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2454 == GlobalFiModInstNr[0]) || (2454 == GlobalFiModInstNr[1]) || (2454 == GlobalFiModInstNr[2]) || (2454 == GlobalFiModInstNr[3]))));
	Tile mesh_3_12(
		.clock(clock),
		.io_in_a_0(r_60_0),
		.io_in_b_0(b_195_0),
		.io_in_d_0(b_451_0),
		.io_in_control_0_dataflow(mesh_3_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_12_io_in_control_0_shift_b),
		.io_in_id_0(r_707_0),
		.io_in_last_0(r_963_0),
		.io_in_valid_0(r_451_0),
		.io_out_a_0(_mesh_3_12_io_out_a_0),
		.io_out_c_0(_mesh_3_12_io_out_c_0),
		.io_out_b_0(_mesh_3_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_12_io_out_id_0),
		.io_out_last_0(_mesh_3_12_io_out_last_0),
		.io_out_valid_0(_mesh_3_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2455 == GlobalFiModInstNr[0]) || (2455 == GlobalFiModInstNr[1]) || (2455 == GlobalFiModInstNr[2]) || (2455 == GlobalFiModInstNr[3]))));
	Tile mesh_3_13(
		.clock(clock),
		.io_in_a_0(r_61_0),
		.io_in_b_0(b_211_0),
		.io_in_d_0(b_467_0),
		.io_in_control_0_dataflow(mesh_3_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_13_io_in_control_0_shift_b),
		.io_in_id_0(r_723_0),
		.io_in_last_0(r_979_0),
		.io_in_valid_0(r_467_0),
		.io_out_a_0(_mesh_3_13_io_out_a_0),
		.io_out_c_0(_mesh_3_13_io_out_c_0),
		.io_out_b_0(_mesh_3_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_13_io_out_id_0),
		.io_out_last_0(_mesh_3_13_io_out_last_0),
		.io_out_valid_0(_mesh_3_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2456 == GlobalFiModInstNr[0]) || (2456 == GlobalFiModInstNr[1]) || (2456 == GlobalFiModInstNr[2]) || (2456 == GlobalFiModInstNr[3]))));
	Tile mesh_3_14(
		.clock(clock),
		.io_in_a_0(r_62_0),
		.io_in_b_0(b_227_0),
		.io_in_d_0(b_483_0),
		.io_in_control_0_dataflow(mesh_3_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_14_io_in_control_0_shift_b),
		.io_in_id_0(r_739_0),
		.io_in_last_0(r_995_0),
		.io_in_valid_0(r_483_0),
		.io_out_a_0(_mesh_3_14_io_out_a_0),
		.io_out_c_0(_mesh_3_14_io_out_c_0),
		.io_out_b_0(_mesh_3_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_14_io_out_id_0),
		.io_out_last_0(_mesh_3_14_io_out_last_0),
		.io_out_valid_0(_mesh_3_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2457 == GlobalFiModInstNr[0]) || (2457 == GlobalFiModInstNr[1]) || (2457 == GlobalFiModInstNr[2]) || (2457 == GlobalFiModInstNr[3]))));
	Tile mesh_3_15(
		.clock(clock),
		.io_in_a_0(r_63_0),
		.io_in_b_0(b_243_0),
		.io_in_d_0(b_499_0),
		.io_in_control_0_dataflow(mesh_3_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_15_io_in_control_0_shift_b),
		.io_in_id_0(r_755_0),
		.io_in_last_0(r_1011_0),
		.io_in_valid_0(r_499_0),
		.io_out_a_0(_mesh_3_15_io_out_a_0),
		.io_out_c_0(_mesh_3_15_io_out_c_0),
		.io_out_b_0(_mesh_3_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_15_io_out_id_0),
		.io_out_last_0(_mesh_3_15_io_out_last_0),
		.io_out_valid_0(_mesh_3_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2458 == GlobalFiModInstNr[0]) || (2458 == GlobalFiModInstNr[1]) || (2458 == GlobalFiModInstNr[2]) || (2458 == GlobalFiModInstNr[3]))));
	Tile mesh_4_0(
		.clock(clock),
		.io_in_a_0(r_64_0),
		.io_in_b_0(b_4_0),
		.io_in_d_0(b_260_0),
		.io_in_control_0_dataflow(mesh_4_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_0_io_in_control_0_shift_b),
		.io_in_id_0(r_516_0),
		.io_in_last_0(r_772_0),
		.io_in_valid_0(r_260_0),
		.io_out_a_0(_mesh_4_0_io_out_a_0),
		.io_out_c_0(_mesh_4_0_io_out_c_0),
		.io_out_b_0(_mesh_4_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_0_io_out_id_0),
		.io_out_last_0(_mesh_4_0_io_out_last_0),
		.io_out_valid_0(_mesh_4_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2459 == GlobalFiModInstNr[0]) || (2459 == GlobalFiModInstNr[1]) || (2459 == GlobalFiModInstNr[2]) || (2459 == GlobalFiModInstNr[3]))));
	Tile mesh_4_1(
		.clock(clock),
		.io_in_a_0(r_65_0),
		.io_in_b_0(b_20_0),
		.io_in_d_0(b_276_0),
		.io_in_control_0_dataflow(mesh_4_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_1_io_in_control_0_shift_b),
		.io_in_id_0(r_532_0),
		.io_in_last_0(r_788_0),
		.io_in_valid_0(r_276_0),
		.io_out_a_0(_mesh_4_1_io_out_a_0),
		.io_out_c_0(_mesh_4_1_io_out_c_0),
		.io_out_b_0(_mesh_4_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_1_io_out_id_0),
		.io_out_last_0(_mesh_4_1_io_out_last_0),
		.io_out_valid_0(_mesh_4_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2460 == GlobalFiModInstNr[0]) || (2460 == GlobalFiModInstNr[1]) || (2460 == GlobalFiModInstNr[2]) || (2460 == GlobalFiModInstNr[3]))));
	Tile mesh_4_2(
		.clock(clock),
		.io_in_a_0(r_66_0),
		.io_in_b_0(b_36_0),
		.io_in_d_0(b_292_0),
		.io_in_control_0_dataflow(mesh_4_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_2_io_in_control_0_shift_b),
		.io_in_id_0(r_548_0),
		.io_in_last_0(r_804_0),
		.io_in_valid_0(r_292_0),
		.io_out_a_0(_mesh_4_2_io_out_a_0),
		.io_out_c_0(_mesh_4_2_io_out_c_0),
		.io_out_b_0(_mesh_4_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_2_io_out_id_0),
		.io_out_last_0(_mesh_4_2_io_out_last_0),
		.io_out_valid_0(_mesh_4_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2461 == GlobalFiModInstNr[0]) || (2461 == GlobalFiModInstNr[1]) || (2461 == GlobalFiModInstNr[2]) || (2461 == GlobalFiModInstNr[3]))));
	Tile mesh_4_3(
		.clock(clock),
		.io_in_a_0(r_67_0),
		.io_in_b_0(b_52_0),
		.io_in_d_0(b_308_0),
		.io_in_control_0_dataflow(mesh_4_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_3_io_in_control_0_shift_b),
		.io_in_id_0(r_564_0),
		.io_in_last_0(r_820_0),
		.io_in_valid_0(r_308_0),
		.io_out_a_0(_mesh_4_3_io_out_a_0),
		.io_out_c_0(_mesh_4_3_io_out_c_0),
		.io_out_b_0(_mesh_4_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_3_io_out_id_0),
		.io_out_last_0(_mesh_4_3_io_out_last_0),
		.io_out_valid_0(_mesh_4_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2462 == GlobalFiModInstNr[0]) || (2462 == GlobalFiModInstNr[1]) || (2462 == GlobalFiModInstNr[2]) || (2462 == GlobalFiModInstNr[3]))));
	Tile mesh_4_4(
		.clock(clock),
		.io_in_a_0(r_68_0),
		.io_in_b_0(b_68_0),
		.io_in_d_0(b_324_0),
		.io_in_control_0_dataflow(mesh_4_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_4_io_in_control_0_shift_b),
		.io_in_id_0(r_580_0),
		.io_in_last_0(r_836_0),
		.io_in_valid_0(r_324_0),
		.io_out_a_0(_mesh_4_4_io_out_a_0),
		.io_out_c_0(_mesh_4_4_io_out_c_0),
		.io_out_b_0(_mesh_4_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_4_io_out_id_0),
		.io_out_last_0(_mesh_4_4_io_out_last_0),
		.io_out_valid_0(_mesh_4_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2463 == GlobalFiModInstNr[0]) || (2463 == GlobalFiModInstNr[1]) || (2463 == GlobalFiModInstNr[2]) || (2463 == GlobalFiModInstNr[3]))));
	Tile mesh_4_5(
		.clock(clock),
		.io_in_a_0(r_69_0),
		.io_in_b_0(b_84_0),
		.io_in_d_0(b_340_0),
		.io_in_control_0_dataflow(mesh_4_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_5_io_in_control_0_shift_b),
		.io_in_id_0(r_596_0),
		.io_in_last_0(r_852_0),
		.io_in_valid_0(r_340_0),
		.io_out_a_0(_mesh_4_5_io_out_a_0),
		.io_out_c_0(_mesh_4_5_io_out_c_0),
		.io_out_b_0(_mesh_4_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_5_io_out_id_0),
		.io_out_last_0(_mesh_4_5_io_out_last_0),
		.io_out_valid_0(_mesh_4_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2464 == GlobalFiModInstNr[0]) || (2464 == GlobalFiModInstNr[1]) || (2464 == GlobalFiModInstNr[2]) || (2464 == GlobalFiModInstNr[3]))));
	Tile mesh_4_6(
		.clock(clock),
		.io_in_a_0(r_70_0),
		.io_in_b_0(b_100_0),
		.io_in_d_0(b_356_0),
		.io_in_control_0_dataflow(mesh_4_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_6_io_in_control_0_shift_b),
		.io_in_id_0(r_612_0),
		.io_in_last_0(r_868_0),
		.io_in_valid_0(r_356_0),
		.io_out_a_0(_mesh_4_6_io_out_a_0),
		.io_out_c_0(_mesh_4_6_io_out_c_0),
		.io_out_b_0(_mesh_4_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_6_io_out_id_0),
		.io_out_last_0(_mesh_4_6_io_out_last_0),
		.io_out_valid_0(_mesh_4_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2465 == GlobalFiModInstNr[0]) || (2465 == GlobalFiModInstNr[1]) || (2465 == GlobalFiModInstNr[2]) || (2465 == GlobalFiModInstNr[3]))));
	Tile mesh_4_7(
		.clock(clock),
		.io_in_a_0(r_71_0),
		.io_in_b_0(b_116_0),
		.io_in_d_0(b_372_0),
		.io_in_control_0_dataflow(mesh_4_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_7_io_in_control_0_shift_b),
		.io_in_id_0(r_628_0),
		.io_in_last_0(r_884_0),
		.io_in_valid_0(r_372_0),
		.io_out_a_0(_mesh_4_7_io_out_a_0),
		.io_out_c_0(_mesh_4_7_io_out_c_0),
		.io_out_b_0(_mesh_4_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_7_io_out_id_0),
		.io_out_last_0(_mesh_4_7_io_out_last_0),
		.io_out_valid_0(_mesh_4_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2466 == GlobalFiModInstNr[0]) || (2466 == GlobalFiModInstNr[1]) || (2466 == GlobalFiModInstNr[2]) || (2466 == GlobalFiModInstNr[3]))));
	Tile mesh_4_8(
		.clock(clock),
		.io_in_a_0(r_72_0),
		.io_in_b_0(b_132_0),
		.io_in_d_0(b_388_0),
		.io_in_control_0_dataflow(mesh_4_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_8_io_in_control_0_shift_b),
		.io_in_id_0(r_644_0),
		.io_in_last_0(r_900_0),
		.io_in_valid_0(r_388_0),
		.io_out_a_0(_mesh_4_8_io_out_a_0),
		.io_out_c_0(_mesh_4_8_io_out_c_0),
		.io_out_b_0(_mesh_4_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_8_io_out_id_0),
		.io_out_last_0(_mesh_4_8_io_out_last_0),
		.io_out_valid_0(_mesh_4_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2467 == GlobalFiModInstNr[0]) || (2467 == GlobalFiModInstNr[1]) || (2467 == GlobalFiModInstNr[2]) || (2467 == GlobalFiModInstNr[3]))));
	Tile mesh_4_9(
		.clock(clock),
		.io_in_a_0(r_73_0),
		.io_in_b_0(b_148_0),
		.io_in_d_0(b_404_0),
		.io_in_control_0_dataflow(mesh_4_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_9_io_in_control_0_shift_b),
		.io_in_id_0(r_660_0),
		.io_in_last_0(r_916_0),
		.io_in_valid_0(r_404_0),
		.io_out_a_0(_mesh_4_9_io_out_a_0),
		.io_out_c_0(_mesh_4_9_io_out_c_0),
		.io_out_b_0(_mesh_4_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_9_io_out_id_0),
		.io_out_last_0(_mesh_4_9_io_out_last_0),
		.io_out_valid_0(_mesh_4_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2468 == GlobalFiModInstNr[0]) || (2468 == GlobalFiModInstNr[1]) || (2468 == GlobalFiModInstNr[2]) || (2468 == GlobalFiModInstNr[3]))));
	Tile mesh_4_10(
		.clock(clock),
		.io_in_a_0(r_74_0),
		.io_in_b_0(b_164_0),
		.io_in_d_0(b_420_0),
		.io_in_control_0_dataflow(mesh_4_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_10_io_in_control_0_shift_b),
		.io_in_id_0(r_676_0),
		.io_in_last_0(r_932_0),
		.io_in_valid_0(r_420_0),
		.io_out_a_0(_mesh_4_10_io_out_a_0),
		.io_out_c_0(_mesh_4_10_io_out_c_0),
		.io_out_b_0(_mesh_4_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_10_io_out_id_0),
		.io_out_last_0(_mesh_4_10_io_out_last_0),
		.io_out_valid_0(_mesh_4_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2469 == GlobalFiModInstNr[0]) || (2469 == GlobalFiModInstNr[1]) || (2469 == GlobalFiModInstNr[2]) || (2469 == GlobalFiModInstNr[3]))));
	Tile mesh_4_11(
		.clock(clock),
		.io_in_a_0(r_75_0),
		.io_in_b_0(b_180_0),
		.io_in_d_0(b_436_0),
		.io_in_control_0_dataflow(mesh_4_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_11_io_in_control_0_shift_b),
		.io_in_id_0(r_692_0),
		.io_in_last_0(r_948_0),
		.io_in_valid_0(r_436_0),
		.io_out_a_0(_mesh_4_11_io_out_a_0),
		.io_out_c_0(_mesh_4_11_io_out_c_0),
		.io_out_b_0(_mesh_4_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_11_io_out_id_0),
		.io_out_last_0(_mesh_4_11_io_out_last_0),
		.io_out_valid_0(_mesh_4_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2470 == GlobalFiModInstNr[0]) || (2470 == GlobalFiModInstNr[1]) || (2470 == GlobalFiModInstNr[2]) || (2470 == GlobalFiModInstNr[3]))));
	Tile mesh_4_12(
		.clock(clock),
		.io_in_a_0(r_76_0),
		.io_in_b_0(b_196_0),
		.io_in_d_0(b_452_0),
		.io_in_control_0_dataflow(mesh_4_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_12_io_in_control_0_shift_b),
		.io_in_id_0(r_708_0),
		.io_in_last_0(r_964_0),
		.io_in_valid_0(r_452_0),
		.io_out_a_0(_mesh_4_12_io_out_a_0),
		.io_out_c_0(_mesh_4_12_io_out_c_0),
		.io_out_b_0(_mesh_4_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_12_io_out_id_0),
		.io_out_last_0(_mesh_4_12_io_out_last_0),
		.io_out_valid_0(_mesh_4_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2471 == GlobalFiModInstNr[0]) || (2471 == GlobalFiModInstNr[1]) || (2471 == GlobalFiModInstNr[2]) || (2471 == GlobalFiModInstNr[3]))));
	Tile mesh_4_13(
		.clock(clock),
		.io_in_a_0(r_77_0),
		.io_in_b_0(b_212_0),
		.io_in_d_0(b_468_0),
		.io_in_control_0_dataflow(mesh_4_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_13_io_in_control_0_shift_b),
		.io_in_id_0(r_724_0),
		.io_in_last_0(r_980_0),
		.io_in_valid_0(r_468_0),
		.io_out_a_0(_mesh_4_13_io_out_a_0),
		.io_out_c_0(_mesh_4_13_io_out_c_0),
		.io_out_b_0(_mesh_4_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_13_io_out_id_0),
		.io_out_last_0(_mesh_4_13_io_out_last_0),
		.io_out_valid_0(_mesh_4_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2472 == GlobalFiModInstNr[0]) || (2472 == GlobalFiModInstNr[1]) || (2472 == GlobalFiModInstNr[2]) || (2472 == GlobalFiModInstNr[3]))));
	Tile mesh_4_14(
		.clock(clock),
		.io_in_a_0(r_78_0),
		.io_in_b_0(b_228_0),
		.io_in_d_0(b_484_0),
		.io_in_control_0_dataflow(mesh_4_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_14_io_in_control_0_shift_b),
		.io_in_id_0(r_740_0),
		.io_in_last_0(r_996_0),
		.io_in_valid_0(r_484_0),
		.io_out_a_0(_mesh_4_14_io_out_a_0),
		.io_out_c_0(_mesh_4_14_io_out_c_0),
		.io_out_b_0(_mesh_4_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_14_io_out_id_0),
		.io_out_last_0(_mesh_4_14_io_out_last_0),
		.io_out_valid_0(_mesh_4_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2473 == GlobalFiModInstNr[0]) || (2473 == GlobalFiModInstNr[1]) || (2473 == GlobalFiModInstNr[2]) || (2473 == GlobalFiModInstNr[3]))));
	Tile mesh_4_15(
		.clock(clock),
		.io_in_a_0(r_79_0),
		.io_in_b_0(b_244_0),
		.io_in_d_0(b_500_0),
		.io_in_control_0_dataflow(mesh_4_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_15_io_in_control_0_shift_b),
		.io_in_id_0(r_756_0),
		.io_in_last_0(r_1012_0),
		.io_in_valid_0(r_500_0),
		.io_out_a_0(_mesh_4_15_io_out_a_0),
		.io_out_c_0(_mesh_4_15_io_out_c_0),
		.io_out_b_0(_mesh_4_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_15_io_out_id_0),
		.io_out_last_0(_mesh_4_15_io_out_last_0),
		.io_out_valid_0(_mesh_4_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2474 == GlobalFiModInstNr[0]) || (2474 == GlobalFiModInstNr[1]) || (2474 == GlobalFiModInstNr[2]) || (2474 == GlobalFiModInstNr[3]))));
	Tile mesh_5_0(
		.clock(clock),
		.io_in_a_0(r_80_0),
		.io_in_b_0(b_5_0),
		.io_in_d_0(b_261_0),
		.io_in_control_0_dataflow(mesh_5_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_0_io_in_control_0_shift_b),
		.io_in_id_0(r_517_0),
		.io_in_last_0(r_773_0),
		.io_in_valid_0(r_261_0),
		.io_out_a_0(_mesh_5_0_io_out_a_0),
		.io_out_c_0(_mesh_5_0_io_out_c_0),
		.io_out_b_0(_mesh_5_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_0_io_out_id_0),
		.io_out_last_0(_mesh_5_0_io_out_last_0),
		.io_out_valid_0(_mesh_5_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2475 == GlobalFiModInstNr[0]) || (2475 == GlobalFiModInstNr[1]) || (2475 == GlobalFiModInstNr[2]) || (2475 == GlobalFiModInstNr[3]))));
	Tile mesh_5_1(
		.clock(clock),
		.io_in_a_0(r_81_0),
		.io_in_b_0(b_21_0),
		.io_in_d_0(b_277_0),
		.io_in_control_0_dataflow(mesh_5_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_1_io_in_control_0_shift_b),
		.io_in_id_0(r_533_0),
		.io_in_last_0(r_789_0),
		.io_in_valid_0(r_277_0),
		.io_out_a_0(_mesh_5_1_io_out_a_0),
		.io_out_c_0(_mesh_5_1_io_out_c_0),
		.io_out_b_0(_mesh_5_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_1_io_out_id_0),
		.io_out_last_0(_mesh_5_1_io_out_last_0),
		.io_out_valid_0(_mesh_5_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2476 == GlobalFiModInstNr[0]) || (2476 == GlobalFiModInstNr[1]) || (2476 == GlobalFiModInstNr[2]) || (2476 == GlobalFiModInstNr[3]))));
	Tile mesh_5_2(
		.clock(clock),
		.io_in_a_0(r_82_0),
		.io_in_b_0(b_37_0),
		.io_in_d_0(b_293_0),
		.io_in_control_0_dataflow(mesh_5_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_2_io_in_control_0_shift_b),
		.io_in_id_0(r_549_0),
		.io_in_last_0(r_805_0),
		.io_in_valid_0(r_293_0),
		.io_out_a_0(_mesh_5_2_io_out_a_0),
		.io_out_c_0(_mesh_5_2_io_out_c_0),
		.io_out_b_0(_mesh_5_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_2_io_out_id_0),
		.io_out_last_0(_mesh_5_2_io_out_last_0),
		.io_out_valid_0(_mesh_5_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2477 == GlobalFiModInstNr[0]) || (2477 == GlobalFiModInstNr[1]) || (2477 == GlobalFiModInstNr[2]) || (2477 == GlobalFiModInstNr[3]))));
	Tile mesh_5_3(
		.clock(clock),
		.io_in_a_0(r_83_0),
		.io_in_b_0(b_53_0),
		.io_in_d_0(b_309_0),
		.io_in_control_0_dataflow(mesh_5_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_3_io_in_control_0_shift_b),
		.io_in_id_0(r_565_0),
		.io_in_last_0(r_821_0),
		.io_in_valid_0(r_309_0),
		.io_out_a_0(_mesh_5_3_io_out_a_0),
		.io_out_c_0(_mesh_5_3_io_out_c_0),
		.io_out_b_0(_mesh_5_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_3_io_out_id_0),
		.io_out_last_0(_mesh_5_3_io_out_last_0),
		.io_out_valid_0(_mesh_5_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2478 == GlobalFiModInstNr[0]) || (2478 == GlobalFiModInstNr[1]) || (2478 == GlobalFiModInstNr[2]) || (2478 == GlobalFiModInstNr[3]))));
	Tile mesh_5_4(
		.clock(clock),
		.io_in_a_0(r_84_0),
		.io_in_b_0(b_69_0),
		.io_in_d_0(b_325_0),
		.io_in_control_0_dataflow(mesh_5_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_4_io_in_control_0_shift_b),
		.io_in_id_0(r_581_0),
		.io_in_last_0(r_837_0),
		.io_in_valid_0(r_325_0),
		.io_out_a_0(_mesh_5_4_io_out_a_0),
		.io_out_c_0(_mesh_5_4_io_out_c_0),
		.io_out_b_0(_mesh_5_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_4_io_out_id_0),
		.io_out_last_0(_mesh_5_4_io_out_last_0),
		.io_out_valid_0(_mesh_5_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2479 == GlobalFiModInstNr[0]) || (2479 == GlobalFiModInstNr[1]) || (2479 == GlobalFiModInstNr[2]) || (2479 == GlobalFiModInstNr[3]))));
	Tile mesh_5_5(
		.clock(clock),
		.io_in_a_0(r_85_0),
		.io_in_b_0(b_85_0),
		.io_in_d_0(b_341_0),
		.io_in_control_0_dataflow(mesh_5_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_5_io_in_control_0_shift_b),
		.io_in_id_0(r_597_0),
		.io_in_last_0(r_853_0),
		.io_in_valid_0(r_341_0),
		.io_out_a_0(_mesh_5_5_io_out_a_0),
		.io_out_c_0(_mesh_5_5_io_out_c_0),
		.io_out_b_0(_mesh_5_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_5_io_out_id_0),
		.io_out_last_0(_mesh_5_5_io_out_last_0),
		.io_out_valid_0(_mesh_5_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2480 == GlobalFiModInstNr[0]) || (2480 == GlobalFiModInstNr[1]) || (2480 == GlobalFiModInstNr[2]) || (2480 == GlobalFiModInstNr[3]))));
	Tile mesh_5_6(
		.clock(clock),
		.io_in_a_0(r_86_0),
		.io_in_b_0(b_101_0),
		.io_in_d_0(b_357_0),
		.io_in_control_0_dataflow(mesh_5_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_6_io_in_control_0_shift_b),
		.io_in_id_0(r_613_0),
		.io_in_last_0(r_869_0),
		.io_in_valid_0(r_357_0),
		.io_out_a_0(_mesh_5_6_io_out_a_0),
		.io_out_c_0(_mesh_5_6_io_out_c_0),
		.io_out_b_0(_mesh_5_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_6_io_out_id_0),
		.io_out_last_0(_mesh_5_6_io_out_last_0),
		.io_out_valid_0(_mesh_5_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2481 == GlobalFiModInstNr[0]) || (2481 == GlobalFiModInstNr[1]) || (2481 == GlobalFiModInstNr[2]) || (2481 == GlobalFiModInstNr[3]))));
	Tile mesh_5_7(
		.clock(clock),
		.io_in_a_0(r_87_0),
		.io_in_b_0(b_117_0),
		.io_in_d_0(b_373_0),
		.io_in_control_0_dataflow(mesh_5_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_7_io_in_control_0_shift_b),
		.io_in_id_0(r_629_0),
		.io_in_last_0(r_885_0),
		.io_in_valid_0(r_373_0),
		.io_out_a_0(_mesh_5_7_io_out_a_0),
		.io_out_c_0(_mesh_5_7_io_out_c_0),
		.io_out_b_0(_mesh_5_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_7_io_out_id_0),
		.io_out_last_0(_mesh_5_7_io_out_last_0),
		.io_out_valid_0(_mesh_5_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2482 == GlobalFiModInstNr[0]) || (2482 == GlobalFiModInstNr[1]) || (2482 == GlobalFiModInstNr[2]) || (2482 == GlobalFiModInstNr[3]))));
	Tile mesh_5_8(
		.clock(clock),
		.io_in_a_0(r_88_0),
		.io_in_b_0(b_133_0),
		.io_in_d_0(b_389_0),
		.io_in_control_0_dataflow(mesh_5_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_8_io_in_control_0_shift_b),
		.io_in_id_0(r_645_0),
		.io_in_last_0(r_901_0),
		.io_in_valid_0(r_389_0),
		.io_out_a_0(_mesh_5_8_io_out_a_0),
		.io_out_c_0(_mesh_5_8_io_out_c_0),
		.io_out_b_0(_mesh_5_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_8_io_out_id_0),
		.io_out_last_0(_mesh_5_8_io_out_last_0),
		.io_out_valid_0(_mesh_5_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2483 == GlobalFiModInstNr[0]) || (2483 == GlobalFiModInstNr[1]) || (2483 == GlobalFiModInstNr[2]) || (2483 == GlobalFiModInstNr[3]))));
	Tile mesh_5_9(
		.clock(clock),
		.io_in_a_0(r_89_0),
		.io_in_b_0(b_149_0),
		.io_in_d_0(b_405_0),
		.io_in_control_0_dataflow(mesh_5_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_9_io_in_control_0_shift_b),
		.io_in_id_0(r_661_0),
		.io_in_last_0(r_917_0),
		.io_in_valid_0(r_405_0),
		.io_out_a_0(_mesh_5_9_io_out_a_0),
		.io_out_c_0(_mesh_5_9_io_out_c_0),
		.io_out_b_0(_mesh_5_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_9_io_out_id_0),
		.io_out_last_0(_mesh_5_9_io_out_last_0),
		.io_out_valid_0(_mesh_5_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2484 == GlobalFiModInstNr[0]) || (2484 == GlobalFiModInstNr[1]) || (2484 == GlobalFiModInstNr[2]) || (2484 == GlobalFiModInstNr[3]))));
	Tile mesh_5_10(
		.clock(clock),
		.io_in_a_0(r_90_0),
		.io_in_b_0(b_165_0),
		.io_in_d_0(b_421_0),
		.io_in_control_0_dataflow(mesh_5_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_10_io_in_control_0_shift_b),
		.io_in_id_0(r_677_0),
		.io_in_last_0(r_933_0),
		.io_in_valid_0(r_421_0),
		.io_out_a_0(_mesh_5_10_io_out_a_0),
		.io_out_c_0(_mesh_5_10_io_out_c_0),
		.io_out_b_0(_mesh_5_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_10_io_out_id_0),
		.io_out_last_0(_mesh_5_10_io_out_last_0),
		.io_out_valid_0(_mesh_5_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2485 == GlobalFiModInstNr[0]) || (2485 == GlobalFiModInstNr[1]) || (2485 == GlobalFiModInstNr[2]) || (2485 == GlobalFiModInstNr[3]))));
	Tile mesh_5_11(
		.clock(clock),
		.io_in_a_0(r_91_0),
		.io_in_b_0(b_181_0),
		.io_in_d_0(b_437_0),
		.io_in_control_0_dataflow(mesh_5_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_11_io_in_control_0_shift_b),
		.io_in_id_0(r_693_0),
		.io_in_last_0(r_949_0),
		.io_in_valid_0(r_437_0),
		.io_out_a_0(_mesh_5_11_io_out_a_0),
		.io_out_c_0(_mesh_5_11_io_out_c_0),
		.io_out_b_0(_mesh_5_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_11_io_out_id_0),
		.io_out_last_0(_mesh_5_11_io_out_last_0),
		.io_out_valid_0(_mesh_5_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2486 == GlobalFiModInstNr[0]) || (2486 == GlobalFiModInstNr[1]) || (2486 == GlobalFiModInstNr[2]) || (2486 == GlobalFiModInstNr[3]))));
	Tile mesh_5_12(
		.clock(clock),
		.io_in_a_0(r_92_0),
		.io_in_b_0(b_197_0),
		.io_in_d_0(b_453_0),
		.io_in_control_0_dataflow(mesh_5_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_12_io_in_control_0_shift_b),
		.io_in_id_0(r_709_0),
		.io_in_last_0(r_965_0),
		.io_in_valid_0(r_453_0),
		.io_out_a_0(_mesh_5_12_io_out_a_0),
		.io_out_c_0(_mesh_5_12_io_out_c_0),
		.io_out_b_0(_mesh_5_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_12_io_out_id_0),
		.io_out_last_0(_mesh_5_12_io_out_last_0),
		.io_out_valid_0(_mesh_5_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2487 == GlobalFiModInstNr[0]) || (2487 == GlobalFiModInstNr[1]) || (2487 == GlobalFiModInstNr[2]) || (2487 == GlobalFiModInstNr[3]))));
	Tile mesh_5_13(
		.clock(clock),
		.io_in_a_0(r_93_0),
		.io_in_b_0(b_213_0),
		.io_in_d_0(b_469_0),
		.io_in_control_0_dataflow(mesh_5_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_13_io_in_control_0_shift_b),
		.io_in_id_0(r_725_0),
		.io_in_last_0(r_981_0),
		.io_in_valid_0(r_469_0),
		.io_out_a_0(_mesh_5_13_io_out_a_0),
		.io_out_c_0(_mesh_5_13_io_out_c_0),
		.io_out_b_0(_mesh_5_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_13_io_out_id_0),
		.io_out_last_0(_mesh_5_13_io_out_last_0),
		.io_out_valid_0(_mesh_5_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2488 == GlobalFiModInstNr[0]) || (2488 == GlobalFiModInstNr[1]) || (2488 == GlobalFiModInstNr[2]) || (2488 == GlobalFiModInstNr[3]))));
	Tile mesh_5_14(
		.clock(clock),
		.io_in_a_0(r_94_0),
		.io_in_b_0(b_229_0),
		.io_in_d_0(b_485_0),
		.io_in_control_0_dataflow(mesh_5_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_14_io_in_control_0_shift_b),
		.io_in_id_0(r_741_0),
		.io_in_last_0(r_997_0),
		.io_in_valid_0(r_485_0),
		.io_out_a_0(_mesh_5_14_io_out_a_0),
		.io_out_c_0(_mesh_5_14_io_out_c_0),
		.io_out_b_0(_mesh_5_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_14_io_out_id_0),
		.io_out_last_0(_mesh_5_14_io_out_last_0),
		.io_out_valid_0(_mesh_5_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2489 == GlobalFiModInstNr[0]) || (2489 == GlobalFiModInstNr[1]) || (2489 == GlobalFiModInstNr[2]) || (2489 == GlobalFiModInstNr[3]))));
	Tile mesh_5_15(
		.clock(clock),
		.io_in_a_0(r_95_0),
		.io_in_b_0(b_245_0),
		.io_in_d_0(b_501_0),
		.io_in_control_0_dataflow(mesh_5_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_15_io_in_control_0_shift_b),
		.io_in_id_0(r_757_0),
		.io_in_last_0(r_1013_0),
		.io_in_valid_0(r_501_0),
		.io_out_a_0(_mesh_5_15_io_out_a_0),
		.io_out_c_0(_mesh_5_15_io_out_c_0),
		.io_out_b_0(_mesh_5_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_15_io_out_id_0),
		.io_out_last_0(_mesh_5_15_io_out_last_0),
		.io_out_valid_0(_mesh_5_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2490 == GlobalFiModInstNr[0]) || (2490 == GlobalFiModInstNr[1]) || (2490 == GlobalFiModInstNr[2]) || (2490 == GlobalFiModInstNr[3]))));
	Tile mesh_6_0(
		.clock(clock),
		.io_in_a_0(r_96_0),
		.io_in_b_0(b_6_0),
		.io_in_d_0(b_262_0),
		.io_in_control_0_dataflow(mesh_6_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_0_io_in_control_0_shift_b),
		.io_in_id_0(r_518_0),
		.io_in_last_0(r_774_0),
		.io_in_valid_0(r_262_0),
		.io_out_a_0(_mesh_6_0_io_out_a_0),
		.io_out_c_0(_mesh_6_0_io_out_c_0),
		.io_out_b_0(_mesh_6_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_0_io_out_id_0),
		.io_out_last_0(_mesh_6_0_io_out_last_0),
		.io_out_valid_0(_mesh_6_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2491 == GlobalFiModInstNr[0]) || (2491 == GlobalFiModInstNr[1]) || (2491 == GlobalFiModInstNr[2]) || (2491 == GlobalFiModInstNr[3]))));
	Tile mesh_6_1(
		.clock(clock),
		.io_in_a_0(r_97_0),
		.io_in_b_0(b_22_0),
		.io_in_d_0(b_278_0),
		.io_in_control_0_dataflow(mesh_6_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_1_io_in_control_0_shift_b),
		.io_in_id_0(r_534_0),
		.io_in_last_0(r_790_0),
		.io_in_valid_0(r_278_0),
		.io_out_a_0(_mesh_6_1_io_out_a_0),
		.io_out_c_0(_mesh_6_1_io_out_c_0),
		.io_out_b_0(_mesh_6_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_1_io_out_id_0),
		.io_out_last_0(_mesh_6_1_io_out_last_0),
		.io_out_valid_0(_mesh_6_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2492 == GlobalFiModInstNr[0]) || (2492 == GlobalFiModInstNr[1]) || (2492 == GlobalFiModInstNr[2]) || (2492 == GlobalFiModInstNr[3]))));
	Tile mesh_6_2(
		.clock(clock),
		.io_in_a_0(r_98_0),
		.io_in_b_0(b_38_0),
		.io_in_d_0(b_294_0),
		.io_in_control_0_dataflow(mesh_6_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_2_io_in_control_0_shift_b),
		.io_in_id_0(r_550_0),
		.io_in_last_0(r_806_0),
		.io_in_valid_0(r_294_0),
		.io_out_a_0(_mesh_6_2_io_out_a_0),
		.io_out_c_0(_mesh_6_2_io_out_c_0),
		.io_out_b_0(_mesh_6_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_2_io_out_id_0),
		.io_out_last_0(_mesh_6_2_io_out_last_0),
		.io_out_valid_0(_mesh_6_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2493 == GlobalFiModInstNr[0]) || (2493 == GlobalFiModInstNr[1]) || (2493 == GlobalFiModInstNr[2]) || (2493 == GlobalFiModInstNr[3]))));
	Tile mesh_6_3(
		.clock(clock),
		.io_in_a_0(r_99_0),
		.io_in_b_0(b_54_0),
		.io_in_d_0(b_310_0),
		.io_in_control_0_dataflow(mesh_6_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_3_io_in_control_0_shift_b),
		.io_in_id_0(r_566_0),
		.io_in_last_0(r_822_0),
		.io_in_valid_0(r_310_0),
		.io_out_a_0(_mesh_6_3_io_out_a_0),
		.io_out_c_0(_mesh_6_3_io_out_c_0),
		.io_out_b_0(_mesh_6_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_3_io_out_id_0),
		.io_out_last_0(_mesh_6_3_io_out_last_0),
		.io_out_valid_0(_mesh_6_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2494 == GlobalFiModInstNr[0]) || (2494 == GlobalFiModInstNr[1]) || (2494 == GlobalFiModInstNr[2]) || (2494 == GlobalFiModInstNr[3]))));
	Tile mesh_6_4(
		.clock(clock),
		.io_in_a_0(r_100_0),
		.io_in_b_0(b_70_0),
		.io_in_d_0(b_326_0),
		.io_in_control_0_dataflow(mesh_6_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_4_io_in_control_0_shift_b),
		.io_in_id_0(r_582_0),
		.io_in_last_0(r_838_0),
		.io_in_valid_0(r_326_0),
		.io_out_a_0(_mesh_6_4_io_out_a_0),
		.io_out_c_0(_mesh_6_4_io_out_c_0),
		.io_out_b_0(_mesh_6_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_4_io_out_id_0),
		.io_out_last_0(_mesh_6_4_io_out_last_0),
		.io_out_valid_0(_mesh_6_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2495 == GlobalFiModInstNr[0]) || (2495 == GlobalFiModInstNr[1]) || (2495 == GlobalFiModInstNr[2]) || (2495 == GlobalFiModInstNr[3]))));
	Tile mesh_6_5(
		.clock(clock),
		.io_in_a_0(r_101_0),
		.io_in_b_0(b_86_0),
		.io_in_d_0(b_342_0),
		.io_in_control_0_dataflow(mesh_6_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_5_io_in_control_0_shift_b),
		.io_in_id_0(r_598_0),
		.io_in_last_0(r_854_0),
		.io_in_valid_0(r_342_0),
		.io_out_a_0(_mesh_6_5_io_out_a_0),
		.io_out_c_0(_mesh_6_5_io_out_c_0),
		.io_out_b_0(_mesh_6_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_5_io_out_id_0),
		.io_out_last_0(_mesh_6_5_io_out_last_0),
		.io_out_valid_0(_mesh_6_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2496 == GlobalFiModInstNr[0]) || (2496 == GlobalFiModInstNr[1]) || (2496 == GlobalFiModInstNr[2]) || (2496 == GlobalFiModInstNr[3]))));
	Tile mesh_6_6(
		.clock(clock),
		.io_in_a_0(r_102_0),
		.io_in_b_0(b_102_0),
		.io_in_d_0(b_358_0),
		.io_in_control_0_dataflow(mesh_6_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_6_io_in_control_0_shift_b),
		.io_in_id_0(r_614_0),
		.io_in_last_0(r_870_0),
		.io_in_valid_0(r_358_0),
		.io_out_a_0(_mesh_6_6_io_out_a_0),
		.io_out_c_0(_mesh_6_6_io_out_c_0),
		.io_out_b_0(_mesh_6_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_6_io_out_id_0),
		.io_out_last_0(_mesh_6_6_io_out_last_0),
		.io_out_valid_0(_mesh_6_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2497 == GlobalFiModInstNr[0]) || (2497 == GlobalFiModInstNr[1]) || (2497 == GlobalFiModInstNr[2]) || (2497 == GlobalFiModInstNr[3]))));
	Tile mesh_6_7(
		.clock(clock),
		.io_in_a_0(r_103_0),
		.io_in_b_0(b_118_0),
		.io_in_d_0(b_374_0),
		.io_in_control_0_dataflow(mesh_6_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_7_io_in_control_0_shift_b),
		.io_in_id_0(r_630_0),
		.io_in_last_0(r_886_0),
		.io_in_valid_0(r_374_0),
		.io_out_a_0(_mesh_6_7_io_out_a_0),
		.io_out_c_0(_mesh_6_7_io_out_c_0),
		.io_out_b_0(_mesh_6_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_7_io_out_id_0),
		.io_out_last_0(_mesh_6_7_io_out_last_0),
		.io_out_valid_0(_mesh_6_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2498 == GlobalFiModInstNr[0]) || (2498 == GlobalFiModInstNr[1]) || (2498 == GlobalFiModInstNr[2]) || (2498 == GlobalFiModInstNr[3]))));
	Tile mesh_6_8(
		.clock(clock),
		.io_in_a_0(r_104_0),
		.io_in_b_0(b_134_0),
		.io_in_d_0(b_390_0),
		.io_in_control_0_dataflow(mesh_6_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_8_io_in_control_0_shift_b),
		.io_in_id_0(r_646_0),
		.io_in_last_0(r_902_0),
		.io_in_valid_0(r_390_0),
		.io_out_a_0(_mesh_6_8_io_out_a_0),
		.io_out_c_0(_mesh_6_8_io_out_c_0),
		.io_out_b_0(_mesh_6_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_8_io_out_id_0),
		.io_out_last_0(_mesh_6_8_io_out_last_0),
		.io_out_valid_0(_mesh_6_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2499 == GlobalFiModInstNr[0]) || (2499 == GlobalFiModInstNr[1]) || (2499 == GlobalFiModInstNr[2]) || (2499 == GlobalFiModInstNr[3]))));
	Tile mesh_6_9(
		.clock(clock),
		.io_in_a_0(r_105_0),
		.io_in_b_0(b_150_0),
		.io_in_d_0(b_406_0),
		.io_in_control_0_dataflow(mesh_6_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_9_io_in_control_0_shift_b),
		.io_in_id_0(r_662_0),
		.io_in_last_0(r_918_0),
		.io_in_valid_0(r_406_0),
		.io_out_a_0(_mesh_6_9_io_out_a_0),
		.io_out_c_0(_mesh_6_9_io_out_c_0),
		.io_out_b_0(_mesh_6_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_9_io_out_id_0),
		.io_out_last_0(_mesh_6_9_io_out_last_0),
		.io_out_valid_0(_mesh_6_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2500 == GlobalFiModInstNr[0]) || (2500 == GlobalFiModInstNr[1]) || (2500 == GlobalFiModInstNr[2]) || (2500 == GlobalFiModInstNr[3]))));
	Tile mesh_6_10(
		.clock(clock),
		.io_in_a_0(r_106_0),
		.io_in_b_0(b_166_0),
		.io_in_d_0(b_422_0),
		.io_in_control_0_dataflow(mesh_6_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_10_io_in_control_0_shift_b),
		.io_in_id_0(r_678_0),
		.io_in_last_0(r_934_0),
		.io_in_valid_0(r_422_0),
		.io_out_a_0(_mesh_6_10_io_out_a_0),
		.io_out_c_0(_mesh_6_10_io_out_c_0),
		.io_out_b_0(_mesh_6_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_10_io_out_id_0),
		.io_out_last_0(_mesh_6_10_io_out_last_0),
		.io_out_valid_0(_mesh_6_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2501 == GlobalFiModInstNr[0]) || (2501 == GlobalFiModInstNr[1]) || (2501 == GlobalFiModInstNr[2]) || (2501 == GlobalFiModInstNr[3]))));
	Tile mesh_6_11(
		.clock(clock),
		.io_in_a_0(r_107_0),
		.io_in_b_0(b_182_0),
		.io_in_d_0(b_438_0),
		.io_in_control_0_dataflow(mesh_6_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_11_io_in_control_0_shift_b),
		.io_in_id_0(r_694_0),
		.io_in_last_0(r_950_0),
		.io_in_valid_0(r_438_0),
		.io_out_a_0(_mesh_6_11_io_out_a_0),
		.io_out_c_0(_mesh_6_11_io_out_c_0),
		.io_out_b_0(_mesh_6_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_11_io_out_id_0),
		.io_out_last_0(_mesh_6_11_io_out_last_0),
		.io_out_valid_0(_mesh_6_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2502 == GlobalFiModInstNr[0]) || (2502 == GlobalFiModInstNr[1]) || (2502 == GlobalFiModInstNr[2]) || (2502 == GlobalFiModInstNr[3]))));
	Tile mesh_6_12(
		.clock(clock),
		.io_in_a_0(r_108_0),
		.io_in_b_0(b_198_0),
		.io_in_d_0(b_454_0),
		.io_in_control_0_dataflow(mesh_6_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_12_io_in_control_0_shift_b),
		.io_in_id_0(r_710_0),
		.io_in_last_0(r_966_0),
		.io_in_valid_0(r_454_0),
		.io_out_a_0(_mesh_6_12_io_out_a_0),
		.io_out_c_0(_mesh_6_12_io_out_c_0),
		.io_out_b_0(_mesh_6_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_12_io_out_id_0),
		.io_out_last_0(_mesh_6_12_io_out_last_0),
		.io_out_valid_0(_mesh_6_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2503 == GlobalFiModInstNr[0]) || (2503 == GlobalFiModInstNr[1]) || (2503 == GlobalFiModInstNr[2]) || (2503 == GlobalFiModInstNr[3]))));
	Tile mesh_6_13(
		.clock(clock),
		.io_in_a_0(r_109_0),
		.io_in_b_0(b_214_0),
		.io_in_d_0(b_470_0),
		.io_in_control_0_dataflow(mesh_6_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_13_io_in_control_0_shift_b),
		.io_in_id_0(r_726_0),
		.io_in_last_0(r_982_0),
		.io_in_valid_0(r_470_0),
		.io_out_a_0(_mesh_6_13_io_out_a_0),
		.io_out_c_0(_mesh_6_13_io_out_c_0),
		.io_out_b_0(_mesh_6_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_13_io_out_id_0),
		.io_out_last_0(_mesh_6_13_io_out_last_0),
		.io_out_valid_0(_mesh_6_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2504 == GlobalFiModInstNr[0]) || (2504 == GlobalFiModInstNr[1]) || (2504 == GlobalFiModInstNr[2]) || (2504 == GlobalFiModInstNr[3]))));
	Tile mesh_6_14(
		.clock(clock),
		.io_in_a_0(r_110_0),
		.io_in_b_0(b_230_0),
		.io_in_d_0(b_486_0),
		.io_in_control_0_dataflow(mesh_6_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_14_io_in_control_0_shift_b),
		.io_in_id_0(r_742_0),
		.io_in_last_0(r_998_0),
		.io_in_valid_0(r_486_0),
		.io_out_a_0(_mesh_6_14_io_out_a_0),
		.io_out_c_0(_mesh_6_14_io_out_c_0),
		.io_out_b_0(_mesh_6_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_14_io_out_id_0),
		.io_out_last_0(_mesh_6_14_io_out_last_0),
		.io_out_valid_0(_mesh_6_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2505 == GlobalFiModInstNr[0]) || (2505 == GlobalFiModInstNr[1]) || (2505 == GlobalFiModInstNr[2]) || (2505 == GlobalFiModInstNr[3]))));
	Tile mesh_6_15(
		.clock(clock),
		.io_in_a_0(r_111_0),
		.io_in_b_0(b_246_0),
		.io_in_d_0(b_502_0),
		.io_in_control_0_dataflow(mesh_6_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_15_io_in_control_0_shift_b),
		.io_in_id_0(r_758_0),
		.io_in_last_0(r_1014_0),
		.io_in_valid_0(r_502_0),
		.io_out_a_0(_mesh_6_15_io_out_a_0),
		.io_out_c_0(_mesh_6_15_io_out_c_0),
		.io_out_b_0(_mesh_6_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_15_io_out_id_0),
		.io_out_last_0(_mesh_6_15_io_out_last_0),
		.io_out_valid_0(_mesh_6_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2506 == GlobalFiModInstNr[0]) || (2506 == GlobalFiModInstNr[1]) || (2506 == GlobalFiModInstNr[2]) || (2506 == GlobalFiModInstNr[3]))));
	Tile mesh_7_0(
		.clock(clock),
		.io_in_a_0(r_112_0),
		.io_in_b_0(b_7_0),
		.io_in_d_0(b_263_0),
		.io_in_control_0_dataflow(mesh_7_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_0_io_in_control_0_shift_b),
		.io_in_id_0(r_519_0),
		.io_in_last_0(r_775_0),
		.io_in_valid_0(r_263_0),
		.io_out_a_0(_mesh_7_0_io_out_a_0),
		.io_out_c_0(_mesh_7_0_io_out_c_0),
		.io_out_b_0(_mesh_7_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_0_io_out_id_0),
		.io_out_last_0(_mesh_7_0_io_out_last_0),
		.io_out_valid_0(_mesh_7_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2507 == GlobalFiModInstNr[0]) || (2507 == GlobalFiModInstNr[1]) || (2507 == GlobalFiModInstNr[2]) || (2507 == GlobalFiModInstNr[3]))));
	Tile mesh_7_1(
		.clock(clock),
		.io_in_a_0(r_113_0),
		.io_in_b_0(b_23_0),
		.io_in_d_0(b_279_0),
		.io_in_control_0_dataflow(mesh_7_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_1_io_in_control_0_shift_b),
		.io_in_id_0(r_535_0),
		.io_in_last_0(r_791_0),
		.io_in_valid_0(r_279_0),
		.io_out_a_0(_mesh_7_1_io_out_a_0),
		.io_out_c_0(_mesh_7_1_io_out_c_0),
		.io_out_b_0(_mesh_7_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_1_io_out_id_0),
		.io_out_last_0(_mesh_7_1_io_out_last_0),
		.io_out_valid_0(_mesh_7_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2508 == GlobalFiModInstNr[0]) || (2508 == GlobalFiModInstNr[1]) || (2508 == GlobalFiModInstNr[2]) || (2508 == GlobalFiModInstNr[3]))));
	Tile mesh_7_2(
		.clock(clock),
		.io_in_a_0(r_114_0),
		.io_in_b_0(b_39_0),
		.io_in_d_0(b_295_0),
		.io_in_control_0_dataflow(mesh_7_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_2_io_in_control_0_shift_b),
		.io_in_id_0(r_551_0),
		.io_in_last_0(r_807_0),
		.io_in_valid_0(r_295_0),
		.io_out_a_0(_mesh_7_2_io_out_a_0),
		.io_out_c_0(_mesh_7_2_io_out_c_0),
		.io_out_b_0(_mesh_7_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_2_io_out_id_0),
		.io_out_last_0(_mesh_7_2_io_out_last_0),
		.io_out_valid_0(_mesh_7_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2509 == GlobalFiModInstNr[0]) || (2509 == GlobalFiModInstNr[1]) || (2509 == GlobalFiModInstNr[2]) || (2509 == GlobalFiModInstNr[3]))));
	Tile mesh_7_3(
		.clock(clock),
		.io_in_a_0(r_115_0),
		.io_in_b_0(b_55_0),
		.io_in_d_0(b_311_0),
		.io_in_control_0_dataflow(mesh_7_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_3_io_in_control_0_shift_b),
		.io_in_id_0(r_567_0),
		.io_in_last_0(r_823_0),
		.io_in_valid_0(r_311_0),
		.io_out_a_0(_mesh_7_3_io_out_a_0),
		.io_out_c_0(_mesh_7_3_io_out_c_0),
		.io_out_b_0(_mesh_7_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_3_io_out_id_0),
		.io_out_last_0(_mesh_7_3_io_out_last_0),
		.io_out_valid_0(_mesh_7_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2510 == GlobalFiModInstNr[0]) || (2510 == GlobalFiModInstNr[1]) || (2510 == GlobalFiModInstNr[2]) || (2510 == GlobalFiModInstNr[3]))));
	Tile mesh_7_4(
		.clock(clock),
		.io_in_a_0(r_116_0),
		.io_in_b_0(b_71_0),
		.io_in_d_0(b_327_0),
		.io_in_control_0_dataflow(mesh_7_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_4_io_in_control_0_shift_b),
		.io_in_id_0(r_583_0),
		.io_in_last_0(r_839_0),
		.io_in_valid_0(r_327_0),
		.io_out_a_0(_mesh_7_4_io_out_a_0),
		.io_out_c_0(_mesh_7_4_io_out_c_0),
		.io_out_b_0(_mesh_7_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_4_io_out_id_0),
		.io_out_last_0(_mesh_7_4_io_out_last_0),
		.io_out_valid_0(_mesh_7_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2511 == GlobalFiModInstNr[0]) || (2511 == GlobalFiModInstNr[1]) || (2511 == GlobalFiModInstNr[2]) || (2511 == GlobalFiModInstNr[3]))));
	Tile mesh_7_5(
		.clock(clock),
		.io_in_a_0(r_117_0),
		.io_in_b_0(b_87_0),
		.io_in_d_0(b_343_0),
		.io_in_control_0_dataflow(mesh_7_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_5_io_in_control_0_shift_b),
		.io_in_id_0(r_599_0),
		.io_in_last_0(r_855_0),
		.io_in_valid_0(r_343_0),
		.io_out_a_0(_mesh_7_5_io_out_a_0),
		.io_out_c_0(_mesh_7_5_io_out_c_0),
		.io_out_b_0(_mesh_7_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_5_io_out_id_0),
		.io_out_last_0(_mesh_7_5_io_out_last_0),
		.io_out_valid_0(_mesh_7_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2512 == GlobalFiModInstNr[0]) || (2512 == GlobalFiModInstNr[1]) || (2512 == GlobalFiModInstNr[2]) || (2512 == GlobalFiModInstNr[3]))));
	Tile mesh_7_6(
		.clock(clock),
		.io_in_a_0(r_118_0),
		.io_in_b_0(b_103_0),
		.io_in_d_0(b_359_0),
		.io_in_control_0_dataflow(mesh_7_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_6_io_in_control_0_shift_b),
		.io_in_id_0(r_615_0),
		.io_in_last_0(r_871_0),
		.io_in_valid_0(r_359_0),
		.io_out_a_0(_mesh_7_6_io_out_a_0),
		.io_out_c_0(_mesh_7_6_io_out_c_0),
		.io_out_b_0(_mesh_7_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_6_io_out_id_0),
		.io_out_last_0(_mesh_7_6_io_out_last_0),
		.io_out_valid_0(_mesh_7_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2513 == GlobalFiModInstNr[0]) || (2513 == GlobalFiModInstNr[1]) || (2513 == GlobalFiModInstNr[2]) || (2513 == GlobalFiModInstNr[3]))));
	Tile mesh_7_7(
		.clock(clock),
		.io_in_a_0(r_119_0),
		.io_in_b_0(b_119_0),
		.io_in_d_0(b_375_0),
		.io_in_control_0_dataflow(mesh_7_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_7_io_in_control_0_shift_b),
		.io_in_id_0(r_631_0),
		.io_in_last_0(r_887_0),
		.io_in_valid_0(r_375_0),
		.io_out_a_0(_mesh_7_7_io_out_a_0),
		.io_out_c_0(_mesh_7_7_io_out_c_0),
		.io_out_b_0(_mesh_7_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_7_io_out_id_0),
		.io_out_last_0(_mesh_7_7_io_out_last_0),
		.io_out_valid_0(_mesh_7_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2514 == GlobalFiModInstNr[0]) || (2514 == GlobalFiModInstNr[1]) || (2514 == GlobalFiModInstNr[2]) || (2514 == GlobalFiModInstNr[3]))));
	Tile mesh_7_8(
		.clock(clock),
		.io_in_a_0(r_120_0),
		.io_in_b_0(b_135_0),
		.io_in_d_0(b_391_0),
		.io_in_control_0_dataflow(mesh_7_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_8_io_in_control_0_shift_b),
		.io_in_id_0(r_647_0),
		.io_in_last_0(r_903_0),
		.io_in_valid_0(r_391_0),
		.io_out_a_0(_mesh_7_8_io_out_a_0),
		.io_out_c_0(_mesh_7_8_io_out_c_0),
		.io_out_b_0(_mesh_7_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_8_io_out_id_0),
		.io_out_last_0(_mesh_7_8_io_out_last_0),
		.io_out_valid_0(_mesh_7_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2515 == GlobalFiModInstNr[0]) || (2515 == GlobalFiModInstNr[1]) || (2515 == GlobalFiModInstNr[2]) || (2515 == GlobalFiModInstNr[3]))));
	Tile mesh_7_9(
		.clock(clock),
		.io_in_a_0(r_121_0),
		.io_in_b_0(b_151_0),
		.io_in_d_0(b_407_0),
		.io_in_control_0_dataflow(mesh_7_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_9_io_in_control_0_shift_b),
		.io_in_id_0(r_663_0),
		.io_in_last_0(r_919_0),
		.io_in_valid_0(r_407_0),
		.io_out_a_0(_mesh_7_9_io_out_a_0),
		.io_out_c_0(_mesh_7_9_io_out_c_0),
		.io_out_b_0(_mesh_7_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_9_io_out_id_0),
		.io_out_last_0(_mesh_7_9_io_out_last_0),
		.io_out_valid_0(_mesh_7_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2516 == GlobalFiModInstNr[0]) || (2516 == GlobalFiModInstNr[1]) || (2516 == GlobalFiModInstNr[2]) || (2516 == GlobalFiModInstNr[3]))));
	Tile mesh_7_10(
		.clock(clock),
		.io_in_a_0(r_122_0),
		.io_in_b_0(b_167_0),
		.io_in_d_0(b_423_0),
		.io_in_control_0_dataflow(mesh_7_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_10_io_in_control_0_shift_b),
		.io_in_id_0(r_679_0),
		.io_in_last_0(r_935_0),
		.io_in_valid_0(r_423_0),
		.io_out_a_0(_mesh_7_10_io_out_a_0),
		.io_out_c_0(_mesh_7_10_io_out_c_0),
		.io_out_b_0(_mesh_7_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_10_io_out_id_0),
		.io_out_last_0(_mesh_7_10_io_out_last_0),
		.io_out_valid_0(_mesh_7_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2517 == GlobalFiModInstNr[0]) || (2517 == GlobalFiModInstNr[1]) || (2517 == GlobalFiModInstNr[2]) || (2517 == GlobalFiModInstNr[3]))));
	Tile mesh_7_11(
		.clock(clock),
		.io_in_a_0(r_123_0),
		.io_in_b_0(b_183_0),
		.io_in_d_0(b_439_0),
		.io_in_control_0_dataflow(mesh_7_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_11_io_in_control_0_shift_b),
		.io_in_id_0(r_695_0),
		.io_in_last_0(r_951_0),
		.io_in_valid_0(r_439_0),
		.io_out_a_0(_mesh_7_11_io_out_a_0),
		.io_out_c_0(_mesh_7_11_io_out_c_0),
		.io_out_b_0(_mesh_7_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_11_io_out_id_0),
		.io_out_last_0(_mesh_7_11_io_out_last_0),
		.io_out_valid_0(_mesh_7_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2518 == GlobalFiModInstNr[0]) || (2518 == GlobalFiModInstNr[1]) || (2518 == GlobalFiModInstNr[2]) || (2518 == GlobalFiModInstNr[3]))));
	Tile mesh_7_12(
		.clock(clock),
		.io_in_a_0(r_124_0),
		.io_in_b_0(b_199_0),
		.io_in_d_0(b_455_0),
		.io_in_control_0_dataflow(mesh_7_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_12_io_in_control_0_shift_b),
		.io_in_id_0(r_711_0),
		.io_in_last_0(r_967_0),
		.io_in_valid_0(r_455_0),
		.io_out_a_0(_mesh_7_12_io_out_a_0),
		.io_out_c_0(_mesh_7_12_io_out_c_0),
		.io_out_b_0(_mesh_7_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_12_io_out_id_0),
		.io_out_last_0(_mesh_7_12_io_out_last_0),
		.io_out_valid_0(_mesh_7_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2519 == GlobalFiModInstNr[0]) || (2519 == GlobalFiModInstNr[1]) || (2519 == GlobalFiModInstNr[2]) || (2519 == GlobalFiModInstNr[3]))));
	Tile mesh_7_13(
		.clock(clock),
		.io_in_a_0(r_125_0),
		.io_in_b_0(b_215_0),
		.io_in_d_0(b_471_0),
		.io_in_control_0_dataflow(mesh_7_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_13_io_in_control_0_shift_b),
		.io_in_id_0(r_727_0),
		.io_in_last_0(r_983_0),
		.io_in_valid_0(r_471_0),
		.io_out_a_0(_mesh_7_13_io_out_a_0),
		.io_out_c_0(_mesh_7_13_io_out_c_0),
		.io_out_b_0(_mesh_7_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_13_io_out_id_0),
		.io_out_last_0(_mesh_7_13_io_out_last_0),
		.io_out_valid_0(_mesh_7_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2520 == GlobalFiModInstNr[0]) || (2520 == GlobalFiModInstNr[1]) || (2520 == GlobalFiModInstNr[2]) || (2520 == GlobalFiModInstNr[3]))));
	Tile mesh_7_14(
		.clock(clock),
		.io_in_a_0(r_126_0),
		.io_in_b_0(b_231_0),
		.io_in_d_0(b_487_0),
		.io_in_control_0_dataflow(mesh_7_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_14_io_in_control_0_shift_b),
		.io_in_id_0(r_743_0),
		.io_in_last_0(r_999_0),
		.io_in_valid_0(r_487_0),
		.io_out_a_0(_mesh_7_14_io_out_a_0),
		.io_out_c_0(_mesh_7_14_io_out_c_0),
		.io_out_b_0(_mesh_7_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_14_io_out_id_0),
		.io_out_last_0(_mesh_7_14_io_out_last_0),
		.io_out_valid_0(_mesh_7_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2521 == GlobalFiModInstNr[0]) || (2521 == GlobalFiModInstNr[1]) || (2521 == GlobalFiModInstNr[2]) || (2521 == GlobalFiModInstNr[3]))));
	Tile mesh_7_15(
		.clock(clock),
		.io_in_a_0(r_127_0),
		.io_in_b_0(b_247_0),
		.io_in_d_0(b_503_0),
		.io_in_control_0_dataflow(mesh_7_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_15_io_in_control_0_shift_b),
		.io_in_id_0(r_759_0),
		.io_in_last_0(r_1015_0),
		.io_in_valid_0(r_503_0),
		.io_out_a_0(_mesh_7_15_io_out_a_0),
		.io_out_c_0(_mesh_7_15_io_out_c_0),
		.io_out_b_0(_mesh_7_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_15_io_out_id_0),
		.io_out_last_0(_mesh_7_15_io_out_last_0),
		.io_out_valid_0(_mesh_7_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2522 == GlobalFiModInstNr[0]) || (2522 == GlobalFiModInstNr[1]) || (2522 == GlobalFiModInstNr[2]) || (2522 == GlobalFiModInstNr[3]))));
	Tile mesh_8_0(
		.clock(clock),
		.io_in_a_0(r_128_0),
		.io_in_b_0(b_8_0),
		.io_in_d_0(b_264_0),
		.io_in_control_0_dataflow(mesh_8_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_0_io_in_control_0_shift_b),
		.io_in_id_0(r_520_0),
		.io_in_last_0(r_776_0),
		.io_in_valid_0(r_264_0),
		.io_out_a_0(_mesh_8_0_io_out_a_0),
		.io_out_c_0(_mesh_8_0_io_out_c_0),
		.io_out_b_0(_mesh_8_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_0_io_out_id_0),
		.io_out_last_0(_mesh_8_0_io_out_last_0),
		.io_out_valid_0(_mesh_8_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2523 == GlobalFiModInstNr[0]) || (2523 == GlobalFiModInstNr[1]) || (2523 == GlobalFiModInstNr[2]) || (2523 == GlobalFiModInstNr[3]))));
	Tile mesh_8_1(
		.clock(clock),
		.io_in_a_0(r_129_0),
		.io_in_b_0(b_24_0),
		.io_in_d_0(b_280_0),
		.io_in_control_0_dataflow(mesh_8_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_1_io_in_control_0_shift_b),
		.io_in_id_0(r_536_0),
		.io_in_last_0(r_792_0),
		.io_in_valid_0(r_280_0),
		.io_out_a_0(_mesh_8_1_io_out_a_0),
		.io_out_c_0(_mesh_8_1_io_out_c_0),
		.io_out_b_0(_mesh_8_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_1_io_out_id_0),
		.io_out_last_0(_mesh_8_1_io_out_last_0),
		.io_out_valid_0(_mesh_8_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2524 == GlobalFiModInstNr[0]) || (2524 == GlobalFiModInstNr[1]) || (2524 == GlobalFiModInstNr[2]) || (2524 == GlobalFiModInstNr[3]))));
	Tile mesh_8_2(
		.clock(clock),
		.io_in_a_0(r_130_0),
		.io_in_b_0(b_40_0),
		.io_in_d_0(b_296_0),
		.io_in_control_0_dataflow(mesh_8_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_2_io_in_control_0_shift_b),
		.io_in_id_0(r_552_0),
		.io_in_last_0(r_808_0),
		.io_in_valid_0(r_296_0),
		.io_out_a_0(_mesh_8_2_io_out_a_0),
		.io_out_c_0(_mesh_8_2_io_out_c_0),
		.io_out_b_0(_mesh_8_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_2_io_out_id_0),
		.io_out_last_0(_mesh_8_2_io_out_last_0),
		.io_out_valid_0(_mesh_8_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2525 == GlobalFiModInstNr[0]) || (2525 == GlobalFiModInstNr[1]) || (2525 == GlobalFiModInstNr[2]) || (2525 == GlobalFiModInstNr[3]))));
	Tile mesh_8_3(
		.clock(clock),
		.io_in_a_0(r_131_0),
		.io_in_b_0(b_56_0),
		.io_in_d_0(b_312_0),
		.io_in_control_0_dataflow(mesh_8_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_3_io_in_control_0_shift_b),
		.io_in_id_0(r_568_0),
		.io_in_last_0(r_824_0),
		.io_in_valid_0(r_312_0),
		.io_out_a_0(_mesh_8_3_io_out_a_0),
		.io_out_c_0(_mesh_8_3_io_out_c_0),
		.io_out_b_0(_mesh_8_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_3_io_out_id_0),
		.io_out_last_0(_mesh_8_3_io_out_last_0),
		.io_out_valid_0(_mesh_8_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2526 == GlobalFiModInstNr[0]) || (2526 == GlobalFiModInstNr[1]) || (2526 == GlobalFiModInstNr[2]) || (2526 == GlobalFiModInstNr[3]))));
	Tile mesh_8_4(
		.clock(clock),
		.io_in_a_0(r_132_0),
		.io_in_b_0(b_72_0),
		.io_in_d_0(b_328_0),
		.io_in_control_0_dataflow(mesh_8_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_4_io_in_control_0_shift_b),
		.io_in_id_0(r_584_0),
		.io_in_last_0(r_840_0),
		.io_in_valid_0(r_328_0),
		.io_out_a_0(_mesh_8_4_io_out_a_0),
		.io_out_c_0(_mesh_8_4_io_out_c_0),
		.io_out_b_0(_mesh_8_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_4_io_out_id_0),
		.io_out_last_0(_mesh_8_4_io_out_last_0),
		.io_out_valid_0(_mesh_8_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2527 == GlobalFiModInstNr[0]) || (2527 == GlobalFiModInstNr[1]) || (2527 == GlobalFiModInstNr[2]) || (2527 == GlobalFiModInstNr[3]))));
	Tile mesh_8_5(
		.clock(clock),
		.io_in_a_0(r_133_0),
		.io_in_b_0(b_88_0),
		.io_in_d_0(b_344_0),
		.io_in_control_0_dataflow(mesh_8_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_5_io_in_control_0_shift_b),
		.io_in_id_0(r_600_0),
		.io_in_last_0(r_856_0),
		.io_in_valid_0(r_344_0),
		.io_out_a_0(_mesh_8_5_io_out_a_0),
		.io_out_c_0(_mesh_8_5_io_out_c_0),
		.io_out_b_0(_mesh_8_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_5_io_out_id_0),
		.io_out_last_0(_mesh_8_5_io_out_last_0),
		.io_out_valid_0(_mesh_8_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2528 == GlobalFiModInstNr[0]) || (2528 == GlobalFiModInstNr[1]) || (2528 == GlobalFiModInstNr[2]) || (2528 == GlobalFiModInstNr[3]))));
	Tile mesh_8_6(
		.clock(clock),
		.io_in_a_0(r_134_0),
		.io_in_b_0(b_104_0),
		.io_in_d_0(b_360_0),
		.io_in_control_0_dataflow(mesh_8_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_6_io_in_control_0_shift_b),
		.io_in_id_0(r_616_0),
		.io_in_last_0(r_872_0),
		.io_in_valid_0(r_360_0),
		.io_out_a_0(_mesh_8_6_io_out_a_0),
		.io_out_c_0(_mesh_8_6_io_out_c_0),
		.io_out_b_0(_mesh_8_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_6_io_out_id_0),
		.io_out_last_0(_mesh_8_6_io_out_last_0),
		.io_out_valid_0(_mesh_8_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2529 == GlobalFiModInstNr[0]) || (2529 == GlobalFiModInstNr[1]) || (2529 == GlobalFiModInstNr[2]) || (2529 == GlobalFiModInstNr[3]))));
	Tile mesh_8_7(
		.clock(clock),
		.io_in_a_0(r_135_0),
		.io_in_b_0(b_120_0),
		.io_in_d_0(b_376_0),
		.io_in_control_0_dataflow(mesh_8_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_7_io_in_control_0_shift_b),
		.io_in_id_0(r_632_0),
		.io_in_last_0(r_888_0),
		.io_in_valid_0(r_376_0),
		.io_out_a_0(_mesh_8_7_io_out_a_0),
		.io_out_c_0(_mesh_8_7_io_out_c_0),
		.io_out_b_0(_mesh_8_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_7_io_out_id_0),
		.io_out_last_0(_mesh_8_7_io_out_last_0),
		.io_out_valid_0(_mesh_8_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2530 == GlobalFiModInstNr[0]) || (2530 == GlobalFiModInstNr[1]) || (2530 == GlobalFiModInstNr[2]) || (2530 == GlobalFiModInstNr[3]))));
	Tile mesh_8_8(
		.clock(clock),
		.io_in_a_0(r_136_0),
		.io_in_b_0(b_136_0),
		.io_in_d_0(b_392_0),
		.io_in_control_0_dataflow(mesh_8_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_8_io_in_control_0_shift_b),
		.io_in_id_0(r_648_0),
		.io_in_last_0(r_904_0),
		.io_in_valid_0(r_392_0),
		.io_out_a_0(_mesh_8_8_io_out_a_0),
		.io_out_c_0(_mesh_8_8_io_out_c_0),
		.io_out_b_0(_mesh_8_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_8_io_out_id_0),
		.io_out_last_0(_mesh_8_8_io_out_last_0),
		.io_out_valid_0(_mesh_8_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2531 == GlobalFiModInstNr[0]) || (2531 == GlobalFiModInstNr[1]) || (2531 == GlobalFiModInstNr[2]) || (2531 == GlobalFiModInstNr[3]))));
	Tile mesh_8_9(
		.clock(clock),
		.io_in_a_0(r_137_0),
		.io_in_b_0(b_152_0),
		.io_in_d_0(b_408_0),
		.io_in_control_0_dataflow(mesh_8_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_9_io_in_control_0_shift_b),
		.io_in_id_0(r_664_0),
		.io_in_last_0(r_920_0),
		.io_in_valid_0(r_408_0),
		.io_out_a_0(_mesh_8_9_io_out_a_0),
		.io_out_c_0(_mesh_8_9_io_out_c_0),
		.io_out_b_0(_mesh_8_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_9_io_out_id_0),
		.io_out_last_0(_mesh_8_9_io_out_last_0),
		.io_out_valid_0(_mesh_8_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2532 == GlobalFiModInstNr[0]) || (2532 == GlobalFiModInstNr[1]) || (2532 == GlobalFiModInstNr[2]) || (2532 == GlobalFiModInstNr[3]))));
	Tile mesh_8_10(
		.clock(clock),
		.io_in_a_0(r_138_0),
		.io_in_b_0(b_168_0),
		.io_in_d_0(b_424_0),
		.io_in_control_0_dataflow(mesh_8_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_10_io_in_control_0_shift_b),
		.io_in_id_0(r_680_0),
		.io_in_last_0(r_936_0),
		.io_in_valid_0(r_424_0),
		.io_out_a_0(_mesh_8_10_io_out_a_0),
		.io_out_c_0(_mesh_8_10_io_out_c_0),
		.io_out_b_0(_mesh_8_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_10_io_out_id_0),
		.io_out_last_0(_mesh_8_10_io_out_last_0),
		.io_out_valid_0(_mesh_8_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2533 == GlobalFiModInstNr[0]) || (2533 == GlobalFiModInstNr[1]) || (2533 == GlobalFiModInstNr[2]) || (2533 == GlobalFiModInstNr[3]))));
	Tile mesh_8_11(
		.clock(clock),
		.io_in_a_0(r_139_0),
		.io_in_b_0(b_184_0),
		.io_in_d_0(b_440_0),
		.io_in_control_0_dataflow(mesh_8_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_11_io_in_control_0_shift_b),
		.io_in_id_0(r_696_0),
		.io_in_last_0(r_952_0),
		.io_in_valid_0(r_440_0),
		.io_out_a_0(_mesh_8_11_io_out_a_0),
		.io_out_c_0(_mesh_8_11_io_out_c_0),
		.io_out_b_0(_mesh_8_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_11_io_out_id_0),
		.io_out_last_0(_mesh_8_11_io_out_last_0),
		.io_out_valid_0(_mesh_8_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2534 == GlobalFiModInstNr[0]) || (2534 == GlobalFiModInstNr[1]) || (2534 == GlobalFiModInstNr[2]) || (2534 == GlobalFiModInstNr[3]))));
	Tile mesh_8_12(
		.clock(clock),
		.io_in_a_0(r_140_0),
		.io_in_b_0(b_200_0),
		.io_in_d_0(b_456_0),
		.io_in_control_0_dataflow(mesh_8_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_12_io_in_control_0_shift_b),
		.io_in_id_0(r_712_0),
		.io_in_last_0(r_968_0),
		.io_in_valid_0(r_456_0),
		.io_out_a_0(_mesh_8_12_io_out_a_0),
		.io_out_c_0(_mesh_8_12_io_out_c_0),
		.io_out_b_0(_mesh_8_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_12_io_out_id_0),
		.io_out_last_0(_mesh_8_12_io_out_last_0),
		.io_out_valid_0(_mesh_8_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2535 == GlobalFiModInstNr[0]) || (2535 == GlobalFiModInstNr[1]) || (2535 == GlobalFiModInstNr[2]) || (2535 == GlobalFiModInstNr[3]))));
	Tile mesh_8_13(
		.clock(clock),
		.io_in_a_0(r_141_0),
		.io_in_b_0(b_216_0),
		.io_in_d_0(b_472_0),
		.io_in_control_0_dataflow(mesh_8_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_13_io_in_control_0_shift_b),
		.io_in_id_0(r_728_0),
		.io_in_last_0(r_984_0),
		.io_in_valid_0(r_472_0),
		.io_out_a_0(_mesh_8_13_io_out_a_0),
		.io_out_c_0(_mesh_8_13_io_out_c_0),
		.io_out_b_0(_mesh_8_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_13_io_out_id_0),
		.io_out_last_0(_mesh_8_13_io_out_last_0),
		.io_out_valid_0(_mesh_8_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2536 == GlobalFiModInstNr[0]) || (2536 == GlobalFiModInstNr[1]) || (2536 == GlobalFiModInstNr[2]) || (2536 == GlobalFiModInstNr[3]))));
	Tile mesh_8_14(
		.clock(clock),
		.io_in_a_0(r_142_0),
		.io_in_b_0(b_232_0),
		.io_in_d_0(b_488_0),
		.io_in_control_0_dataflow(mesh_8_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_14_io_in_control_0_shift_b),
		.io_in_id_0(r_744_0),
		.io_in_last_0(r_1000_0),
		.io_in_valid_0(r_488_0),
		.io_out_a_0(_mesh_8_14_io_out_a_0),
		.io_out_c_0(_mesh_8_14_io_out_c_0),
		.io_out_b_0(_mesh_8_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_14_io_out_id_0),
		.io_out_last_0(_mesh_8_14_io_out_last_0),
		.io_out_valid_0(_mesh_8_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2537 == GlobalFiModInstNr[0]) || (2537 == GlobalFiModInstNr[1]) || (2537 == GlobalFiModInstNr[2]) || (2537 == GlobalFiModInstNr[3]))));
	Tile mesh_8_15(
		.clock(clock),
		.io_in_a_0(r_143_0),
		.io_in_b_0(b_248_0),
		.io_in_d_0(b_504_0),
		.io_in_control_0_dataflow(mesh_8_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_15_io_in_control_0_shift_b),
		.io_in_id_0(r_760_0),
		.io_in_last_0(r_1016_0),
		.io_in_valid_0(r_504_0),
		.io_out_a_0(_mesh_8_15_io_out_a_0),
		.io_out_c_0(_mesh_8_15_io_out_c_0),
		.io_out_b_0(_mesh_8_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_15_io_out_id_0),
		.io_out_last_0(_mesh_8_15_io_out_last_0),
		.io_out_valid_0(_mesh_8_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2538 == GlobalFiModInstNr[0]) || (2538 == GlobalFiModInstNr[1]) || (2538 == GlobalFiModInstNr[2]) || (2538 == GlobalFiModInstNr[3]))));
	Tile mesh_9_0(
		.clock(clock),
		.io_in_a_0(r_144_0),
		.io_in_b_0(b_9_0),
		.io_in_d_0(b_265_0),
		.io_in_control_0_dataflow(mesh_9_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_0_io_in_control_0_shift_b),
		.io_in_id_0(r_521_0),
		.io_in_last_0(r_777_0),
		.io_in_valid_0(r_265_0),
		.io_out_a_0(_mesh_9_0_io_out_a_0),
		.io_out_c_0(_mesh_9_0_io_out_c_0),
		.io_out_b_0(_mesh_9_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_0_io_out_id_0),
		.io_out_last_0(_mesh_9_0_io_out_last_0),
		.io_out_valid_0(_mesh_9_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2539 == GlobalFiModInstNr[0]) || (2539 == GlobalFiModInstNr[1]) || (2539 == GlobalFiModInstNr[2]) || (2539 == GlobalFiModInstNr[3]))));
	Tile mesh_9_1(
		.clock(clock),
		.io_in_a_0(r_145_0),
		.io_in_b_0(b_25_0),
		.io_in_d_0(b_281_0),
		.io_in_control_0_dataflow(mesh_9_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_1_io_in_control_0_shift_b),
		.io_in_id_0(r_537_0),
		.io_in_last_0(r_793_0),
		.io_in_valid_0(r_281_0),
		.io_out_a_0(_mesh_9_1_io_out_a_0),
		.io_out_c_0(_mesh_9_1_io_out_c_0),
		.io_out_b_0(_mesh_9_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_1_io_out_id_0),
		.io_out_last_0(_mesh_9_1_io_out_last_0),
		.io_out_valid_0(_mesh_9_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2540 == GlobalFiModInstNr[0]) || (2540 == GlobalFiModInstNr[1]) || (2540 == GlobalFiModInstNr[2]) || (2540 == GlobalFiModInstNr[3]))));
	Tile mesh_9_2(
		.clock(clock),
		.io_in_a_0(r_146_0),
		.io_in_b_0(b_41_0),
		.io_in_d_0(b_297_0),
		.io_in_control_0_dataflow(mesh_9_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_2_io_in_control_0_shift_b),
		.io_in_id_0(r_553_0),
		.io_in_last_0(r_809_0),
		.io_in_valid_0(r_297_0),
		.io_out_a_0(_mesh_9_2_io_out_a_0),
		.io_out_c_0(_mesh_9_2_io_out_c_0),
		.io_out_b_0(_mesh_9_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_2_io_out_id_0),
		.io_out_last_0(_mesh_9_2_io_out_last_0),
		.io_out_valid_0(_mesh_9_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2541 == GlobalFiModInstNr[0]) || (2541 == GlobalFiModInstNr[1]) || (2541 == GlobalFiModInstNr[2]) || (2541 == GlobalFiModInstNr[3]))));
	Tile mesh_9_3(
		.clock(clock),
		.io_in_a_0(r_147_0),
		.io_in_b_0(b_57_0),
		.io_in_d_0(b_313_0),
		.io_in_control_0_dataflow(mesh_9_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_3_io_in_control_0_shift_b),
		.io_in_id_0(r_569_0),
		.io_in_last_0(r_825_0),
		.io_in_valid_0(r_313_0),
		.io_out_a_0(_mesh_9_3_io_out_a_0),
		.io_out_c_0(_mesh_9_3_io_out_c_0),
		.io_out_b_0(_mesh_9_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_3_io_out_id_0),
		.io_out_last_0(_mesh_9_3_io_out_last_0),
		.io_out_valid_0(_mesh_9_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2542 == GlobalFiModInstNr[0]) || (2542 == GlobalFiModInstNr[1]) || (2542 == GlobalFiModInstNr[2]) || (2542 == GlobalFiModInstNr[3]))));
	Tile mesh_9_4(
		.clock(clock),
		.io_in_a_0(r_148_0),
		.io_in_b_0(b_73_0),
		.io_in_d_0(b_329_0),
		.io_in_control_0_dataflow(mesh_9_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_4_io_in_control_0_shift_b),
		.io_in_id_0(r_585_0),
		.io_in_last_0(r_841_0),
		.io_in_valid_0(r_329_0),
		.io_out_a_0(_mesh_9_4_io_out_a_0),
		.io_out_c_0(_mesh_9_4_io_out_c_0),
		.io_out_b_0(_mesh_9_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_4_io_out_id_0),
		.io_out_last_0(_mesh_9_4_io_out_last_0),
		.io_out_valid_0(_mesh_9_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2543 == GlobalFiModInstNr[0]) || (2543 == GlobalFiModInstNr[1]) || (2543 == GlobalFiModInstNr[2]) || (2543 == GlobalFiModInstNr[3]))));
	Tile mesh_9_5(
		.clock(clock),
		.io_in_a_0(r_149_0),
		.io_in_b_0(b_89_0),
		.io_in_d_0(b_345_0),
		.io_in_control_0_dataflow(mesh_9_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_5_io_in_control_0_shift_b),
		.io_in_id_0(r_601_0),
		.io_in_last_0(r_857_0),
		.io_in_valid_0(r_345_0),
		.io_out_a_0(_mesh_9_5_io_out_a_0),
		.io_out_c_0(_mesh_9_5_io_out_c_0),
		.io_out_b_0(_mesh_9_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_5_io_out_id_0),
		.io_out_last_0(_mesh_9_5_io_out_last_0),
		.io_out_valid_0(_mesh_9_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2544 == GlobalFiModInstNr[0]) || (2544 == GlobalFiModInstNr[1]) || (2544 == GlobalFiModInstNr[2]) || (2544 == GlobalFiModInstNr[3]))));
	Tile mesh_9_6(
		.clock(clock),
		.io_in_a_0(r_150_0),
		.io_in_b_0(b_105_0),
		.io_in_d_0(b_361_0),
		.io_in_control_0_dataflow(mesh_9_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_6_io_in_control_0_shift_b),
		.io_in_id_0(r_617_0),
		.io_in_last_0(r_873_0),
		.io_in_valid_0(r_361_0),
		.io_out_a_0(_mesh_9_6_io_out_a_0),
		.io_out_c_0(_mesh_9_6_io_out_c_0),
		.io_out_b_0(_mesh_9_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_6_io_out_id_0),
		.io_out_last_0(_mesh_9_6_io_out_last_0),
		.io_out_valid_0(_mesh_9_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2545 == GlobalFiModInstNr[0]) || (2545 == GlobalFiModInstNr[1]) || (2545 == GlobalFiModInstNr[2]) || (2545 == GlobalFiModInstNr[3]))));
	Tile mesh_9_7(
		.clock(clock),
		.io_in_a_0(r_151_0),
		.io_in_b_0(b_121_0),
		.io_in_d_0(b_377_0),
		.io_in_control_0_dataflow(mesh_9_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_7_io_in_control_0_shift_b),
		.io_in_id_0(r_633_0),
		.io_in_last_0(r_889_0),
		.io_in_valid_0(r_377_0),
		.io_out_a_0(_mesh_9_7_io_out_a_0),
		.io_out_c_0(_mesh_9_7_io_out_c_0),
		.io_out_b_0(_mesh_9_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_7_io_out_id_0),
		.io_out_last_0(_mesh_9_7_io_out_last_0),
		.io_out_valid_0(_mesh_9_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2546 == GlobalFiModInstNr[0]) || (2546 == GlobalFiModInstNr[1]) || (2546 == GlobalFiModInstNr[2]) || (2546 == GlobalFiModInstNr[3]))));
	Tile mesh_9_8(
		.clock(clock),
		.io_in_a_0(r_152_0),
		.io_in_b_0(b_137_0),
		.io_in_d_0(b_393_0),
		.io_in_control_0_dataflow(mesh_9_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_8_io_in_control_0_shift_b),
		.io_in_id_0(r_649_0),
		.io_in_last_0(r_905_0),
		.io_in_valid_0(r_393_0),
		.io_out_a_0(_mesh_9_8_io_out_a_0),
		.io_out_c_0(_mesh_9_8_io_out_c_0),
		.io_out_b_0(_mesh_9_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_8_io_out_id_0),
		.io_out_last_0(_mesh_9_8_io_out_last_0),
		.io_out_valid_0(_mesh_9_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2547 == GlobalFiModInstNr[0]) || (2547 == GlobalFiModInstNr[1]) || (2547 == GlobalFiModInstNr[2]) || (2547 == GlobalFiModInstNr[3]))));
	Tile mesh_9_9(
		.clock(clock),
		.io_in_a_0(r_153_0),
		.io_in_b_0(b_153_0),
		.io_in_d_0(b_409_0),
		.io_in_control_0_dataflow(mesh_9_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_9_io_in_control_0_shift_b),
		.io_in_id_0(r_665_0),
		.io_in_last_0(r_921_0),
		.io_in_valid_0(r_409_0),
		.io_out_a_0(_mesh_9_9_io_out_a_0),
		.io_out_c_0(_mesh_9_9_io_out_c_0),
		.io_out_b_0(_mesh_9_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_9_io_out_id_0),
		.io_out_last_0(_mesh_9_9_io_out_last_0),
		.io_out_valid_0(_mesh_9_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2548 == GlobalFiModInstNr[0]) || (2548 == GlobalFiModInstNr[1]) || (2548 == GlobalFiModInstNr[2]) || (2548 == GlobalFiModInstNr[3]))));
	Tile mesh_9_10(
		.clock(clock),
		.io_in_a_0(r_154_0),
		.io_in_b_0(b_169_0),
		.io_in_d_0(b_425_0),
		.io_in_control_0_dataflow(mesh_9_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_10_io_in_control_0_shift_b),
		.io_in_id_0(r_681_0),
		.io_in_last_0(r_937_0),
		.io_in_valid_0(r_425_0),
		.io_out_a_0(_mesh_9_10_io_out_a_0),
		.io_out_c_0(_mesh_9_10_io_out_c_0),
		.io_out_b_0(_mesh_9_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_10_io_out_id_0),
		.io_out_last_0(_mesh_9_10_io_out_last_0),
		.io_out_valid_0(_mesh_9_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2549 == GlobalFiModInstNr[0]) || (2549 == GlobalFiModInstNr[1]) || (2549 == GlobalFiModInstNr[2]) || (2549 == GlobalFiModInstNr[3]))));
	Tile mesh_9_11(
		.clock(clock),
		.io_in_a_0(r_155_0),
		.io_in_b_0(b_185_0),
		.io_in_d_0(b_441_0),
		.io_in_control_0_dataflow(mesh_9_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_11_io_in_control_0_shift_b),
		.io_in_id_0(r_697_0),
		.io_in_last_0(r_953_0),
		.io_in_valid_0(r_441_0),
		.io_out_a_0(_mesh_9_11_io_out_a_0),
		.io_out_c_0(_mesh_9_11_io_out_c_0),
		.io_out_b_0(_mesh_9_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_11_io_out_id_0),
		.io_out_last_0(_mesh_9_11_io_out_last_0),
		.io_out_valid_0(_mesh_9_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2550 == GlobalFiModInstNr[0]) || (2550 == GlobalFiModInstNr[1]) || (2550 == GlobalFiModInstNr[2]) || (2550 == GlobalFiModInstNr[3]))));
	Tile mesh_9_12(
		.clock(clock),
		.io_in_a_0(r_156_0),
		.io_in_b_0(b_201_0),
		.io_in_d_0(b_457_0),
		.io_in_control_0_dataflow(mesh_9_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_12_io_in_control_0_shift_b),
		.io_in_id_0(r_713_0),
		.io_in_last_0(r_969_0),
		.io_in_valid_0(r_457_0),
		.io_out_a_0(_mesh_9_12_io_out_a_0),
		.io_out_c_0(_mesh_9_12_io_out_c_0),
		.io_out_b_0(_mesh_9_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_12_io_out_id_0),
		.io_out_last_0(_mesh_9_12_io_out_last_0),
		.io_out_valid_0(_mesh_9_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2551 == GlobalFiModInstNr[0]) || (2551 == GlobalFiModInstNr[1]) || (2551 == GlobalFiModInstNr[2]) || (2551 == GlobalFiModInstNr[3]))));
	Tile mesh_9_13(
		.clock(clock),
		.io_in_a_0(r_157_0),
		.io_in_b_0(b_217_0),
		.io_in_d_0(b_473_0),
		.io_in_control_0_dataflow(mesh_9_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_13_io_in_control_0_shift_b),
		.io_in_id_0(r_729_0),
		.io_in_last_0(r_985_0),
		.io_in_valid_0(r_473_0),
		.io_out_a_0(_mesh_9_13_io_out_a_0),
		.io_out_c_0(_mesh_9_13_io_out_c_0),
		.io_out_b_0(_mesh_9_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_13_io_out_id_0),
		.io_out_last_0(_mesh_9_13_io_out_last_0),
		.io_out_valid_0(_mesh_9_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2552 == GlobalFiModInstNr[0]) || (2552 == GlobalFiModInstNr[1]) || (2552 == GlobalFiModInstNr[2]) || (2552 == GlobalFiModInstNr[3]))));
	Tile mesh_9_14(
		.clock(clock),
		.io_in_a_0(r_158_0),
		.io_in_b_0(b_233_0),
		.io_in_d_0(b_489_0),
		.io_in_control_0_dataflow(mesh_9_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_14_io_in_control_0_shift_b),
		.io_in_id_0(r_745_0),
		.io_in_last_0(r_1001_0),
		.io_in_valid_0(r_489_0),
		.io_out_a_0(_mesh_9_14_io_out_a_0),
		.io_out_c_0(_mesh_9_14_io_out_c_0),
		.io_out_b_0(_mesh_9_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_14_io_out_id_0),
		.io_out_last_0(_mesh_9_14_io_out_last_0),
		.io_out_valid_0(_mesh_9_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2553 == GlobalFiModInstNr[0]) || (2553 == GlobalFiModInstNr[1]) || (2553 == GlobalFiModInstNr[2]) || (2553 == GlobalFiModInstNr[3]))));
	Tile mesh_9_15(
		.clock(clock),
		.io_in_a_0(r_159_0),
		.io_in_b_0(b_249_0),
		.io_in_d_0(b_505_0),
		.io_in_control_0_dataflow(mesh_9_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_15_io_in_control_0_shift_b),
		.io_in_id_0(r_761_0),
		.io_in_last_0(r_1017_0),
		.io_in_valid_0(r_505_0),
		.io_out_a_0(_mesh_9_15_io_out_a_0),
		.io_out_c_0(_mesh_9_15_io_out_c_0),
		.io_out_b_0(_mesh_9_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_15_io_out_id_0),
		.io_out_last_0(_mesh_9_15_io_out_last_0),
		.io_out_valid_0(_mesh_9_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2554 == GlobalFiModInstNr[0]) || (2554 == GlobalFiModInstNr[1]) || (2554 == GlobalFiModInstNr[2]) || (2554 == GlobalFiModInstNr[3]))));
	Tile mesh_10_0(
		.clock(clock),
		.io_in_a_0(r_160_0),
		.io_in_b_0(b_10_0),
		.io_in_d_0(b_266_0),
		.io_in_control_0_dataflow(mesh_10_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_0_io_in_control_0_shift_b),
		.io_in_id_0(r_522_0),
		.io_in_last_0(r_778_0),
		.io_in_valid_0(r_266_0),
		.io_out_a_0(_mesh_10_0_io_out_a_0),
		.io_out_c_0(_mesh_10_0_io_out_c_0),
		.io_out_b_0(_mesh_10_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_0_io_out_id_0),
		.io_out_last_0(_mesh_10_0_io_out_last_0),
		.io_out_valid_0(_mesh_10_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2555 == GlobalFiModInstNr[0]) || (2555 == GlobalFiModInstNr[1]) || (2555 == GlobalFiModInstNr[2]) || (2555 == GlobalFiModInstNr[3]))));
	Tile mesh_10_1(
		.clock(clock),
		.io_in_a_0(r_161_0),
		.io_in_b_0(b_26_0),
		.io_in_d_0(b_282_0),
		.io_in_control_0_dataflow(mesh_10_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_1_io_in_control_0_shift_b),
		.io_in_id_0(r_538_0),
		.io_in_last_0(r_794_0),
		.io_in_valid_0(r_282_0),
		.io_out_a_0(_mesh_10_1_io_out_a_0),
		.io_out_c_0(_mesh_10_1_io_out_c_0),
		.io_out_b_0(_mesh_10_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_1_io_out_id_0),
		.io_out_last_0(_mesh_10_1_io_out_last_0),
		.io_out_valid_0(_mesh_10_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2556 == GlobalFiModInstNr[0]) || (2556 == GlobalFiModInstNr[1]) || (2556 == GlobalFiModInstNr[2]) || (2556 == GlobalFiModInstNr[3]))));
	Tile mesh_10_2(
		.clock(clock),
		.io_in_a_0(r_162_0),
		.io_in_b_0(b_42_0),
		.io_in_d_0(b_298_0),
		.io_in_control_0_dataflow(mesh_10_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_2_io_in_control_0_shift_b),
		.io_in_id_0(r_554_0),
		.io_in_last_0(r_810_0),
		.io_in_valid_0(r_298_0),
		.io_out_a_0(_mesh_10_2_io_out_a_0),
		.io_out_c_0(_mesh_10_2_io_out_c_0),
		.io_out_b_0(_mesh_10_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_2_io_out_id_0),
		.io_out_last_0(_mesh_10_2_io_out_last_0),
		.io_out_valid_0(_mesh_10_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2557 == GlobalFiModInstNr[0]) || (2557 == GlobalFiModInstNr[1]) || (2557 == GlobalFiModInstNr[2]) || (2557 == GlobalFiModInstNr[3]))));
	Tile mesh_10_3(
		.clock(clock),
		.io_in_a_0(r_163_0),
		.io_in_b_0(b_58_0),
		.io_in_d_0(b_314_0),
		.io_in_control_0_dataflow(mesh_10_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_3_io_in_control_0_shift_b),
		.io_in_id_0(r_570_0),
		.io_in_last_0(r_826_0),
		.io_in_valid_0(r_314_0),
		.io_out_a_0(_mesh_10_3_io_out_a_0),
		.io_out_c_0(_mesh_10_3_io_out_c_0),
		.io_out_b_0(_mesh_10_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_3_io_out_id_0),
		.io_out_last_0(_mesh_10_3_io_out_last_0),
		.io_out_valid_0(_mesh_10_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2558 == GlobalFiModInstNr[0]) || (2558 == GlobalFiModInstNr[1]) || (2558 == GlobalFiModInstNr[2]) || (2558 == GlobalFiModInstNr[3]))));
	Tile mesh_10_4(
		.clock(clock),
		.io_in_a_0(r_164_0),
		.io_in_b_0(b_74_0),
		.io_in_d_0(b_330_0),
		.io_in_control_0_dataflow(mesh_10_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_4_io_in_control_0_shift_b),
		.io_in_id_0(r_586_0),
		.io_in_last_0(r_842_0),
		.io_in_valid_0(r_330_0),
		.io_out_a_0(_mesh_10_4_io_out_a_0),
		.io_out_c_0(_mesh_10_4_io_out_c_0),
		.io_out_b_0(_mesh_10_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_4_io_out_id_0),
		.io_out_last_0(_mesh_10_4_io_out_last_0),
		.io_out_valid_0(_mesh_10_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2559 == GlobalFiModInstNr[0]) || (2559 == GlobalFiModInstNr[1]) || (2559 == GlobalFiModInstNr[2]) || (2559 == GlobalFiModInstNr[3]))));
	Tile mesh_10_5(
		.clock(clock),
		.io_in_a_0(r_165_0),
		.io_in_b_0(b_90_0),
		.io_in_d_0(b_346_0),
		.io_in_control_0_dataflow(mesh_10_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_5_io_in_control_0_shift_b),
		.io_in_id_0(r_602_0),
		.io_in_last_0(r_858_0),
		.io_in_valid_0(r_346_0),
		.io_out_a_0(_mesh_10_5_io_out_a_0),
		.io_out_c_0(_mesh_10_5_io_out_c_0),
		.io_out_b_0(_mesh_10_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_5_io_out_id_0),
		.io_out_last_0(_mesh_10_5_io_out_last_0),
		.io_out_valid_0(_mesh_10_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2560 == GlobalFiModInstNr[0]) || (2560 == GlobalFiModInstNr[1]) || (2560 == GlobalFiModInstNr[2]) || (2560 == GlobalFiModInstNr[3]))));
	Tile mesh_10_6(
		.clock(clock),
		.io_in_a_0(r_166_0),
		.io_in_b_0(b_106_0),
		.io_in_d_0(b_362_0),
		.io_in_control_0_dataflow(mesh_10_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_6_io_in_control_0_shift_b),
		.io_in_id_0(r_618_0),
		.io_in_last_0(r_874_0),
		.io_in_valid_0(r_362_0),
		.io_out_a_0(_mesh_10_6_io_out_a_0),
		.io_out_c_0(_mesh_10_6_io_out_c_0),
		.io_out_b_0(_mesh_10_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_6_io_out_id_0),
		.io_out_last_0(_mesh_10_6_io_out_last_0),
		.io_out_valid_0(_mesh_10_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2561 == GlobalFiModInstNr[0]) || (2561 == GlobalFiModInstNr[1]) || (2561 == GlobalFiModInstNr[2]) || (2561 == GlobalFiModInstNr[3]))));
	Tile mesh_10_7(
		.clock(clock),
		.io_in_a_0(r_167_0),
		.io_in_b_0(b_122_0),
		.io_in_d_0(b_378_0),
		.io_in_control_0_dataflow(mesh_10_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_7_io_in_control_0_shift_b),
		.io_in_id_0(r_634_0),
		.io_in_last_0(r_890_0),
		.io_in_valid_0(r_378_0),
		.io_out_a_0(_mesh_10_7_io_out_a_0),
		.io_out_c_0(_mesh_10_7_io_out_c_0),
		.io_out_b_0(_mesh_10_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_7_io_out_id_0),
		.io_out_last_0(_mesh_10_7_io_out_last_0),
		.io_out_valid_0(_mesh_10_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2562 == GlobalFiModInstNr[0]) || (2562 == GlobalFiModInstNr[1]) || (2562 == GlobalFiModInstNr[2]) || (2562 == GlobalFiModInstNr[3]))));
	Tile mesh_10_8(
		.clock(clock),
		.io_in_a_0(r_168_0),
		.io_in_b_0(b_138_0),
		.io_in_d_0(b_394_0),
		.io_in_control_0_dataflow(mesh_10_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_8_io_in_control_0_shift_b),
		.io_in_id_0(r_650_0),
		.io_in_last_0(r_906_0),
		.io_in_valid_0(r_394_0),
		.io_out_a_0(_mesh_10_8_io_out_a_0),
		.io_out_c_0(_mesh_10_8_io_out_c_0),
		.io_out_b_0(_mesh_10_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_8_io_out_id_0),
		.io_out_last_0(_mesh_10_8_io_out_last_0),
		.io_out_valid_0(_mesh_10_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2563 == GlobalFiModInstNr[0]) || (2563 == GlobalFiModInstNr[1]) || (2563 == GlobalFiModInstNr[2]) || (2563 == GlobalFiModInstNr[3]))));
	Tile mesh_10_9(
		.clock(clock),
		.io_in_a_0(r_169_0),
		.io_in_b_0(b_154_0),
		.io_in_d_0(b_410_0),
		.io_in_control_0_dataflow(mesh_10_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_9_io_in_control_0_shift_b),
		.io_in_id_0(r_666_0),
		.io_in_last_0(r_922_0),
		.io_in_valid_0(r_410_0),
		.io_out_a_0(_mesh_10_9_io_out_a_0),
		.io_out_c_0(_mesh_10_9_io_out_c_0),
		.io_out_b_0(_mesh_10_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_9_io_out_id_0),
		.io_out_last_0(_mesh_10_9_io_out_last_0),
		.io_out_valid_0(_mesh_10_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2564 == GlobalFiModInstNr[0]) || (2564 == GlobalFiModInstNr[1]) || (2564 == GlobalFiModInstNr[2]) || (2564 == GlobalFiModInstNr[3]))));
	Tile mesh_10_10(
		.clock(clock),
		.io_in_a_0(r_170_0),
		.io_in_b_0(b_170_0),
		.io_in_d_0(b_426_0),
		.io_in_control_0_dataflow(mesh_10_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_10_io_in_control_0_shift_b),
		.io_in_id_0(r_682_0),
		.io_in_last_0(r_938_0),
		.io_in_valid_0(r_426_0),
		.io_out_a_0(_mesh_10_10_io_out_a_0),
		.io_out_c_0(_mesh_10_10_io_out_c_0),
		.io_out_b_0(_mesh_10_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_10_io_out_id_0),
		.io_out_last_0(_mesh_10_10_io_out_last_0),
		.io_out_valid_0(_mesh_10_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2565 == GlobalFiModInstNr[0]) || (2565 == GlobalFiModInstNr[1]) || (2565 == GlobalFiModInstNr[2]) || (2565 == GlobalFiModInstNr[3]))));
	Tile mesh_10_11(
		.clock(clock),
		.io_in_a_0(r_171_0),
		.io_in_b_0(b_186_0),
		.io_in_d_0(b_442_0),
		.io_in_control_0_dataflow(mesh_10_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_11_io_in_control_0_shift_b),
		.io_in_id_0(r_698_0),
		.io_in_last_0(r_954_0),
		.io_in_valid_0(r_442_0),
		.io_out_a_0(_mesh_10_11_io_out_a_0),
		.io_out_c_0(_mesh_10_11_io_out_c_0),
		.io_out_b_0(_mesh_10_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_11_io_out_id_0),
		.io_out_last_0(_mesh_10_11_io_out_last_0),
		.io_out_valid_0(_mesh_10_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2566 == GlobalFiModInstNr[0]) || (2566 == GlobalFiModInstNr[1]) || (2566 == GlobalFiModInstNr[2]) || (2566 == GlobalFiModInstNr[3]))));
	Tile mesh_10_12(
		.clock(clock),
		.io_in_a_0(r_172_0),
		.io_in_b_0(b_202_0),
		.io_in_d_0(b_458_0),
		.io_in_control_0_dataflow(mesh_10_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_12_io_in_control_0_shift_b),
		.io_in_id_0(r_714_0),
		.io_in_last_0(r_970_0),
		.io_in_valid_0(r_458_0),
		.io_out_a_0(_mesh_10_12_io_out_a_0),
		.io_out_c_0(_mesh_10_12_io_out_c_0),
		.io_out_b_0(_mesh_10_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_12_io_out_id_0),
		.io_out_last_0(_mesh_10_12_io_out_last_0),
		.io_out_valid_0(_mesh_10_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2567 == GlobalFiModInstNr[0]) || (2567 == GlobalFiModInstNr[1]) || (2567 == GlobalFiModInstNr[2]) || (2567 == GlobalFiModInstNr[3]))));
	Tile mesh_10_13(
		.clock(clock),
		.io_in_a_0(r_173_0),
		.io_in_b_0(b_218_0),
		.io_in_d_0(b_474_0),
		.io_in_control_0_dataflow(mesh_10_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_13_io_in_control_0_shift_b),
		.io_in_id_0(r_730_0),
		.io_in_last_0(r_986_0),
		.io_in_valid_0(r_474_0),
		.io_out_a_0(_mesh_10_13_io_out_a_0),
		.io_out_c_0(_mesh_10_13_io_out_c_0),
		.io_out_b_0(_mesh_10_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_13_io_out_id_0),
		.io_out_last_0(_mesh_10_13_io_out_last_0),
		.io_out_valid_0(_mesh_10_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2568 == GlobalFiModInstNr[0]) || (2568 == GlobalFiModInstNr[1]) || (2568 == GlobalFiModInstNr[2]) || (2568 == GlobalFiModInstNr[3]))));
	Tile mesh_10_14(
		.clock(clock),
		.io_in_a_0(r_174_0),
		.io_in_b_0(b_234_0),
		.io_in_d_0(b_490_0),
		.io_in_control_0_dataflow(mesh_10_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_14_io_in_control_0_shift_b),
		.io_in_id_0(r_746_0),
		.io_in_last_0(r_1002_0),
		.io_in_valid_0(r_490_0),
		.io_out_a_0(_mesh_10_14_io_out_a_0),
		.io_out_c_0(_mesh_10_14_io_out_c_0),
		.io_out_b_0(_mesh_10_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_14_io_out_id_0),
		.io_out_last_0(_mesh_10_14_io_out_last_0),
		.io_out_valid_0(_mesh_10_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2569 == GlobalFiModInstNr[0]) || (2569 == GlobalFiModInstNr[1]) || (2569 == GlobalFiModInstNr[2]) || (2569 == GlobalFiModInstNr[3]))));
	Tile mesh_10_15(
		.clock(clock),
		.io_in_a_0(r_175_0),
		.io_in_b_0(b_250_0),
		.io_in_d_0(b_506_0),
		.io_in_control_0_dataflow(mesh_10_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_15_io_in_control_0_shift_b),
		.io_in_id_0(r_762_0),
		.io_in_last_0(r_1018_0),
		.io_in_valid_0(r_506_0),
		.io_out_a_0(_mesh_10_15_io_out_a_0),
		.io_out_c_0(_mesh_10_15_io_out_c_0),
		.io_out_b_0(_mesh_10_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_15_io_out_id_0),
		.io_out_last_0(_mesh_10_15_io_out_last_0),
		.io_out_valid_0(_mesh_10_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2570 == GlobalFiModInstNr[0]) || (2570 == GlobalFiModInstNr[1]) || (2570 == GlobalFiModInstNr[2]) || (2570 == GlobalFiModInstNr[3]))));
	Tile mesh_11_0(
		.clock(clock),
		.io_in_a_0(r_176_0),
		.io_in_b_0(b_11_0),
		.io_in_d_0(b_267_0),
		.io_in_control_0_dataflow(mesh_11_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_0_io_in_control_0_shift_b),
		.io_in_id_0(r_523_0),
		.io_in_last_0(r_779_0),
		.io_in_valid_0(r_267_0),
		.io_out_a_0(_mesh_11_0_io_out_a_0),
		.io_out_c_0(_mesh_11_0_io_out_c_0),
		.io_out_b_0(_mesh_11_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_0_io_out_id_0),
		.io_out_last_0(_mesh_11_0_io_out_last_0),
		.io_out_valid_0(_mesh_11_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2571 == GlobalFiModInstNr[0]) || (2571 == GlobalFiModInstNr[1]) || (2571 == GlobalFiModInstNr[2]) || (2571 == GlobalFiModInstNr[3]))));
	Tile mesh_11_1(
		.clock(clock),
		.io_in_a_0(r_177_0),
		.io_in_b_0(b_27_0),
		.io_in_d_0(b_283_0),
		.io_in_control_0_dataflow(mesh_11_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_1_io_in_control_0_shift_b),
		.io_in_id_0(r_539_0),
		.io_in_last_0(r_795_0),
		.io_in_valid_0(r_283_0),
		.io_out_a_0(_mesh_11_1_io_out_a_0),
		.io_out_c_0(_mesh_11_1_io_out_c_0),
		.io_out_b_0(_mesh_11_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_1_io_out_id_0),
		.io_out_last_0(_mesh_11_1_io_out_last_0),
		.io_out_valid_0(_mesh_11_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2572 == GlobalFiModInstNr[0]) || (2572 == GlobalFiModInstNr[1]) || (2572 == GlobalFiModInstNr[2]) || (2572 == GlobalFiModInstNr[3]))));
	Tile mesh_11_2(
		.clock(clock),
		.io_in_a_0(r_178_0),
		.io_in_b_0(b_43_0),
		.io_in_d_0(b_299_0),
		.io_in_control_0_dataflow(mesh_11_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_2_io_in_control_0_shift_b),
		.io_in_id_0(r_555_0),
		.io_in_last_0(r_811_0),
		.io_in_valid_0(r_299_0),
		.io_out_a_0(_mesh_11_2_io_out_a_0),
		.io_out_c_0(_mesh_11_2_io_out_c_0),
		.io_out_b_0(_mesh_11_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_2_io_out_id_0),
		.io_out_last_0(_mesh_11_2_io_out_last_0),
		.io_out_valid_0(_mesh_11_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2573 == GlobalFiModInstNr[0]) || (2573 == GlobalFiModInstNr[1]) || (2573 == GlobalFiModInstNr[2]) || (2573 == GlobalFiModInstNr[3]))));
	Tile mesh_11_3(
		.clock(clock),
		.io_in_a_0(r_179_0),
		.io_in_b_0(b_59_0),
		.io_in_d_0(b_315_0),
		.io_in_control_0_dataflow(mesh_11_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_3_io_in_control_0_shift_b),
		.io_in_id_0(r_571_0),
		.io_in_last_0(r_827_0),
		.io_in_valid_0(r_315_0),
		.io_out_a_0(_mesh_11_3_io_out_a_0),
		.io_out_c_0(_mesh_11_3_io_out_c_0),
		.io_out_b_0(_mesh_11_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_3_io_out_id_0),
		.io_out_last_0(_mesh_11_3_io_out_last_0),
		.io_out_valid_0(_mesh_11_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2574 == GlobalFiModInstNr[0]) || (2574 == GlobalFiModInstNr[1]) || (2574 == GlobalFiModInstNr[2]) || (2574 == GlobalFiModInstNr[3]))));
	Tile mesh_11_4(
		.clock(clock),
		.io_in_a_0(r_180_0),
		.io_in_b_0(b_75_0),
		.io_in_d_0(b_331_0),
		.io_in_control_0_dataflow(mesh_11_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_4_io_in_control_0_shift_b),
		.io_in_id_0(r_587_0),
		.io_in_last_0(r_843_0),
		.io_in_valid_0(r_331_0),
		.io_out_a_0(_mesh_11_4_io_out_a_0),
		.io_out_c_0(_mesh_11_4_io_out_c_0),
		.io_out_b_0(_mesh_11_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_4_io_out_id_0),
		.io_out_last_0(_mesh_11_4_io_out_last_0),
		.io_out_valid_0(_mesh_11_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2575 == GlobalFiModInstNr[0]) || (2575 == GlobalFiModInstNr[1]) || (2575 == GlobalFiModInstNr[2]) || (2575 == GlobalFiModInstNr[3]))));
	Tile mesh_11_5(
		.clock(clock),
		.io_in_a_0(r_181_0),
		.io_in_b_0(b_91_0),
		.io_in_d_0(b_347_0),
		.io_in_control_0_dataflow(mesh_11_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_5_io_in_control_0_shift_b),
		.io_in_id_0(r_603_0),
		.io_in_last_0(r_859_0),
		.io_in_valid_0(r_347_0),
		.io_out_a_0(_mesh_11_5_io_out_a_0),
		.io_out_c_0(_mesh_11_5_io_out_c_0),
		.io_out_b_0(_mesh_11_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_5_io_out_id_0),
		.io_out_last_0(_mesh_11_5_io_out_last_0),
		.io_out_valid_0(_mesh_11_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2576 == GlobalFiModInstNr[0]) || (2576 == GlobalFiModInstNr[1]) || (2576 == GlobalFiModInstNr[2]) || (2576 == GlobalFiModInstNr[3]))));
	Tile mesh_11_6(
		.clock(clock),
		.io_in_a_0(r_182_0),
		.io_in_b_0(b_107_0),
		.io_in_d_0(b_363_0),
		.io_in_control_0_dataflow(mesh_11_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_6_io_in_control_0_shift_b),
		.io_in_id_0(r_619_0),
		.io_in_last_0(r_875_0),
		.io_in_valid_0(r_363_0),
		.io_out_a_0(_mesh_11_6_io_out_a_0),
		.io_out_c_0(_mesh_11_6_io_out_c_0),
		.io_out_b_0(_mesh_11_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_6_io_out_id_0),
		.io_out_last_0(_mesh_11_6_io_out_last_0),
		.io_out_valid_0(_mesh_11_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2577 == GlobalFiModInstNr[0]) || (2577 == GlobalFiModInstNr[1]) || (2577 == GlobalFiModInstNr[2]) || (2577 == GlobalFiModInstNr[3]))));
	Tile mesh_11_7(
		.clock(clock),
		.io_in_a_0(r_183_0),
		.io_in_b_0(b_123_0),
		.io_in_d_0(b_379_0),
		.io_in_control_0_dataflow(mesh_11_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_7_io_in_control_0_shift_b),
		.io_in_id_0(r_635_0),
		.io_in_last_0(r_891_0),
		.io_in_valid_0(r_379_0),
		.io_out_a_0(_mesh_11_7_io_out_a_0),
		.io_out_c_0(_mesh_11_7_io_out_c_0),
		.io_out_b_0(_mesh_11_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_7_io_out_id_0),
		.io_out_last_0(_mesh_11_7_io_out_last_0),
		.io_out_valid_0(_mesh_11_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2578 == GlobalFiModInstNr[0]) || (2578 == GlobalFiModInstNr[1]) || (2578 == GlobalFiModInstNr[2]) || (2578 == GlobalFiModInstNr[3]))));
	Tile mesh_11_8(
		.clock(clock),
		.io_in_a_0(r_184_0),
		.io_in_b_0(b_139_0),
		.io_in_d_0(b_395_0),
		.io_in_control_0_dataflow(mesh_11_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_8_io_in_control_0_shift_b),
		.io_in_id_0(r_651_0),
		.io_in_last_0(r_907_0),
		.io_in_valid_0(r_395_0),
		.io_out_a_0(_mesh_11_8_io_out_a_0),
		.io_out_c_0(_mesh_11_8_io_out_c_0),
		.io_out_b_0(_mesh_11_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_8_io_out_id_0),
		.io_out_last_0(_mesh_11_8_io_out_last_0),
		.io_out_valid_0(_mesh_11_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2579 == GlobalFiModInstNr[0]) || (2579 == GlobalFiModInstNr[1]) || (2579 == GlobalFiModInstNr[2]) || (2579 == GlobalFiModInstNr[3]))));
	Tile mesh_11_9(
		.clock(clock),
		.io_in_a_0(r_185_0),
		.io_in_b_0(b_155_0),
		.io_in_d_0(b_411_0),
		.io_in_control_0_dataflow(mesh_11_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_9_io_in_control_0_shift_b),
		.io_in_id_0(r_667_0),
		.io_in_last_0(r_923_0),
		.io_in_valid_0(r_411_0),
		.io_out_a_0(_mesh_11_9_io_out_a_0),
		.io_out_c_0(_mesh_11_9_io_out_c_0),
		.io_out_b_0(_mesh_11_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_9_io_out_id_0),
		.io_out_last_0(_mesh_11_9_io_out_last_0),
		.io_out_valid_0(_mesh_11_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2580 == GlobalFiModInstNr[0]) || (2580 == GlobalFiModInstNr[1]) || (2580 == GlobalFiModInstNr[2]) || (2580 == GlobalFiModInstNr[3]))));
	Tile mesh_11_10(
		.clock(clock),
		.io_in_a_0(r_186_0),
		.io_in_b_0(b_171_0),
		.io_in_d_0(b_427_0),
		.io_in_control_0_dataflow(mesh_11_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_10_io_in_control_0_shift_b),
		.io_in_id_0(r_683_0),
		.io_in_last_0(r_939_0),
		.io_in_valid_0(r_427_0),
		.io_out_a_0(_mesh_11_10_io_out_a_0),
		.io_out_c_0(_mesh_11_10_io_out_c_0),
		.io_out_b_0(_mesh_11_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_10_io_out_id_0),
		.io_out_last_0(_mesh_11_10_io_out_last_0),
		.io_out_valid_0(_mesh_11_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2581 == GlobalFiModInstNr[0]) || (2581 == GlobalFiModInstNr[1]) || (2581 == GlobalFiModInstNr[2]) || (2581 == GlobalFiModInstNr[3]))));
	Tile mesh_11_11(
		.clock(clock),
		.io_in_a_0(r_187_0),
		.io_in_b_0(b_187_0),
		.io_in_d_0(b_443_0),
		.io_in_control_0_dataflow(mesh_11_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_11_io_in_control_0_shift_b),
		.io_in_id_0(r_699_0),
		.io_in_last_0(r_955_0),
		.io_in_valid_0(r_443_0),
		.io_out_a_0(_mesh_11_11_io_out_a_0),
		.io_out_c_0(_mesh_11_11_io_out_c_0),
		.io_out_b_0(_mesh_11_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_11_io_out_id_0),
		.io_out_last_0(_mesh_11_11_io_out_last_0),
		.io_out_valid_0(_mesh_11_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2582 == GlobalFiModInstNr[0]) || (2582 == GlobalFiModInstNr[1]) || (2582 == GlobalFiModInstNr[2]) || (2582 == GlobalFiModInstNr[3]))));
	Tile mesh_11_12(
		.clock(clock),
		.io_in_a_0(r_188_0),
		.io_in_b_0(b_203_0),
		.io_in_d_0(b_459_0),
		.io_in_control_0_dataflow(mesh_11_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_12_io_in_control_0_shift_b),
		.io_in_id_0(r_715_0),
		.io_in_last_0(r_971_0),
		.io_in_valid_0(r_459_0),
		.io_out_a_0(_mesh_11_12_io_out_a_0),
		.io_out_c_0(_mesh_11_12_io_out_c_0),
		.io_out_b_0(_mesh_11_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_12_io_out_id_0),
		.io_out_last_0(_mesh_11_12_io_out_last_0),
		.io_out_valid_0(_mesh_11_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2583 == GlobalFiModInstNr[0]) || (2583 == GlobalFiModInstNr[1]) || (2583 == GlobalFiModInstNr[2]) || (2583 == GlobalFiModInstNr[3]))));
	Tile mesh_11_13(
		.clock(clock),
		.io_in_a_0(r_189_0),
		.io_in_b_0(b_219_0),
		.io_in_d_0(b_475_0),
		.io_in_control_0_dataflow(mesh_11_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_13_io_in_control_0_shift_b),
		.io_in_id_0(r_731_0),
		.io_in_last_0(r_987_0),
		.io_in_valid_0(r_475_0),
		.io_out_a_0(_mesh_11_13_io_out_a_0),
		.io_out_c_0(_mesh_11_13_io_out_c_0),
		.io_out_b_0(_mesh_11_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_13_io_out_id_0),
		.io_out_last_0(_mesh_11_13_io_out_last_0),
		.io_out_valid_0(_mesh_11_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2584 == GlobalFiModInstNr[0]) || (2584 == GlobalFiModInstNr[1]) || (2584 == GlobalFiModInstNr[2]) || (2584 == GlobalFiModInstNr[3]))));
	Tile mesh_11_14(
		.clock(clock),
		.io_in_a_0(r_190_0),
		.io_in_b_0(b_235_0),
		.io_in_d_0(b_491_0),
		.io_in_control_0_dataflow(mesh_11_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_14_io_in_control_0_shift_b),
		.io_in_id_0(r_747_0),
		.io_in_last_0(r_1003_0),
		.io_in_valid_0(r_491_0),
		.io_out_a_0(_mesh_11_14_io_out_a_0),
		.io_out_c_0(_mesh_11_14_io_out_c_0),
		.io_out_b_0(_mesh_11_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_14_io_out_id_0),
		.io_out_last_0(_mesh_11_14_io_out_last_0),
		.io_out_valid_0(_mesh_11_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2585 == GlobalFiModInstNr[0]) || (2585 == GlobalFiModInstNr[1]) || (2585 == GlobalFiModInstNr[2]) || (2585 == GlobalFiModInstNr[3]))));
	Tile mesh_11_15(
		.clock(clock),
		.io_in_a_0(r_191_0),
		.io_in_b_0(b_251_0),
		.io_in_d_0(b_507_0),
		.io_in_control_0_dataflow(mesh_11_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_15_io_in_control_0_shift_b),
		.io_in_id_0(r_763_0),
		.io_in_last_0(r_1019_0),
		.io_in_valid_0(r_507_0),
		.io_out_a_0(_mesh_11_15_io_out_a_0),
		.io_out_c_0(_mesh_11_15_io_out_c_0),
		.io_out_b_0(_mesh_11_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_15_io_out_id_0),
		.io_out_last_0(_mesh_11_15_io_out_last_0),
		.io_out_valid_0(_mesh_11_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2586 == GlobalFiModInstNr[0]) || (2586 == GlobalFiModInstNr[1]) || (2586 == GlobalFiModInstNr[2]) || (2586 == GlobalFiModInstNr[3]))));
	Tile mesh_12_0(
		.clock(clock),
		.io_in_a_0(r_192_0),
		.io_in_b_0(b_12_0),
		.io_in_d_0(b_268_0),
		.io_in_control_0_dataflow(mesh_12_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_0_io_in_control_0_shift_b),
		.io_in_id_0(r_524_0),
		.io_in_last_0(r_780_0),
		.io_in_valid_0(r_268_0),
		.io_out_a_0(_mesh_12_0_io_out_a_0),
		.io_out_c_0(_mesh_12_0_io_out_c_0),
		.io_out_b_0(_mesh_12_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_0_io_out_id_0),
		.io_out_last_0(_mesh_12_0_io_out_last_0),
		.io_out_valid_0(_mesh_12_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2587 == GlobalFiModInstNr[0]) || (2587 == GlobalFiModInstNr[1]) || (2587 == GlobalFiModInstNr[2]) || (2587 == GlobalFiModInstNr[3]))));
	Tile mesh_12_1(
		.clock(clock),
		.io_in_a_0(r_193_0),
		.io_in_b_0(b_28_0),
		.io_in_d_0(b_284_0),
		.io_in_control_0_dataflow(mesh_12_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_1_io_in_control_0_shift_b),
		.io_in_id_0(r_540_0),
		.io_in_last_0(r_796_0),
		.io_in_valid_0(r_284_0),
		.io_out_a_0(_mesh_12_1_io_out_a_0),
		.io_out_c_0(_mesh_12_1_io_out_c_0),
		.io_out_b_0(_mesh_12_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_1_io_out_id_0),
		.io_out_last_0(_mesh_12_1_io_out_last_0),
		.io_out_valid_0(_mesh_12_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2588 == GlobalFiModInstNr[0]) || (2588 == GlobalFiModInstNr[1]) || (2588 == GlobalFiModInstNr[2]) || (2588 == GlobalFiModInstNr[3]))));
	Tile mesh_12_2(
		.clock(clock),
		.io_in_a_0(r_194_0),
		.io_in_b_0(b_44_0),
		.io_in_d_0(b_300_0),
		.io_in_control_0_dataflow(mesh_12_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_2_io_in_control_0_shift_b),
		.io_in_id_0(r_556_0),
		.io_in_last_0(r_812_0),
		.io_in_valid_0(r_300_0),
		.io_out_a_0(_mesh_12_2_io_out_a_0),
		.io_out_c_0(_mesh_12_2_io_out_c_0),
		.io_out_b_0(_mesh_12_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_2_io_out_id_0),
		.io_out_last_0(_mesh_12_2_io_out_last_0),
		.io_out_valid_0(_mesh_12_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2589 == GlobalFiModInstNr[0]) || (2589 == GlobalFiModInstNr[1]) || (2589 == GlobalFiModInstNr[2]) || (2589 == GlobalFiModInstNr[3]))));
	Tile mesh_12_3(
		.clock(clock),
		.io_in_a_0(r_195_0),
		.io_in_b_0(b_60_0),
		.io_in_d_0(b_316_0),
		.io_in_control_0_dataflow(mesh_12_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_3_io_in_control_0_shift_b),
		.io_in_id_0(r_572_0),
		.io_in_last_0(r_828_0),
		.io_in_valid_0(r_316_0),
		.io_out_a_0(_mesh_12_3_io_out_a_0),
		.io_out_c_0(_mesh_12_3_io_out_c_0),
		.io_out_b_0(_mesh_12_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_3_io_out_id_0),
		.io_out_last_0(_mesh_12_3_io_out_last_0),
		.io_out_valid_0(_mesh_12_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2590 == GlobalFiModInstNr[0]) || (2590 == GlobalFiModInstNr[1]) || (2590 == GlobalFiModInstNr[2]) || (2590 == GlobalFiModInstNr[3]))));
	Tile mesh_12_4(
		.clock(clock),
		.io_in_a_0(r_196_0),
		.io_in_b_0(b_76_0),
		.io_in_d_0(b_332_0),
		.io_in_control_0_dataflow(mesh_12_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_4_io_in_control_0_shift_b),
		.io_in_id_0(r_588_0),
		.io_in_last_0(r_844_0),
		.io_in_valid_0(r_332_0),
		.io_out_a_0(_mesh_12_4_io_out_a_0),
		.io_out_c_0(_mesh_12_4_io_out_c_0),
		.io_out_b_0(_mesh_12_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_4_io_out_id_0),
		.io_out_last_0(_mesh_12_4_io_out_last_0),
		.io_out_valid_0(_mesh_12_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2591 == GlobalFiModInstNr[0]) || (2591 == GlobalFiModInstNr[1]) || (2591 == GlobalFiModInstNr[2]) || (2591 == GlobalFiModInstNr[3]))));
	Tile mesh_12_5(
		.clock(clock),
		.io_in_a_0(r_197_0),
		.io_in_b_0(b_92_0),
		.io_in_d_0(b_348_0),
		.io_in_control_0_dataflow(mesh_12_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_5_io_in_control_0_shift_b),
		.io_in_id_0(r_604_0),
		.io_in_last_0(r_860_0),
		.io_in_valid_0(r_348_0),
		.io_out_a_0(_mesh_12_5_io_out_a_0),
		.io_out_c_0(_mesh_12_5_io_out_c_0),
		.io_out_b_0(_mesh_12_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_5_io_out_id_0),
		.io_out_last_0(_mesh_12_5_io_out_last_0),
		.io_out_valid_0(_mesh_12_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2592 == GlobalFiModInstNr[0]) || (2592 == GlobalFiModInstNr[1]) || (2592 == GlobalFiModInstNr[2]) || (2592 == GlobalFiModInstNr[3]))));
	Tile mesh_12_6(
		.clock(clock),
		.io_in_a_0(r_198_0),
		.io_in_b_0(b_108_0),
		.io_in_d_0(b_364_0),
		.io_in_control_0_dataflow(mesh_12_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_6_io_in_control_0_shift_b),
		.io_in_id_0(r_620_0),
		.io_in_last_0(r_876_0),
		.io_in_valid_0(r_364_0),
		.io_out_a_0(_mesh_12_6_io_out_a_0),
		.io_out_c_0(_mesh_12_6_io_out_c_0),
		.io_out_b_0(_mesh_12_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_6_io_out_id_0),
		.io_out_last_0(_mesh_12_6_io_out_last_0),
		.io_out_valid_0(_mesh_12_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2593 == GlobalFiModInstNr[0]) || (2593 == GlobalFiModInstNr[1]) || (2593 == GlobalFiModInstNr[2]) || (2593 == GlobalFiModInstNr[3]))));
	Tile mesh_12_7(
		.clock(clock),
		.io_in_a_0(r_199_0),
		.io_in_b_0(b_124_0),
		.io_in_d_0(b_380_0),
		.io_in_control_0_dataflow(mesh_12_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_7_io_in_control_0_shift_b),
		.io_in_id_0(r_636_0),
		.io_in_last_0(r_892_0),
		.io_in_valid_0(r_380_0),
		.io_out_a_0(_mesh_12_7_io_out_a_0),
		.io_out_c_0(_mesh_12_7_io_out_c_0),
		.io_out_b_0(_mesh_12_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_7_io_out_id_0),
		.io_out_last_0(_mesh_12_7_io_out_last_0),
		.io_out_valid_0(_mesh_12_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2594 == GlobalFiModInstNr[0]) || (2594 == GlobalFiModInstNr[1]) || (2594 == GlobalFiModInstNr[2]) || (2594 == GlobalFiModInstNr[3]))));
	Tile mesh_12_8(
		.clock(clock),
		.io_in_a_0(r_200_0),
		.io_in_b_0(b_140_0),
		.io_in_d_0(b_396_0),
		.io_in_control_0_dataflow(mesh_12_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_8_io_in_control_0_shift_b),
		.io_in_id_0(r_652_0),
		.io_in_last_0(r_908_0),
		.io_in_valid_0(r_396_0),
		.io_out_a_0(_mesh_12_8_io_out_a_0),
		.io_out_c_0(_mesh_12_8_io_out_c_0),
		.io_out_b_0(_mesh_12_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_8_io_out_id_0),
		.io_out_last_0(_mesh_12_8_io_out_last_0),
		.io_out_valid_0(_mesh_12_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2595 == GlobalFiModInstNr[0]) || (2595 == GlobalFiModInstNr[1]) || (2595 == GlobalFiModInstNr[2]) || (2595 == GlobalFiModInstNr[3]))));
	Tile mesh_12_9(
		.clock(clock),
		.io_in_a_0(r_201_0),
		.io_in_b_0(b_156_0),
		.io_in_d_0(b_412_0),
		.io_in_control_0_dataflow(mesh_12_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_9_io_in_control_0_shift_b),
		.io_in_id_0(r_668_0),
		.io_in_last_0(r_924_0),
		.io_in_valid_0(r_412_0),
		.io_out_a_0(_mesh_12_9_io_out_a_0),
		.io_out_c_0(_mesh_12_9_io_out_c_0),
		.io_out_b_0(_mesh_12_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_9_io_out_id_0),
		.io_out_last_0(_mesh_12_9_io_out_last_0),
		.io_out_valid_0(_mesh_12_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2596 == GlobalFiModInstNr[0]) || (2596 == GlobalFiModInstNr[1]) || (2596 == GlobalFiModInstNr[2]) || (2596 == GlobalFiModInstNr[3]))));
	Tile mesh_12_10(
		.clock(clock),
		.io_in_a_0(r_202_0),
		.io_in_b_0(b_172_0),
		.io_in_d_0(b_428_0),
		.io_in_control_0_dataflow(mesh_12_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_10_io_in_control_0_shift_b),
		.io_in_id_0(r_684_0),
		.io_in_last_0(r_940_0),
		.io_in_valid_0(r_428_0),
		.io_out_a_0(_mesh_12_10_io_out_a_0),
		.io_out_c_0(_mesh_12_10_io_out_c_0),
		.io_out_b_0(_mesh_12_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_10_io_out_id_0),
		.io_out_last_0(_mesh_12_10_io_out_last_0),
		.io_out_valid_0(_mesh_12_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2597 == GlobalFiModInstNr[0]) || (2597 == GlobalFiModInstNr[1]) || (2597 == GlobalFiModInstNr[2]) || (2597 == GlobalFiModInstNr[3]))));
	Tile mesh_12_11(
		.clock(clock),
		.io_in_a_0(r_203_0),
		.io_in_b_0(b_188_0),
		.io_in_d_0(b_444_0),
		.io_in_control_0_dataflow(mesh_12_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_11_io_in_control_0_shift_b),
		.io_in_id_0(r_700_0),
		.io_in_last_0(r_956_0),
		.io_in_valid_0(r_444_0),
		.io_out_a_0(_mesh_12_11_io_out_a_0),
		.io_out_c_0(_mesh_12_11_io_out_c_0),
		.io_out_b_0(_mesh_12_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_11_io_out_id_0),
		.io_out_last_0(_mesh_12_11_io_out_last_0),
		.io_out_valid_0(_mesh_12_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2598 == GlobalFiModInstNr[0]) || (2598 == GlobalFiModInstNr[1]) || (2598 == GlobalFiModInstNr[2]) || (2598 == GlobalFiModInstNr[3]))));
	Tile mesh_12_12(
		.clock(clock),
		.io_in_a_0(r_204_0),
		.io_in_b_0(b_204_0),
		.io_in_d_0(b_460_0),
		.io_in_control_0_dataflow(mesh_12_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_12_io_in_control_0_shift_b),
		.io_in_id_0(r_716_0),
		.io_in_last_0(r_972_0),
		.io_in_valid_0(r_460_0),
		.io_out_a_0(_mesh_12_12_io_out_a_0),
		.io_out_c_0(_mesh_12_12_io_out_c_0),
		.io_out_b_0(_mesh_12_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_12_io_out_id_0),
		.io_out_last_0(_mesh_12_12_io_out_last_0),
		.io_out_valid_0(_mesh_12_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2599 == GlobalFiModInstNr[0]) || (2599 == GlobalFiModInstNr[1]) || (2599 == GlobalFiModInstNr[2]) || (2599 == GlobalFiModInstNr[3]))));
	Tile mesh_12_13(
		.clock(clock),
		.io_in_a_0(r_205_0),
		.io_in_b_0(b_220_0),
		.io_in_d_0(b_476_0),
		.io_in_control_0_dataflow(mesh_12_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_13_io_in_control_0_shift_b),
		.io_in_id_0(r_732_0),
		.io_in_last_0(r_988_0),
		.io_in_valid_0(r_476_0),
		.io_out_a_0(_mesh_12_13_io_out_a_0),
		.io_out_c_0(_mesh_12_13_io_out_c_0),
		.io_out_b_0(_mesh_12_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_13_io_out_id_0),
		.io_out_last_0(_mesh_12_13_io_out_last_0),
		.io_out_valid_0(_mesh_12_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2600 == GlobalFiModInstNr[0]) || (2600 == GlobalFiModInstNr[1]) || (2600 == GlobalFiModInstNr[2]) || (2600 == GlobalFiModInstNr[3]))));
	Tile mesh_12_14(
		.clock(clock),
		.io_in_a_0(r_206_0),
		.io_in_b_0(b_236_0),
		.io_in_d_0(b_492_0),
		.io_in_control_0_dataflow(mesh_12_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_14_io_in_control_0_shift_b),
		.io_in_id_0(r_748_0),
		.io_in_last_0(r_1004_0),
		.io_in_valid_0(r_492_0),
		.io_out_a_0(_mesh_12_14_io_out_a_0),
		.io_out_c_0(_mesh_12_14_io_out_c_0),
		.io_out_b_0(_mesh_12_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_14_io_out_id_0),
		.io_out_last_0(_mesh_12_14_io_out_last_0),
		.io_out_valid_0(_mesh_12_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2601 == GlobalFiModInstNr[0]) || (2601 == GlobalFiModInstNr[1]) || (2601 == GlobalFiModInstNr[2]) || (2601 == GlobalFiModInstNr[3]))));
	Tile mesh_12_15(
		.clock(clock),
		.io_in_a_0(r_207_0),
		.io_in_b_0(b_252_0),
		.io_in_d_0(b_508_0),
		.io_in_control_0_dataflow(mesh_12_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_15_io_in_control_0_shift_b),
		.io_in_id_0(r_764_0),
		.io_in_last_0(r_1020_0),
		.io_in_valid_0(r_508_0),
		.io_out_a_0(_mesh_12_15_io_out_a_0),
		.io_out_c_0(_mesh_12_15_io_out_c_0),
		.io_out_b_0(_mesh_12_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_15_io_out_id_0),
		.io_out_last_0(_mesh_12_15_io_out_last_0),
		.io_out_valid_0(_mesh_12_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2602 == GlobalFiModInstNr[0]) || (2602 == GlobalFiModInstNr[1]) || (2602 == GlobalFiModInstNr[2]) || (2602 == GlobalFiModInstNr[3]))));
	Tile mesh_13_0(
		.clock(clock),
		.io_in_a_0(r_208_0),
		.io_in_b_0(b_13_0),
		.io_in_d_0(b_269_0),
		.io_in_control_0_dataflow(mesh_13_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_0_io_in_control_0_shift_b),
		.io_in_id_0(r_525_0),
		.io_in_last_0(r_781_0),
		.io_in_valid_0(r_269_0),
		.io_out_a_0(_mesh_13_0_io_out_a_0),
		.io_out_c_0(_mesh_13_0_io_out_c_0),
		.io_out_b_0(_mesh_13_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_0_io_out_id_0),
		.io_out_last_0(_mesh_13_0_io_out_last_0),
		.io_out_valid_0(_mesh_13_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2603 == GlobalFiModInstNr[0]) || (2603 == GlobalFiModInstNr[1]) || (2603 == GlobalFiModInstNr[2]) || (2603 == GlobalFiModInstNr[3]))));
	Tile mesh_13_1(
		.clock(clock),
		.io_in_a_0(r_209_0),
		.io_in_b_0(b_29_0),
		.io_in_d_0(b_285_0),
		.io_in_control_0_dataflow(mesh_13_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_1_io_in_control_0_shift_b),
		.io_in_id_0(r_541_0),
		.io_in_last_0(r_797_0),
		.io_in_valid_0(r_285_0),
		.io_out_a_0(_mesh_13_1_io_out_a_0),
		.io_out_c_0(_mesh_13_1_io_out_c_0),
		.io_out_b_0(_mesh_13_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_1_io_out_id_0),
		.io_out_last_0(_mesh_13_1_io_out_last_0),
		.io_out_valid_0(_mesh_13_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2604 == GlobalFiModInstNr[0]) || (2604 == GlobalFiModInstNr[1]) || (2604 == GlobalFiModInstNr[2]) || (2604 == GlobalFiModInstNr[3]))));
	Tile mesh_13_2(
		.clock(clock),
		.io_in_a_0(r_210_0),
		.io_in_b_0(b_45_0),
		.io_in_d_0(b_301_0),
		.io_in_control_0_dataflow(mesh_13_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_2_io_in_control_0_shift_b),
		.io_in_id_0(r_557_0),
		.io_in_last_0(r_813_0),
		.io_in_valid_0(r_301_0),
		.io_out_a_0(_mesh_13_2_io_out_a_0),
		.io_out_c_0(_mesh_13_2_io_out_c_0),
		.io_out_b_0(_mesh_13_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_2_io_out_id_0),
		.io_out_last_0(_mesh_13_2_io_out_last_0),
		.io_out_valid_0(_mesh_13_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2605 == GlobalFiModInstNr[0]) || (2605 == GlobalFiModInstNr[1]) || (2605 == GlobalFiModInstNr[2]) || (2605 == GlobalFiModInstNr[3]))));
	Tile mesh_13_3(
		.clock(clock),
		.io_in_a_0(r_211_0),
		.io_in_b_0(b_61_0),
		.io_in_d_0(b_317_0),
		.io_in_control_0_dataflow(mesh_13_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_3_io_in_control_0_shift_b),
		.io_in_id_0(r_573_0),
		.io_in_last_0(r_829_0),
		.io_in_valid_0(r_317_0),
		.io_out_a_0(_mesh_13_3_io_out_a_0),
		.io_out_c_0(_mesh_13_3_io_out_c_0),
		.io_out_b_0(_mesh_13_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_3_io_out_id_0),
		.io_out_last_0(_mesh_13_3_io_out_last_0),
		.io_out_valid_0(_mesh_13_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2606 == GlobalFiModInstNr[0]) || (2606 == GlobalFiModInstNr[1]) || (2606 == GlobalFiModInstNr[2]) || (2606 == GlobalFiModInstNr[3]))));
	Tile mesh_13_4(
		.clock(clock),
		.io_in_a_0(r_212_0),
		.io_in_b_0(b_77_0),
		.io_in_d_0(b_333_0),
		.io_in_control_0_dataflow(mesh_13_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_4_io_in_control_0_shift_b),
		.io_in_id_0(r_589_0),
		.io_in_last_0(r_845_0),
		.io_in_valid_0(r_333_0),
		.io_out_a_0(_mesh_13_4_io_out_a_0),
		.io_out_c_0(_mesh_13_4_io_out_c_0),
		.io_out_b_0(_mesh_13_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_4_io_out_id_0),
		.io_out_last_0(_mesh_13_4_io_out_last_0),
		.io_out_valid_0(_mesh_13_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2607 == GlobalFiModInstNr[0]) || (2607 == GlobalFiModInstNr[1]) || (2607 == GlobalFiModInstNr[2]) || (2607 == GlobalFiModInstNr[3]))));
	Tile mesh_13_5(
		.clock(clock),
		.io_in_a_0(r_213_0),
		.io_in_b_0(b_93_0),
		.io_in_d_0(b_349_0),
		.io_in_control_0_dataflow(mesh_13_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_5_io_in_control_0_shift_b),
		.io_in_id_0(r_605_0),
		.io_in_last_0(r_861_0),
		.io_in_valid_0(r_349_0),
		.io_out_a_0(_mesh_13_5_io_out_a_0),
		.io_out_c_0(_mesh_13_5_io_out_c_0),
		.io_out_b_0(_mesh_13_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_5_io_out_id_0),
		.io_out_last_0(_mesh_13_5_io_out_last_0),
		.io_out_valid_0(_mesh_13_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2608 == GlobalFiModInstNr[0]) || (2608 == GlobalFiModInstNr[1]) || (2608 == GlobalFiModInstNr[2]) || (2608 == GlobalFiModInstNr[3]))));
	Tile mesh_13_6(
		.clock(clock),
		.io_in_a_0(r_214_0),
		.io_in_b_0(b_109_0),
		.io_in_d_0(b_365_0),
		.io_in_control_0_dataflow(mesh_13_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_6_io_in_control_0_shift_b),
		.io_in_id_0(r_621_0),
		.io_in_last_0(r_877_0),
		.io_in_valid_0(r_365_0),
		.io_out_a_0(_mesh_13_6_io_out_a_0),
		.io_out_c_0(_mesh_13_6_io_out_c_0),
		.io_out_b_0(_mesh_13_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_6_io_out_id_0),
		.io_out_last_0(_mesh_13_6_io_out_last_0),
		.io_out_valid_0(_mesh_13_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2609 == GlobalFiModInstNr[0]) || (2609 == GlobalFiModInstNr[1]) || (2609 == GlobalFiModInstNr[2]) || (2609 == GlobalFiModInstNr[3]))));
	Tile mesh_13_7(
		.clock(clock),
		.io_in_a_0(r_215_0),
		.io_in_b_0(b_125_0),
		.io_in_d_0(b_381_0),
		.io_in_control_0_dataflow(mesh_13_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_7_io_in_control_0_shift_b),
		.io_in_id_0(r_637_0),
		.io_in_last_0(r_893_0),
		.io_in_valid_0(r_381_0),
		.io_out_a_0(_mesh_13_7_io_out_a_0),
		.io_out_c_0(_mesh_13_7_io_out_c_0),
		.io_out_b_0(_mesh_13_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_7_io_out_id_0),
		.io_out_last_0(_mesh_13_7_io_out_last_0),
		.io_out_valid_0(_mesh_13_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2610 == GlobalFiModInstNr[0]) || (2610 == GlobalFiModInstNr[1]) || (2610 == GlobalFiModInstNr[2]) || (2610 == GlobalFiModInstNr[3]))));
	Tile mesh_13_8(
		.clock(clock),
		.io_in_a_0(r_216_0),
		.io_in_b_0(b_141_0),
		.io_in_d_0(b_397_0),
		.io_in_control_0_dataflow(mesh_13_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_8_io_in_control_0_shift_b),
		.io_in_id_0(r_653_0),
		.io_in_last_0(r_909_0),
		.io_in_valid_0(r_397_0),
		.io_out_a_0(_mesh_13_8_io_out_a_0),
		.io_out_c_0(_mesh_13_8_io_out_c_0),
		.io_out_b_0(_mesh_13_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_8_io_out_id_0),
		.io_out_last_0(_mesh_13_8_io_out_last_0),
		.io_out_valid_0(_mesh_13_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2611 == GlobalFiModInstNr[0]) || (2611 == GlobalFiModInstNr[1]) || (2611 == GlobalFiModInstNr[2]) || (2611 == GlobalFiModInstNr[3]))));
	Tile mesh_13_9(
		.clock(clock),
		.io_in_a_0(r_217_0),
		.io_in_b_0(b_157_0),
		.io_in_d_0(b_413_0),
		.io_in_control_0_dataflow(mesh_13_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_9_io_in_control_0_shift_b),
		.io_in_id_0(r_669_0),
		.io_in_last_0(r_925_0),
		.io_in_valid_0(r_413_0),
		.io_out_a_0(_mesh_13_9_io_out_a_0),
		.io_out_c_0(_mesh_13_9_io_out_c_0),
		.io_out_b_0(_mesh_13_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_9_io_out_id_0),
		.io_out_last_0(_mesh_13_9_io_out_last_0),
		.io_out_valid_0(_mesh_13_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2612 == GlobalFiModInstNr[0]) || (2612 == GlobalFiModInstNr[1]) || (2612 == GlobalFiModInstNr[2]) || (2612 == GlobalFiModInstNr[3]))));
	Tile mesh_13_10(
		.clock(clock),
		.io_in_a_0(r_218_0),
		.io_in_b_0(b_173_0),
		.io_in_d_0(b_429_0),
		.io_in_control_0_dataflow(mesh_13_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_10_io_in_control_0_shift_b),
		.io_in_id_0(r_685_0),
		.io_in_last_0(r_941_0),
		.io_in_valid_0(r_429_0),
		.io_out_a_0(_mesh_13_10_io_out_a_0),
		.io_out_c_0(_mesh_13_10_io_out_c_0),
		.io_out_b_0(_mesh_13_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_10_io_out_id_0),
		.io_out_last_0(_mesh_13_10_io_out_last_0),
		.io_out_valid_0(_mesh_13_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2613 == GlobalFiModInstNr[0]) || (2613 == GlobalFiModInstNr[1]) || (2613 == GlobalFiModInstNr[2]) || (2613 == GlobalFiModInstNr[3]))));
	Tile mesh_13_11(
		.clock(clock),
		.io_in_a_0(r_219_0),
		.io_in_b_0(b_189_0),
		.io_in_d_0(b_445_0),
		.io_in_control_0_dataflow(mesh_13_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_11_io_in_control_0_shift_b),
		.io_in_id_0(r_701_0),
		.io_in_last_0(r_957_0),
		.io_in_valid_0(r_445_0),
		.io_out_a_0(_mesh_13_11_io_out_a_0),
		.io_out_c_0(_mesh_13_11_io_out_c_0),
		.io_out_b_0(_mesh_13_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_11_io_out_id_0),
		.io_out_last_0(_mesh_13_11_io_out_last_0),
		.io_out_valid_0(_mesh_13_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2614 == GlobalFiModInstNr[0]) || (2614 == GlobalFiModInstNr[1]) || (2614 == GlobalFiModInstNr[2]) || (2614 == GlobalFiModInstNr[3]))));
	Tile mesh_13_12(
		.clock(clock),
		.io_in_a_0(r_220_0),
		.io_in_b_0(b_205_0),
		.io_in_d_0(b_461_0),
		.io_in_control_0_dataflow(mesh_13_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_12_io_in_control_0_shift_b),
		.io_in_id_0(r_717_0),
		.io_in_last_0(r_973_0),
		.io_in_valid_0(r_461_0),
		.io_out_a_0(_mesh_13_12_io_out_a_0),
		.io_out_c_0(_mesh_13_12_io_out_c_0),
		.io_out_b_0(_mesh_13_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_12_io_out_id_0),
		.io_out_last_0(_mesh_13_12_io_out_last_0),
		.io_out_valid_0(_mesh_13_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2615 == GlobalFiModInstNr[0]) || (2615 == GlobalFiModInstNr[1]) || (2615 == GlobalFiModInstNr[2]) || (2615 == GlobalFiModInstNr[3]))));
	Tile mesh_13_13(
		.clock(clock),
		.io_in_a_0(r_221_0),
		.io_in_b_0(b_221_0),
		.io_in_d_0(b_477_0),
		.io_in_control_0_dataflow(mesh_13_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_13_io_in_control_0_shift_b),
		.io_in_id_0(r_733_0),
		.io_in_last_0(r_989_0),
		.io_in_valid_0(r_477_0),
		.io_out_a_0(_mesh_13_13_io_out_a_0),
		.io_out_c_0(_mesh_13_13_io_out_c_0),
		.io_out_b_0(_mesh_13_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_13_io_out_id_0),
		.io_out_last_0(_mesh_13_13_io_out_last_0),
		.io_out_valid_0(_mesh_13_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2616 == GlobalFiModInstNr[0]) || (2616 == GlobalFiModInstNr[1]) || (2616 == GlobalFiModInstNr[2]) || (2616 == GlobalFiModInstNr[3]))));
	Tile mesh_13_14(
		.clock(clock),
		.io_in_a_0(r_222_0),
		.io_in_b_0(b_237_0),
		.io_in_d_0(b_493_0),
		.io_in_control_0_dataflow(mesh_13_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_14_io_in_control_0_shift_b),
		.io_in_id_0(r_749_0),
		.io_in_last_0(r_1005_0),
		.io_in_valid_0(r_493_0),
		.io_out_a_0(_mesh_13_14_io_out_a_0),
		.io_out_c_0(_mesh_13_14_io_out_c_0),
		.io_out_b_0(_mesh_13_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_14_io_out_id_0),
		.io_out_last_0(_mesh_13_14_io_out_last_0),
		.io_out_valid_0(_mesh_13_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2617 == GlobalFiModInstNr[0]) || (2617 == GlobalFiModInstNr[1]) || (2617 == GlobalFiModInstNr[2]) || (2617 == GlobalFiModInstNr[3]))));
	Tile mesh_13_15(
		.clock(clock),
		.io_in_a_0(r_223_0),
		.io_in_b_0(b_253_0),
		.io_in_d_0(b_509_0),
		.io_in_control_0_dataflow(mesh_13_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_15_io_in_control_0_shift_b),
		.io_in_id_0(r_765_0),
		.io_in_last_0(r_1021_0),
		.io_in_valid_0(r_509_0),
		.io_out_a_0(_mesh_13_15_io_out_a_0),
		.io_out_c_0(_mesh_13_15_io_out_c_0),
		.io_out_b_0(_mesh_13_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_15_io_out_id_0),
		.io_out_last_0(_mesh_13_15_io_out_last_0),
		.io_out_valid_0(_mesh_13_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2618 == GlobalFiModInstNr[0]) || (2618 == GlobalFiModInstNr[1]) || (2618 == GlobalFiModInstNr[2]) || (2618 == GlobalFiModInstNr[3]))));
	Tile mesh_14_0(
		.clock(clock),
		.io_in_a_0(r_224_0),
		.io_in_b_0(b_14_0),
		.io_in_d_0(b_270_0),
		.io_in_control_0_dataflow(mesh_14_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_0_io_in_control_0_shift_b),
		.io_in_id_0(r_526_0),
		.io_in_last_0(r_782_0),
		.io_in_valid_0(r_270_0),
		.io_out_a_0(_mesh_14_0_io_out_a_0),
		.io_out_c_0(_mesh_14_0_io_out_c_0),
		.io_out_b_0(_mesh_14_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_0_io_out_id_0),
		.io_out_last_0(_mesh_14_0_io_out_last_0),
		.io_out_valid_0(_mesh_14_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2619 == GlobalFiModInstNr[0]) || (2619 == GlobalFiModInstNr[1]) || (2619 == GlobalFiModInstNr[2]) || (2619 == GlobalFiModInstNr[3]))));
	Tile mesh_14_1(
		.clock(clock),
		.io_in_a_0(r_225_0),
		.io_in_b_0(b_30_0),
		.io_in_d_0(b_286_0),
		.io_in_control_0_dataflow(mesh_14_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_1_io_in_control_0_shift_b),
		.io_in_id_0(r_542_0),
		.io_in_last_0(r_798_0),
		.io_in_valid_0(r_286_0),
		.io_out_a_0(_mesh_14_1_io_out_a_0),
		.io_out_c_0(_mesh_14_1_io_out_c_0),
		.io_out_b_0(_mesh_14_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_1_io_out_id_0),
		.io_out_last_0(_mesh_14_1_io_out_last_0),
		.io_out_valid_0(_mesh_14_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2620 == GlobalFiModInstNr[0]) || (2620 == GlobalFiModInstNr[1]) || (2620 == GlobalFiModInstNr[2]) || (2620 == GlobalFiModInstNr[3]))));
	Tile mesh_14_2(
		.clock(clock),
		.io_in_a_0(r_226_0),
		.io_in_b_0(b_46_0),
		.io_in_d_0(b_302_0),
		.io_in_control_0_dataflow(mesh_14_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_2_io_in_control_0_shift_b),
		.io_in_id_0(r_558_0),
		.io_in_last_0(r_814_0),
		.io_in_valid_0(r_302_0),
		.io_out_a_0(_mesh_14_2_io_out_a_0),
		.io_out_c_0(_mesh_14_2_io_out_c_0),
		.io_out_b_0(_mesh_14_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_2_io_out_id_0),
		.io_out_last_0(_mesh_14_2_io_out_last_0),
		.io_out_valid_0(_mesh_14_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2621 == GlobalFiModInstNr[0]) || (2621 == GlobalFiModInstNr[1]) || (2621 == GlobalFiModInstNr[2]) || (2621 == GlobalFiModInstNr[3]))));
	Tile mesh_14_3(
		.clock(clock),
		.io_in_a_0(r_227_0),
		.io_in_b_0(b_62_0),
		.io_in_d_0(b_318_0),
		.io_in_control_0_dataflow(mesh_14_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_3_io_in_control_0_shift_b),
		.io_in_id_0(r_574_0),
		.io_in_last_0(r_830_0),
		.io_in_valid_0(r_318_0),
		.io_out_a_0(_mesh_14_3_io_out_a_0),
		.io_out_c_0(_mesh_14_3_io_out_c_0),
		.io_out_b_0(_mesh_14_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_3_io_out_id_0),
		.io_out_last_0(_mesh_14_3_io_out_last_0),
		.io_out_valid_0(_mesh_14_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2622 == GlobalFiModInstNr[0]) || (2622 == GlobalFiModInstNr[1]) || (2622 == GlobalFiModInstNr[2]) || (2622 == GlobalFiModInstNr[3]))));
	Tile mesh_14_4(
		.clock(clock),
		.io_in_a_0(r_228_0),
		.io_in_b_0(b_78_0),
		.io_in_d_0(b_334_0),
		.io_in_control_0_dataflow(mesh_14_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_4_io_in_control_0_shift_b),
		.io_in_id_0(r_590_0),
		.io_in_last_0(r_846_0),
		.io_in_valid_0(r_334_0),
		.io_out_a_0(_mesh_14_4_io_out_a_0),
		.io_out_c_0(_mesh_14_4_io_out_c_0),
		.io_out_b_0(_mesh_14_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_4_io_out_id_0),
		.io_out_last_0(_mesh_14_4_io_out_last_0),
		.io_out_valid_0(_mesh_14_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2623 == GlobalFiModInstNr[0]) || (2623 == GlobalFiModInstNr[1]) || (2623 == GlobalFiModInstNr[2]) || (2623 == GlobalFiModInstNr[3]))));
	Tile mesh_14_5(
		.clock(clock),
		.io_in_a_0(r_229_0),
		.io_in_b_0(b_94_0),
		.io_in_d_0(b_350_0),
		.io_in_control_0_dataflow(mesh_14_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_5_io_in_control_0_shift_b),
		.io_in_id_0(r_606_0),
		.io_in_last_0(r_862_0),
		.io_in_valid_0(r_350_0),
		.io_out_a_0(_mesh_14_5_io_out_a_0),
		.io_out_c_0(_mesh_14_5_io_out_c_0),
		.io_out_b_0(_mesh_14_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_5_io_out_id_0),
		.io_out_last_0(_mesh_14_5_io_out_last_0),
		.io_out_valid_0(_mesh_14_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2624 == GlobalFiModInstNr[0]) || (2624 == GlobalFiModInstNr[1]) || (2624 == GlobalFiModInstNr[2]) || (2624 == GlobalFiModInstNr[3]))));
	Tile mesh_14_6(
		.clock(clock),
		.io_in_a_0(r_230_0),
		.io_in_b_0(b_110_0),
		.io_in_d_0(b_366_0),
		.io_in_control_0_dataflow(mesh_14_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_6_io_in_control_0_shift_b),
		.io_in_id_0(r_622_0),
		.io_in_last_0(r_878_0),
		.io_in_valid_0(r_366_0),
		.io_out_a_0(_mesh_14_6_io_out_a_0),
		.io_out_c_0(_mesh_14_6_io_out_c_0),
		.io_out_b_0(_mesh_14_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_6_io_out_id_0),
		.io_out_last_0(_mesh_14_6_io_out_last_0),
		.io_out_valid_0(_mesh_14_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2625 == GlobalFiModInstNr[0]) || (2625 == GlobalFiModInstNr[1]) || (2625 == GlobalFiModInstNr[2]) || (2625 == GlobalFiModInstNr[3]))));
	Tile mesh_14_7(
		.clock(clock),
		.io_in_a_0(r_231_0),
		.io_in_b_0(b_126_0),
		.io_in_d_0(b_382_0),
		.io_in_control_0_dataflow(mesh_14_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_7_io_in_control_0_shift_b),
		.io_in_id_0(r_638_0),
		.io_in_last_0(r_894_0),
		.io_in_valid_0(r_382_0),
		.io_out_a_0(_mesh_14_7_io_out_a_0),
		.io_out_c_0(_mesh_14_7_io_out_c_0),
		.io_out_b_0(_mesh_14_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_7_io_out_id_0),
		.io_out_last_0(_mesh_14_7_io_out_last_0),
		.io_out_valid_0(_mesh_14_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2626 == GlobalFiModInstNr[0]) || (2626 == GlobalFiModInstNr[1]) || (2626 == GlobalFiModInstNr[2]) || (2626 == GlobalFiModInstNr[3]))));
	Tile mesh_14_8(
		.clock(clock),
		.io_in_a_0(r_232_0),
		.io_in_b_0(b_142_0),
		.io_in_d_0(b_398_0),
		.io_in_control_0_dataflow(mesh_14_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_8_io_in_control_0_shift_b),
		.io_in_id_0(r_654_0),
		.io_in_last_0(r_910_0),
		.io_in_valid_0(r_398_0),
		.io_out_a_0(_mesh_14_8_io_out_a_0),
		.io_out_c_0(_mesh_14_8_io_out_c_0),
		.io_out_b_0(_mesh_14_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_8_io_out_id_0),
		.io_out_last_0(_mesh_14_8_io_out_last_0),
		.io_out_valid_0(_mesh_14_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2627 == GlobalFiModInstNr[0]) || (2627 == GlobalFiModInstNr[1]) || (2627 == GlobalFiModInstNr[2]) || (2627 == GlobalFiModInstNr[3]))));
	Tile mesh_14_9(
		.clock(clock),
		.io_in_a_0(r_233_0),
		.io_in_b_0(b_158_0),
		.io_in_d_0(b_414_0),
		.io_in_control_0_dataflow(mesh_14_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_9_io_in_control_0_shift_b),
		.io_in_id_0(r_670_0),
		.io_in_last_0(r_926_0),
		.io_in_valid_0(r_414_0),
		.io_out_a_0(_mesh_14_9_io_out_a_0),
		.io_out_c_0(_mesh_14_9_io_out_c_0),
		.io_out_b_0(_mesh_14_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_9_io_out_id_0),
		.io_out_last_0(_mesh_14_9_io_out_last_0),
		.io_out_valid_0(_mesh_14_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2628 == GlobalFiModInstNr[0]) || (2628 == GlobalFiModInstNr[1]) || (2628 == GlobalFiModInstNr[2]) || (2628 == GlobalFiModInstNr[3]))));
	Tile mesh_14_10(
		.clock(clock),
		.io_in_a_0(r_234_0),
		.io_in_b_0(b_174_0),
		.io_in_d_0(b_430_0),
		.io_in_control_0_dataflow(mesh_14_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_10_io_in_control_0_shift_b),
		.io_in_id_0(r_686_0),
		.io_in_last_0(r_942_0),
		.io_in_valid_0(r_430_0),
		.io_out_a_0(_mesh_14_10_io_out_a_0),
		.io_out_c_0(_mesh_14_10_io_out_c_0),
		.io_out_b_0(_mesh_14_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_10_io_out_id_0),
		.io_out_last_0(_mesh_14_10_io_out_last_0),
		.io_out_valid_0(_mesh_14_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2629 == GlobalFiModInstNr[0]) || (2629 == GlobalFiModInstNr[1]) || (2629 == GlobalFiModInstNr[2]) || (2629 == GlobalFiModInstNr[3]))));
	Tile mesh_14_11(
		.clock(clock),
		.io_in_a_0(r_235_0),
		.io_in_b_0(b_190_0),
		.io_in_d_0(b_446_0),
		.io_in_control_0_dataflow(mesh_14_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_11_io_in_control_0_shift_b),
		.io_in_id_0(r_702_0),
		.io_in_last_0(r_958_0),
		.io_in_valid_0(r_446_0),
		.io_out_a_0(_mesh_14_11_io_out_a_0),
		.io_out_c_0(_mesh_14_11_io_out_c_0),
		.io_out_b_0(_mesh_14_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_11_io_out_id_0),
		.io_out_last_0(_mesh_14_11_io_out_last_0),
		.io_out_valid_0(_mesh_14_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2630 == GlobalFiModInstNr[0]) || (2630 == GlobalFiModInstNr[1]) || (2630 == GlobalFiModInstNr[2]) || (2630 == GlobalFiModInstNr[3]))));
	Tile mesh_14_12(
		.clock(clock),
		.io_in_a_0(r_236_0),
		.io_in_b_0(b_206_0),
		.io_in_d_0(b_462_0),
		.io_in_control_0_dataflow(mesh_14_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_12_io_in_control_0_shift_b),
		.io_in_id_0(r_718_0),
		.io_in_last_0(r_974_0),
		.io_in_valid_0(r_462_0),
		.io_out_a_0(_mesh_14_12_io_out_a_0),
		.io_out_c_0(_mesh_14_12_io_out_c_0),
		.io_out_b_0(_mesh_14_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_12_io_out_id_0),
		.io_out_last_0(_mesh_14_12_io_out_last_0),
		.io_out_valid_0(_mesh_14_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2631 == GlobalFiModInstNr[0]) || (2631 == GlobalFiModInstNr[1]) || (2631 == GlobalFiModInstNr[2]) || (2631 == GlobalFiModInstNr[3]))));
	Tile mesh_14_13(
		.clock(clock),
		.io_in_a_0(r_237_0),
		.io_in_b_0(b_222_0),
		.io_in_d_0(b_478_0),
		.io_in_control_0_dataflow(mesh_14_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_13_io_in_control_0_shift_b),
		.io_in_id_0(r_734_0),
		.io_in_last_0(r_990_0),
		.io_in_valid_0(r_478_0),
		.io_out_a_0(_mesh_14_13_io_out_a_0),
		.io_out_c_0(_mesh_14_13_io_out_c_0),
		.io_out_b_0(_mesh_14_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_13_io_out_id_0),
		.io_out_last_0(_mesh_14_13_io_out_last_0),
		.io_out_valid_0(_mesh_14_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2632 == GlobalFiModInstNr[0]) || (2632 == GlobalFiModInstNr[1]) || (2632 == GlobalFiModInstNr[2]) || (2632 == GlobalFiModInstNr[3]))));
	Tile mesh_14_14(
		.clock(clock),
		.io_in_a_0(r_238_0),
		.io_in_b_0(b_238_0),
		.io_in_d_0(b_494_0),
		.io_in_control_0_dataflow(mesh_14_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_14_io_in_control_0_shift_b),
		.io_in_id_0(r_750_0),
		.io_in_last_0(r_1006_0),
		.io_in_valid_0(r_494_0),
		.io_out_a_0(_mesh_14_14_io_out_a_0),
		.io_out_c_0(_mesh_14_14_io_out_c_0),
		.io_out_b_0(_mesh_14_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_14_io_out_id_0),
		.io_out_last_0(_mesh_14_14_io_out_last_0),
		.io_out_valid_0(_mesh_14_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2633 == GlobalFiModInstNr[0]) || (2633 == GlobalFiModInstNr[1]) || (2633 == GlobalFiModInstNr[2]) || (2633 == GlobalFiModInstNr[3]))));
	Tile mesh_14_15(
		.clock(clock),
		.io_in_a_0(r_239_0),
		.io_in_b_0(b_254_0),
		.io_in_d_0(b_510_0),
		.io_in_control_0_dataflow(mesh_14_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_15_io_in_control_0_shift_b),
		.io_in_id_0(r_766_0),
		.io_in_last_0(r_1022_0),
		.io_in_valid_0(r_510_0),
		.io_out_a_0(_mesh_14_15_io_out_a_0),
		.io_out_c_0(_mesh_14_15_io_out_c_0),
		.io_out_b_0(_mesh_14_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_15_io_out_id_0),
		.io_out_last_0(_mesh_14_15_io_out_last_0),
		.io_out_valid_0(_mesh_14_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2634 == GlobalFiModInstNr[0]) || (2634 == GlobalFiModInstNr[1]) || (2634 == GlobalFiModInstNr[2]) || (2634 == GlobalFiModInstNr[3]))));
	Tile mesh_15_0(
		.clock(clock),
		.io_in_a_0(r_240_0),
		.io_in_b_0(b_15_0),
		.io_in_d_0(b_271_0),
		.io_in_control_0_dataflow(mesh_15_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_0_io_in_control_0_shift_b),
		.io_in_id_0(r_527_0),
		.io_in_last_0(r_783_0),
		.io_in_valid_0(r_271_0),
		.io_out_a_0(_mesh_15_0_io_out_a_0),
		.io_out_c_0(_mesh_15_0_io_out_c_0),
		.io_out_b_0(_mesh_15_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_0_io_out_id_0),
		.io_out_last_0(_mesh_15_0_io_out_last_0),
		.io_out_valid_0(_mesh_15_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2635 == GlobalFiModInstNr[0]) || (2635 == GlobalFiModInstNr[1]) || (2635 == GlobalFiModInstNr[2]) || (2635 == GlobalFiModInstNr[3]))));
	Tile mesh_15_1(
		.clock(clock),
		.io_in_a_0(r_241_0),
		.io_in_b_0(b_31_0),
		.io_in_d_0(b_287_0),
		.io_in_control_0_dataflow(mesh_15_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_1_io_in_control_0_shift_b),
		.io_in_id_0(r_543_0),
		.io_in_last_0(r_799_0),
		.io_in_valid_0(r_287_0),
		.io_out_a_0(_mesh_15_1_io_out_a_0),
		.io_out_c_0(_mesh_15_1_io_out_c_0),
		.io_out_b_0(_mesh_15_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_1_io_out_id_0),
		.io_out_last_0(_mesh_15_1_io_out_last_0),
		.io_out_valid_0(_mesh_15_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2636 == GlobalFiModInstNr[0]) || (2636 == GlobalFiModInstNr[1]) || (2636 == GlobalFiModInstNr[2]) || (2636 == GlobalFiModInstNr[3]))));
	Tile mesh_15_2(
		.clock(clock),
		.io_in_a_0(r_242_0),
		.io_in_b_0(b_47_0),
		.io_in_d_0(b_303_0),
		.io_in_control_0_dataflow(mesh_15_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_2_io_in_control_0_shift_b),
		.io_in_id_0(r_559_0),
		.io_in_last_0(r_815_0),
		.io_in_valid_0(r_303_0),
		.io_out_a_0(_mesh_15_2_io_out_a_0),
		.io_out_c_0(_mesh_15_2_io_out_c_0),
		.io_out_b_0(_mesh_15_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_2_io_out_id_0),
		.io_out_last_0(_mesh_15_2_io_out_last_0),
		.io_out_valid_0(_mesh_15_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2637 == GlobalFiModInstNr[0]) || (2637 == GlobalFiModInstNr[1]) || (2637 == GlobalFiModInstNr[2]) || (2637 == GlobalFiModInstNr[3]))));
	Tile mesh_15_3(
		.clock(clock),
		.io_in_a_0(r_243_0),
		.io_in_b_0(b_63_0),
		.io_in_d_0(b_319_0),
		.io_in_control_0_dataflow(mesh_15_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_3_io_in_control_0_shift_b),
		.io_in_id_0(r_575_0),
		.io_in_last_0(r_831_0),
		.io_in_valid_0(r_319_0),
		.io_out_a_0(_mesh_15_3_io_out_a_0),
		.io_out_c_0(_mesh_15_3_io_out_c_0),
		.io_out_b_0(_mesh_15_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_3_io_out_id_0),
		.io_out_last_0(_mesh_15_3_io_out_last_0),
		.io_out_valid_0(_mesh_15_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2638 == GlobalFiModInstNr[0]) || (2638 == GlobalFiModInstNr[1]) || (2638 == GlobalFiModInstNr[2]) || (2638 == GlobalFiModInstNr[3]))));
	Tile mesh_15_4(
		.clock(clock),
		.io_in_a_0(r_244_0),
		.io_in_b_0(b_79_0),
		.io_in_d_0(b_335_0),
		.io_in_control_0_dataflow(mesh_15_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_4_io_in_control_0_shift_b),
		.io_in_id_0(r_591_0),
		.io_in_last_0(r_847_0),
		.io_in_valid_0(r_335_0),
		.io_out_a_0(_mesh_15_4_io_out_a_0),
		.io_out_c_0(_mesh_15_4_io_out_c_0),
		.io_out_b_0(_mesh_15_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_4_io_out_id_0),
		.io_out_last_0(_mesh_15_4_io_out_last_0),
		.io_out_valid_0(_mesh_15_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2639 == GlobalFiModInstNr[0]) || (2639 == GlobalFiModInstNr[1]) || (2639 == GlobalFiModInstNr[2]) || (2639 == GlobalFiModInstNr[3]))));
	Tile mesh_15_5(
		.clock(clock),
		.io_in_a_0(r_245_0),
		.io_in_b_0(b_95_0),
		.io_in_d_0(b_351_0),
		.io_in_control_0_dataflow(mesh_15_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_5_io_in_control_0_shift_b),
		.io_in_id_0(r_607_0),
		.io_in_last_0(r_863_0),
		.io_in_valid_0(r_351_0),
		.io_out_a_0(_mesh_15_5_io_out_a_0),
		.io_out_c_0(_mesh_15_5_io_out_c_0),
		.io_out_b_0(_mesh_15_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_5_io_out_id_0),
		.io_out_last_0(_mesh_15_5_io_out_last_0),
		.io_out_valid_0(_mesh_15_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2640 == GlobalFiModInstNr[0]) || (2640 == GlobalFiModInstNr[1]) || (2640 == GlobalFiModInstNr[2]) || (2640 == GlobalFiModInstNr[3]))));
	Tile mesh_15_6(
		.clock(clock),
		.io_in_a_0(r_246_0),
		.io_in_b_0(b_111_0),
		.io_in_d_0(b_367_0),
		.io_in_control_0_dataflow(mesh_15_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_6_io_in_control_0_shift_b),
		.io_in_id_0(r_623_0),
		.io_in_last_0(r_879_0),
		.io_in_valid_0(r_367_0),
		.io_out_a_0(_mesh_15_6_io_out_a_0),
		.io_out_c_0(_mesh_15_6_io_out_c_0),
		.io_out_b_0(_mesh_15_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_6_io_out_id_0),
		.io_out_last_0(_mesh_15_6_io_out_last_0),
		.io_out_valid_0(_mesh_15_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2641 == GlobalFiModInstNr[0]) || (2641 == GlobalFiModInstNr[1]) || (2641 == GlobalFiModInstNr[2]) || (2641 == GlobalFiModInstNr[3]))));
	Tile mesh_15_7(
		.clock(clock),
		.io_in_a_0(r_247_0),
		.io_in_b_0(b_127_0),
		.io_in_d_0(b_383_0),
		.io_in_control_0_dataflow(mesh_15_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_7_io_in_control_0_shift_b),
		.io_in_id_0(r_639_0),
		.io_in_last_0(r_895_0),
		.io_in_valid_0(r_383_0),
		.io_out_a_0(_mesh_15_7_io_out_a_0),
		.io_out_c_0(_mesh_15_7_io_out_c_0),
		.io_out_b_0(_mesh_15_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_7_io_out_id_0),
		.io_out_last_0(_mesh_15_7_io_out_last_0),
		.io_out_valid_0(_mesh_15_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2642 == GlobalFiModInstNr[0]) || (2642 == GlobalFiModInstNr[1]) || (2642 == GlobalFiModInstNr[2]) || (2642 == GlobalFiModInstNr[3]))));
	Tile mesh_15_8(
		.clock(clock),
		.io_in_a_0(r_248_0),
		.io_in_b_0(b_143_0),
		.io_in_d_0(b_399_0),
		.io_in_control_0_dataflow(mesh_15_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_8_io_in_control_0_shift_b),
		.io_in_id_0(r_655_0),
		.io_in_last_0(r_911_0),
		.io_in_valid_0(r_399_0),
		.io_out_a_0(_mesh_15_8_io_out_a_0),
		.io_out_c_0(_mesh_15_8_io_out_c_0),
		.io_out_b_0(_mesh_15_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_8_io_out_id_0),
		.io_out_last_0(_mesh_15_8_io_out_last_0),
		.io_out_valid_0(_mesh_15_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2643 == GlobalFiModInstNr[0]) || (2643 == GlobalFiModInstNr[1]) || (2643 == GlobalFiModInstNr[2]) || (2643 == GlobalFiModInstNr[3]))));
	Tile mesh_15_9(
		.clock(clock),
		.io_in_a_0(r_249_0),
		.io_in_b_0(b_159_0),
		.io_in_d_0(b_415_0),
		.io_in_control_0_dataflow(mesh_15_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_9_io_in_control_0_shift_b),
		.io_in_id_0(r_671_0),
		.io_in_last_0(r_927_0),
		.io_in_valid_0(r_415_0),
		.io_out_a_0(_mesh_15_9_io_out_a_0),
		.io_out_c_0(_mesh_15_9_io_out_c_0),
		.io_out_b_0(_mesh_15_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_9_io_out_id_0),
		.io_out_last_0(_mesh_15_9_io_out_last_0),
		.io_out_valid_0(_mesh_15_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2644 == GlobalFiModInstNr[0]) || (2644 == GlobalFiModInstNr[1]) || (2644 == GlobalFiModInstNr[2]) || (2644 == GlobalFiModInstNr[3]))));
	Tile mesh_15_10(
		.clock(clock),
		.io_in_a_0(r_250_0),
		.io_in_b_0(b_175_0),
		.io_in_d_0(b_431_0),
		.io_in_control_0_dataflow(mesh_15_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_10_io_in_control_0_shift_b),
		.io_in_id_0(r_687_0),
		.io_in_last_0(r_943_0),
		.io_in_valid_0(r_431_0),
		.io_out_a_0(_mesh_15_10_io_out_a_0),
		.io_out_c_0(_mesh_15_10_io_out_c_0),
		.io_out_b_0(_mesh_15_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_10_io_out_id_0),
		.io_out_last_0(_mesh_15_10_io_out_last_0),
		.io_out_valid_0(_mesh_15_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2645 == GlobalFiModInstNr[0]) || (2645 == GlobalFiModInstNr[1]) || (2645 == GlobalFiModInstNr[2]) || (2645 == GlobalFiModInstNr[3]))));
	Tile mesh_15_11(
		.clock(clock),
		.io_in_a_0(r_251_0),
		.io_in_b_0(b_191_0),
		.io_in_d_0(b_447_0),
		.io_in_control_0_dataflow(mesh_15_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_11_io_in_control_0_shift_b),
		.io_in_id_0(r_703_0),
		.io_in_last_0(r_959_0),
		.io_in_valid_0(r_447_0),
		.io_out_a_0(_mesh_15_11_io_out_a_0),
		.io_out_c_0(_mesh_15_11_io_out_c_0),
		.io_out_b_0(_mesh_15_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_11_io_out_id_0),
		.io_out_last_0(_mesh_15_11_io_out_last_0),
		.io_out_valid_0(_mesh_15_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2646 == GlobalFiModInstNr[0]) || (2646 == GlobalFiModInstNr[1]) || (2646 == GlobalFiModInstNr[2]) || (2646 == GlobalFiModInstNr[3]))));
	Tile mesh_15_12(
		.clock(clock),
		.io_in_a_0(r_252_0),
		.io_in_b_0(b_207_0),
		.io_in_d_0(b_463_0),
		.io_in_control_0_dataflow(mesh_15_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_12_io_in_control_0_shift_b),
		.io_in_id_0(r_719_0),
		.io_in_last_0(r_975_0),
		.io_in_valid_0(r_463_0),
		.io_out_a_0(_mesh_15_12_io_out_a_0),
		.io_out_c_0(_mesh_15_12_io_out_c_0),
		.io_out_b_0(_mesh_15_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_12_io_out_id_0),
		.io_out_last_0(_mesh_15_12_io_out_last_0),
		.io_out_valid_0(_mesh_15_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2647 == GlobalFiModInstNr[0]) || (2647 == GlobalFiModInstNr[1]) || (2647 == GlobalFiModInstNr[2]) || (2647 == GlobalFiModInstNr[3]))));
	Tile mesh_15_13(
		.clock(clock),
		.io_in_a_0(r_253_0),
		.io_in_b_0(b_223_0),
		.io_in_d_0(b_479_0),
		.io_in_control_0_dataflow(mesh_15_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_13_io_in_control_0_shift_b),
		.io_in_id_0(r_735_0),
		.io_in_last_0(r_991_0),
		.io_in_valid_0(r_479_0),
		.io_out_a_0(_mesh_15_13_io_out_a_0),
		.io_out_c_0(_mesh_15_13_io_out_c_0),
		.io_out_b_0(_mesh_15_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_13_io_out_id_0),
		.io_out_last_0(_mesh_15_13_io_out_last_0),
		.io_out_valid_0(_mesh_15_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2648 == GlobalFiModInstNr[0]) || (2648 == GlobalFiModInstNr[1]) || (2648 == GlobalFiModInstNr[2]) || (2648 == GlobalFiModInstNr[3]))));
	Tile mesh_15_14(
		.clock(clock),
		.io_in_a_0(r_254_0),
		.io_in_b_0(b_239_0),
		.io_in_d_0(b_495_0),
		.io_in_control_0_dataflow(mesh_15_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_14_io_in_control_0_shift_b),
		.io_in_id_0(r_751_0),
		.io_in_last_0(r_1007_0),
		.io_in_valid_0(r_495_0),
		.io_out_a_0(_mesh_15_14_io_out_a_0),
		.io_out_c_0(_mesh_15_14_io_out_c_0),
		.io_out_b_0(_mesh_15_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_14_io_out_id_0),
		.io_out_last_0(_mesh_15_14_io_out_last_0),
		.io_out_valid_0(_mesh_15_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2649 == GlobalFiModInstNr[0]) || (2649 == GlobalFiModInstNr[1]) || (2649 == GlobalFiModInstNr[2]) || (2649 == GlobalFiModInstNr[3]))));
	Tile mesh_15_15(
		.clock(clock),
		.io_in_a_0(r_255_0),
		.io_in_b_0(b_255_0),
		.io_in_d_0(b_511_0),
		.io_in_control_0_dataflow(mesh_15_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_15_io_in_control_0_shift_b),
		.io_in_id_0(r_767_0),
		.io_in_last_0(r_1023_0),
		.io_in_valid_0(r_511_0),
		.io_out_a_0(_mesh_15_15_io_out_a_0),
		.io_out_c_0(_mesh_15_15_io_out_c_0),
		.io_out_b_0(_mesh_15_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_15_io_out_id_0),
		.io_out_last_0(_mesh_15_15_io_out_last_0),
		.io_out_valid_0(_mesh_15_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((2650 == GlobalFiModInstNr[0]) || (2650 == GlobalFiModInstNr[1]) || (2650 == GlobalFiModInstNr[2]) || (2650 == GlobalFiModInstNr[3]))));
	assign io_out_b_0_0 =( r_1024_0) ^ ((fiEnable && (2357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_1_0 =( r_1030_0) ^ ((fiEnable && (2358 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_2_0 =( r_1036_0) ^ ((fiEnable && (2359 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_3_0 =( r_1042_0) ^ ((fiEnable && (2360 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_4_0 =( r_1048_0) ^ ((fiEnable && (2361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_5_0 =( r_1054_0) ^ ((fiEnable && (2362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_6_0 =( r_1060_0) ^ ((fiEnable && (2363 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_7_0 =( r_1066_0) ^ ((fiEnable && (2364 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_8_0 =( r_1072_0) ^ ((fiEnable && (2365 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_9_0 =( r_1078_0) ^ ((fiEnable && (2366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_10_0 =( r_1084_0) ^ ((fiEnable && (2367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_11_0 =( r_1090_0) ^ ((fiEnable && (2368 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_12_0 =( r_1096_0) ^ ((fiEnable && (2369 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_13_0 =( r_1102_0) ^ ((fiEnable && (2370 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_14_0 =( r_1108_0) ^ ((fiEnable && (2371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_15_0 =( r_1114_0) ^ ((fiEnable && (2372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_0_0 =( r_1025_0) ^ ((fiEnable && (2373 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_1_0 =( r_1031_0) ^ ((fiEnable && (2374 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_2_0 =( r_1037_0) ^ ((fiEnable && (2375 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_3_0 =( r_1043_0) ^ ((fiEnable && (2376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_4_0 =( r_1049_0) ^ ((fiEnable && (2377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_5_0 =( r_1055_0) ^ ((fiEnable && (2378 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_6_0 =( r_1061_0) ^ ((fiEnable && (2379 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_7_0 =( r_1067_0) ^ ((fiEnable && (2380 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_8_0 =( r_1073_0) ^ ((fiEnable && (2381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_9_0 =( r_1079_0) ^ ((fiEnable && (2382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_10_0 =( r_1085_0) ^ ((fiEnable && (2383 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_11_0 =( r_1091_0) ^ ((fiEnable && (2384 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_12_0 =( r_1097_0) ^ ((fiEnable && (2385 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_13_0 =( r_1103_0) ^ ((fiEnable && (2386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_14_0 =( r_1109_0) ^ ((fiEnable && (2387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_15_0 =( r_1115_0) ^ ((fiEnable && (2388 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_valid_0_0 =( r_1026_0) ^ ((fiEnable && (2389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_0_0_dataflow =( r_1027_0_dataflow) ^ ((fiEnable && (2390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_id_0_0 =( r_1028_0) ^ ((fiEnable && (2391 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last_0_0 =( r_1029_0) ^ ((fiEnable && (2392 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
endmodule