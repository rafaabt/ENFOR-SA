module MacUnit (
	io_in_a,
	io_in_b,
	io_in_c,
	io_out_d
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_c;
	output logic [31:0] io_out_d;
	assign io_out_d =( (io_in_a * io_in_b) + io_in_c) ^ ((fiEnable && (2 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
endmodule
module PE_16 (
	clock,
	io_in_a,
	io_in_b,
	io_in_d,
	io_in_control_dataflow,
	io_in_control_propagate,
	io_in_control_shift,
	io_in_id,
	io_in_last,
	io_in_valid,
	io_out_a,
	io_out_b,
	io_out_c,
	io_out_control_dataflow,
	io_out_control_propagate,
	io_out_control_shift,
	io_out_id,
	io_out_last,
	io_out_valid
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_d;
	input io_in_control_dataflow;
	input io_in_control_propagate;
	input [4:0] io_in_control_shift;
	input [2:0] io_in_id;
	input io_in_last;
	input io_in_valid;
	output logic [31:0] io_out_a;
	output logic [31:0] io_out_b;
	output logic [31:0] io_out_c;
	output logic io_out_control_dataflow;
	output logic io_out_control_propagate;
	output logic [4:0] io_out_control_shift;
	output logic [2:0] io_out_id;
	output logic io_out_last;
	output logic io_out_valid;
	wire [31:0] _mac_unit_io_out_d;
	reg [31:0] c1;
	reg [31:0] c2;
	reg last_s;
	wire [4:0] shift_offset = (last_s != io_in_control_propagate ? io_in_control_shift : 5'h00);
	wire [31:0] _GEN = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_3 = $signed($signed(c1) >>> _GEN);
	wire [31:0] _GEN_0 = {27'h0000000, shift_offset};
	wire [31:0] _io_out_c_T = $signed($signed(c1) >>> _GEN_0);
	wire [31:0] _GEN_1 = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_8 = $signed($signed(c2) >>> _GEN_1);
	wire [31:0] _io_out_c_T_11 = $signed($signed(c2) >>> _GEN_0);
	always @(posedge clock)
		if (io_in_valid) begin
			if (io_in_control_propagate) begin
				c1 <=( io_in_d) ^ ((fiEnable && (3 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( _mac_unit_io_out_d) ^ ((fiEnable && (4 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			end
			else begin
				c1 <=( _mac_unit_io_out_d) ^ ((fiEnable && (5 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( io_in_d) ^ ((fiEnable && (6 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			end
			last_s <=( io_in_control_propagate) ^ ((fiEnable && (7 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
		end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	MacUnit mac_unit(
		.io_in_a(io_in_a),
		.io_in_b(io_in_b),
		.io_in_c((io_in_control_propagate ? c2 : c1)),
		.io_out_d(_mac_unit_io_out_d)
	,
    .fiEnable(fiEnable && ((185 == Mesh.GlobalFiModInstNr[0]) || (185 == Mesh.GlobalFiModInstNr[1]) || (185 == Mesh.GlobalFiModInstNr[2]) || (185 == Mesh.GlobalFiModInstNr[3]))));
    
	assign io_out_a =( io_in_a) ^ ((fiEnable && (8 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b =( io_in_b) ^ ((fiEnable && (9 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c =( (io_in_control_propagate ? _io_out_c_T + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_3[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c1 & ((32'h00000001 << _GEN) - 32'h00000001)) | _io_out_c_T[0])} : _io_out_c_T_11 + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_8[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c2 & ((32'h00000001 << _GEN_1) - 32'h00000001)) | _io_out_c_T_11[0])})) ^ ((fiEnable && (10 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_control_dataflow =( io_in_control_dataflow) ^ ((fiEnable && (11 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_propagate =( io_in_control_propagate) ^ ((fiEnable && (12 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_shift =( io_in_control_shift) ^ ((fiEnable && (13 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[4:0] : {5{1'b0}});
	assign io_out_id =( io_in_id) ^ ((fiEnable && (14 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last =( io_in_last) ^ ((fiEnable && (15 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_valid =( io_in_valid) ^ ((fiEnable && (16 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
endmodule
module Tile (
	clock,
	io_in_a_0,
	io_in_b_0,
	io_in_d_0,
	io_in_control_0_dataflow,
	io_in_control_0_propagate,
	io_in_control_0_shift,
	io_in_id_0,
	io_in_last_0,
	io_in_valid_0,
	io_out_a_0,
	io_out_c_0,
	io_out_b_0,
	io_out_control_0_dataflow,
	io_out_control_0_propagate,
	io_out_control_0_shift,
	io_out_id_0,
	io_out_last_0,
	io_out_valid_0
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a_0;
	input [31:0] io_in_b_0;
	input [31:0] io_in_d_0;
	input io_in_control_0_dataflow;
	input io_in_control_0_propagate;
	input [4:0] io_in_control_0_shift;
	input [2:0] io_in_id_0;
	input io_in_last_0;
	input io_in_valid_0;
	output logic [31:0] io_out_a_0;
	output logic [31:0] io_out_c_0;
	output logic [31:0] io_out_b_0;
	output logic io_out_control_0_dataflow;
	output logic io_out_control_0_propagate;
	output logic [4:0] io_out_control_0_shift;
	output logic [2:0] io_out_id_0;
	output logic io_out_last_0;
	output logic io_out_valid_0;
	PE_16 tile_0_0(
		.clock(clock),
		.io_in_a(io_in_a_0),
		.io_in_b(io_in_b_0),
		.io_in_d(io_in_d_0),
		.io_in_control_dataflow(io_in_control_0_dataflow),
		.io_in_control_propagate(io_in_control_0_propagate),
		.io_in_control_shift(io_in_control_0_shift),
		.io_in_id(io_in_id_0),
		.io_in_last(io_in_last_0),
		.io_in_valid(io_in_valid_0),
		.io_out_a(io_out_a_0),
		.io_out_b(io_out_b_0),
		.io_out_c(io_out_c_0),
		.io_out_control_dataflow(io_out_control_0_dataflow),
		.io_out_control_propagate(io_out_control_0_propagate),
		.io_out_control_shift(io_out_control_0_shift),
		.io_out_id(io_out_id_0),
		.io_out_last(io_out_last_0),
		.io_out_valid(io_out_valid_0)
	,
    .fiEnable(fiEnable && ((186 == Mesh.GlobalFiModInstNr[0]) || (186 == Mesh.GlobalFiModInstNr[1]) || (186 == Mesh.GlobalFiModInstNr[2]) || (186 == Mesh.GlobalFiModInstNr[3]))));
endmodule



module Mesh (
	clock,
	io_in_a_0_0,
	io_in_a_1_0,
	io_in_a_2_0,
	io_in_a_3_0,
	io_in_b_0_0,
	io_in_b_1_0,
	io_in_b_2_0,
	io_in_b_3_0,
	io_in_d_0_0,
	io_in_d_1_0,
	io_in_d_2_0,
	io_in_d_3_0,
	io_in_control_0_0_dataflow,
	io_in_control_0_0_propagate,
	io_in_control_0_0_shift,
	io_in_control_1_0_dataflow,
	io_in_control_1_0_propagate,
	io_in_control_1_0_shift,
	io_in_control_2_0_dataflow,
	io_in_control_2_0_propagate,
	io_in_control_2_0_shift,
	io_in_control_3_0_dataflow,
	io_in_control_3_0_propagate,
	io_in_control_3_0_shift,
	io_in_id_0_0,
	io_in_id_1_0,
	io_in_id_2_0,
	io_in_id_3_0,
	io_in_last_0_0,
	io_in_last_1_0,
	io_in_last_2_0,
	io_in_last_3_0,
	io_in_valid_0_0,
	io_in_valid_1_0,
	io_in_valid_2_0,
	io_in_valid_3_0,
	io_out_b_0_0,
	io_out_b_1_0,
	io_out_b_2_0,
	io_out_b_3_0,
	io_out_c_0_0,
	io_out_c_1_0,
	io_out_c_2_0,
	io_out_c_3_0,
	io_out_valid_0_0,
	io_out_control_0_0_dataflow,
	io_out_id_0_0,
	io_out_last_0_0
, GlobalFiSignal, GlobalFiNumber, GlobalFiModInstNr);
input GlobalFiSignal;
wire [31:0] GlobalFiSignal;
input GlobalFiNumber;
wire [31:0] GlobalFiNumber;
input GlobalFiModInstNr;
wire [15:0] GlobalFiModInstNr[4];
wire fiEnable;
assign fiEnable = (1 == GlobalFiModInstNr[0]) || (1 == GlobalFiModInstNr[1]) || (1 == GlobalFiModInstNr[2]) || (1 == GlobalFiModInstNr[3]);

	input clock;
	input [31:0] io_in_a_0_0;
	input [31:0] io_in_a_1_0;
	input [31:0] io_in_a_2_0;
	input [31:0] io_in_a_3_0;
	input [31:0] io_in_b_0_0;
	input [31:0] io_in_b_1_0;
	input [31:0] io_in_b_2_0;
	input [31:0] io_in_b_3_0;
	input [31:0] io_in_d_0_0;
	input [31:0] io_in_d_1_0;
	input [31:0] io_in_d_2_0;
	input [31:0] io_in_d_3_0;
	input io_in_control_0_0_dataflow;
	input io_in_control_0_0_propagate;
	input [4:0] io_in_control_0_0_shift;
	input io_in_control_1_0_dataflow;
	input io_in_control_1_0_propagate;
	input [4:0] io_in_control_1_0_shift;
	input io_in_control_2_0_dataflow;
	input io_in_control_2_0_propagate;
	input [4:0] io_in_control_2_0_shift;
	input io_in_control_3_0_dataflow;
	input io_in_control_3_0_propagate;
	input [4:0] io_in_control_3_0_shift;
	input [2:0] io_in_id_0_0;
	input [2:0] io_in_id_1_0;
	input [2:0] io_in_id_2_0;
	input [2:0] io_in_id_3_0;
	input io_in_last_0_0;
	input io_in_last_1_0;
	input io_in_last_2_0;
	input io_in_last_3_0;
	input io_in_valid_0_0;
	input io_in_valid_1_0;
	input io_in_valid_2_0;
	input io_in_valid_3_0;
	output logic [31:0] io_out_b_0_0;
	output logic [31:0] io_out_b_1_0;
	output logic [31:0] io_out_b_2_0;
	output logic [31:0] io_out_b_3_0;
	output logic [31:0] io_out_c_0_0;
	output logic [31:0] io_out_c_1_0;
	output logic [31:0] io_out_c_2_0;
	output logic [31:0] io_out_c_3_0;
	output logic io_out_valid_0_0;
	output logic io_out_control_0_0_dataflow;
	output logic [2:0] io_out_id_0_0;
	output logic io_out_last_0_0;
	wire [31:0] _mesh_3_3_io_out_a_0;
	wire [31:0] _mesh_3_3_io_out_c_0;
	wire [31:0] _mesh_3_3_io_out_b_0;
	wire _mesh_3_3_io_out_control_0_dataflow;
	wire _mesh_3_3_io_out_control_0_propagate;
	wire [4:0] _mesh_3_3_io_out_control_0_shift;
	wire [2:0] _mesh_3_3_io_out_id_0;
	wire _mesh_3_3_io_out_last_0;
	wire _mesh_3_3_io_out_valid_0;
	wire [31:0] _mesh_3_2_io_out_a_0;
	wire [31:0] _mesh_3_2_io_out_c_0;
	wire [31:0] _mesh_3_2_io_out_b_0;
	wire _mesh_3_2_io_out_control_0_dataflow;
	wire _mesh_3_2_io_out_control_0_propagate;
	wire [4:0] _mesh_3_2_io_out_control_0_shift;
	wire [2:0] _mesh_3_2_io_out_id_0;
	wire _mesh_3_2_io_out_last_0;
	wire _mesh_3_2_io_out_valid_0;
	wire [31:0] _mesh_3_1_io_out_a_0;
	wire [31:0] _mesh_3_1_io_out_c_0;
	wire [31:0] _mesh_3_1_io_out_b_0;
	wire _mesh_3_1_io_out_control_0_dataflow;
	wire _mesh_3_1_io_out_control_0_propagate;
	wire [4:0] _mesh_3_1_io_out_control_0_shift;
	wire [2:0] _mesh_3_1_io_out_id_0;
	wire _mesh_3_1_io_out_last_0;
	wire _mesh_3_1_io_out_valid_0;
	wire [31:0] _mesh_3_0_io_out_a_0;
	wire [31:0] _mesh_3_0_io_out_c_0;
	wire [31:0] _mesh_3_0_io_out_b_0;
	wire _mesh_3_0_io_out_control_0_dataflow;
	wire _mesh_3_0_io_out_control_0_propagate;
	wire [4:0] _mesh_3_0_io_out_control_0_shift;
	wire [2:0] _mesh_3_0_io_out_id_0;
	wire _mesh_3_0_io_out_last_0;
	wire _mesh_3_0_io_out_valid_0;
	wire [31:0] _mesh_2_3_io_out_a_0;
	wire [31:0] _mesh_2_3_io_out_c_0;
	wire [31:0] _mesh_2_3_io_out_b_0;
	wire _mesh_2_3_io_out_control_0_dataflow;
	wire _mesh_2_3_io_out_control_0_propagate;
	wire [4:0] _mesh_2_3_io_out_control_0_shift;
	wire [2:0] _mesh_2_3_io_out_id_0;
	wire _mesh_2_3_io_out_last_0;
	wire _mesh_2_3_io_out_valid_0;
	wire [31:0] _mesh_2_2_io_out_a_0;
	wire [31:0] _mesh_2_2_io_out_c_0;
	wire [31:0] _mesh_2_2_io_out_b_0;
	wire _mesh_2_2_io_out_control_0_dataflow;
	wire _mesh_2_2_io_out_control_0_propagate;
	wire [4:0] _mesh_2_2_io_out_control_0_shift;
	wire [2:0] _mesh_2_2_io_out_id_0;
	wire _mesh_2_2_io_out_last_0;
	wire _mesh_2_2_io_out_valid_0;
	wire [31:0] _mesh_2_1_io_out_a_0;
	wire [31:0] _mesh_2_1_io_out_c_0;
	wire [31:0] _mesh_2_1_io_out_b_0;
	wire _mesh_2_1_io_out_control_0_dataflow;
	wire _mesh_2_1_io_out_control_0_propagate;
	wire [4:0] _mesh_2_1_io_out_control_0_shift;
	wire [2:0] _mesh_2_1_io_out_id_0;
	wire _mesh_2_1_io_out_last_0;
	wire _mesh_2_1_io_out_valid_0;
	wire [31:0] _mesh_2_0_io_out_a_0;
	wire [31:0] _mesh_2_0_io_out_c_0;
	wire [31:0] _mesh_2_0_io_out_b_0;
	wire _mesh_2_0_io_out_control_0_dataflow;
	wire _mesh_2_0_io_out_control_0_propagate;
	wire [4:0] _mesh_2_0_io_out_control_0_shift;
	wire [2:0] _mesh_2_0_io_out_id_0;
	wire _mesh_2_0_io_out_last_0;
	wire _mesh_2_0_io_out_valid_0;
	wire [31:0] _mesh_1_3_io_out_a_0;
	wire [31:0] _mesh_1_3_io_out_c_0;
	wire [31:0] _mesh_1_3_io_out_b_0;
	wire _mesh_1_3_io_out_control_0_dataflow;
	wire _mesh_1_3_io_out_control_0_propagate;
	wire [4:0] _mesh_1_3_io_out_control_0_shift;
	wire [2:0] _mesh_1_3_io_out_id_0;
	wire _mesh_1_3_io_out_last_0;
	wire _mesh_1_3_io_out_valid_0;
	wire [31:0] _mesh_1_2_io_out_a_0;
	wire [31:0] _mesh_1_2_io_out_c_0;
	wire [31:0] _mesh_1_2_io_out_b_0;
	wire _mesh_1_2_io_out_control_0_dataflow;
	wire _mesh_1_2_io_out_control_0_propagate;
	wire [4:0] _mesh_1_2_io_out_control_0_shift;
	wire [2:0] _mesh_1_2_io_out_id_0;
	wire _mesh_1_2_io_out_last_0;
	wire _mesh_1_2_io_out_valid_0;
	wire [31:0] _mesh_1_1_io_out_a_0;
	wire [31:0] _mesh_1_1_io_out_c_0;
	wire [31:0] _mesh_1_1_io_out_b_0;
	wire _mesh_1_1_io_out_control_0_dataflow;
	wire _mesh_1_1_io_out_control_0_propagate;
	wire [4:0] _mesh_1_1_io_out_control_0_shift;
	wire [2:0] _mesh_1_1_io_out_id_0;
	wire _mesh_1_1_io_out_last_0;
	wire _mesh_1_1_io_out_valid_0;
	wire [31:0] _mesh_1_0_io_out_a_0;
	wire [31:0] _mesh_1_0_io_out_c_0;
	wire [31:0] _mesh_1_0_io_out_b_0;
	wire _mesh_1_0_io_out_control_0_dataflow;
	wire _mesh_1_0_io_out_control_0_propagate;
	wire [4:0] _mesh_1_0_io_out_control_0_shift;
	wire [2:0] _mesh_1_0_io_out_id_0;
	wire _mesh_1_0_io_out_last_0;
	wire _mesh_1_0_io_out_valid_0;
	wire [31:0] _mesh_0_3_io_out_a_0;
	wire [31:0] _mesh_0_3_io_out_c_0;
	wire [31:0] _mesh_0_3_io_out_b_0;
	wire _mesh_0_3_io_out_control_0_dataflow;
	wire _mesh_0_3_io_out_control_0_propagate;
	wire [4:0] _mesh_0_3_io_out_control_0_shift;
	wire [2:0] _mesh_0_3_io_out_id_0;
	wire _mesh_0_3_io_out_last_0;
	wire _mesh_0_3_io_out_valid_0;
	wire [31:0] _mesh_0_2_io_out_a_0;
	wire [31:0] _mesh_0_2_io_out_c_0;
	wire [31:0] _mesh_0_2_io_out_b_0;
	wire _mesh_0_2_io_out_control_0_dataflow;
	wire _mesh_0_2_io_out_control_0_propagate;
	wire [4:0] _mesh_0_2_io_out_control_0_shift;
	wire [2:0] _mesh_0_2_io_out_id_0;
	wire _mesh_0_2_io_out_last_0;
	wire _mesh_0_2_io_out_valid_0;
	wire [31:0] _mesh_0_1_io_out_a_0;
	wire [31:0] _mesh_0_1_io_out_c_0;
	wire [31:0] _mesh_0_1_io_out_b_0;
	wire _mesh_0_1_io_out_control_0_dataflow;
	wire _mesh_0_1_io_out_control_0_propagate;
	wire [4:0] _mesh_0_1_io_out_control_0_shift;
	wire [2:0] _mesh_0_1_io_out_id_0;
	wire _mesh_0_1_io_out_last_0;
	wire _mesh_0_1_io_out_valid_0;
	wire [31:0] _mesh_0_0_io_out_a_0;
	wire [31:0] _mesh_0_0_io_out_c_0;
	wire [31:0] _mesh_0_0_io_out_b_0;
	wire _mesh_0_0_io_out_control_0_dataflow;
	wire _mesh_0_0_io_out_control_0_propagate;
	wire [4:0] _mesh_0_0_io_out_control_0_shift;
	wire [2:0] _mesh_0_0_io_out_id_0;
	wire _mesh_0_0_io_out_last_0;
	wire _mesh_0_0_io_out_valid_0;
	reg [31:0] r_0;
	reg [31:0] r_1_0;
	reg [31:0] r_2_0;
	reg [31:0] r_3_0;
	reg [31:0] r_4_0;
	reg [31:0] r_5_0;
	reg [31:0] r_6_0;
	reg [31:0] r_7_0;
	reg [31:0] r_8_0;
	reg [31:0] r_9_0;
	reg [31:0] r_10_0;
	reg [31:0] r_11_0;
	reg [31:0] r_12_0;
	reg [31:0] r_13_0;
	reg [31:0] r_14_0;
	reg [31:0] r_15_0;
	reg [31:0] b_0;
	reg [31:0] b_1_0;
	reg [31:0] b_2_0;
	reg [31:0] b_3_0;
	reg [31:0] b_4_0;
	reg [31:0] b_5_0;
	reg [31:0] b_6_0;
	reg [31:0] b_7_0;
	reg [31:0] b_8_0;
	reg [31:0] b_9_0;
	reg [31:0] b_10_0;
	reg [31:0] b_11_0;
	reg [31:0] b_12_0;
	reg [31:0] b_13_0;
	reg [31:0] b_14_0;
	reg [31:0] b_15_0;
	reg [31:0] b_16_0;
	reg [31:0] b_17_0;
	reg [31:0] b_18_0;
	reg [31:0] b_19_0;
	reg [31:0] b_20_0;
	reg [31:0] b_21_0;
	reg [31:0] b_22_0;
	reg [31:0] b_23_0;
	reg [31:0] b_24_0;
	reg [31:0] b_25_0;
	reg [31:0] b_26_0;
	reg [31:0] b_27_0;
	reg [31:0] b_28_0;
	reg [31:0] b_29_0;
	reg [31:0] b_30_0;
	reg [31:0] b_31_0;
	reg [4:0] mesh_0_0_io_in_control_0_shift_b;
	reg mesh_0_0_io_in_control_0_dataflow_b;
	reg mesh_0_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_0_io_in_control_0_shift_b;
	reg mesh_1_0_io_in_control_0_dataflow_b;
	reg mesh_1_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_0_io_in_control_0_shift_b;
	reg mesh_2_0_io_in_control_0_dataflow_b;
	reg mesh_2_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_0_io_in_control_0_shift_b;
	reg mesh_3_0_io_in_control_0_dataflow_b;
	reg mesh_3_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_1_io_in_control_0_shift_b;
	reg mesh_0_1_io_in_control_0_dataflow_b;
	reg mesh_0_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_1_io_in_control_0_shift_b;
	reg mesh_1_1_io_in_control_0_dataflow_b;
	reg mesh_1_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_1_io_in_control_0_shift_b;
	reg mesh_2_1_io_in_control_0_dataflow_b;
	reg mesh_2_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_1_io_in_control_0_shift_b;
	reg mesh_3_1_io_in_control_0_dataflow_b;
	reg mesh_3_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_2_io_in_control_0_shift_b;
	reg mesh_0_2_io_in_control_0_dataflow_b;
	reg mesh_0_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_2_io_in_control_0_shift_b;
	reg mesh_1_2_io_in_control_0_dataflow_b;
	reg mesh_1_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_2_io_in_control_0_shift_b;
	reg mesh_2_2_io_in_control_0_dataflow_b;
	reg mesh_2_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_2_io_in_control_0_shift_b;
	reg mesh_3_2_io_in_control_0_dataflow_b;
	reg mesh_3_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_3_io_in_control_0_shift_b;
	reg mesh_0_3_io_in_control_0_dataflow_b;
	reg mesh_0_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_3_io_in_control_0_shift_b;
	reg mesh_1_3_io_in_control_0_dataflow_b;
	reg mesh_1_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_3_io_in_control_0_shift_b;
	reg mesh_2_3_io_in_control_0_dataflow_b;
	reg mesh_2_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_3_io_in_control_0_shift_b;
	reg mesh_3_3_io_in_control_0_dataflow_b;
	reg mesh_3_3_io_in_control_0_propagate_b;
	reg r_16_0;
	reg r_17_0;
	reg r_18_0;
	reg r_19_0;
	reg r_20_0;
	reg r_21_0;
	reg r_22_0;
	reg r_23_0;
	reg r_24_0;
	reg r_25_0;
	reg r_26_0;
	reg r_27_0;
	reg r_28_0;
	reg r_29_0;
	reg r_30_0;
	reg r_31_0;
	reg [2:0] r_32_0;
	reg [2:0] r_33_0;
	reg [2:0] r_34_0;
	reg [2:0] r_35_0;
	reg [2:0] r_36_0;
	reg [2:0] r_37_0;
	reg [2:0] r_38_0;
	reg [2:0] r_39_0;
	reg [2:0] r_40_0;
	reg [2:0] r_41_0;
	reg [2:0] r_42_0;
	reg [2:0] r_43_0;
	reg [2:0] r_44_0;
	reg [2:0] r_45_0;
	reg [2:0] r_46_0;
	reg [2:0] r_47_0;
	reg r_48_0;
	reg r_49_0;
	reg r_50_0;
	reg r_51_0;
	reg r_52_0;
	reg r_53_0;
	reg r_54_0;
	reg r_55_0;
	reg r_56_0;
	reg r_57_0;
	reg r_58_0;
	reg r_59_0;
	reg r_60_0;
	reg r_61_0;
	reg r_62_0;
	reg r_63_0;
	reg [31:0] r_64_0;
	reg [31:0] r_65_0;
	reg r_66_0;
	reg r_67_0_dataflow;
	reg [2:0] r_68_0;
	reg r_69_0;
	reg [31:0] r_70_0;
	reg [31:0] r_71_0;
	reg [31:0] r_76_0;
	reg [31:0] r_77_0;
	reg [31:0] r_82_0;
	reg [31:0] r_83_0;
	always @(posedge clock) begin
		r_0 <=( io_in_a_0_0) ^ ((fiEnable && (17 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1_0 <=( _mesh_0_0_io_out_a_0) ^ ((fiEnable && (18 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_2_0 <=( _mesh_0_1_io_out_a_0) ^ ((fiEnable && (19 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_3_0 <=( _mesh_0_2_io_out_a_0) ^ ((fiEnable && (20 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4_0 <=( io_in_a_1_0) ^ ((fiEnable && (21 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_5_0 <=( _mesh_1_0_io_out_a_0) ^ ((fiEnable && (22 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_6_0 <=( _mesh_1_1_io_out_a_0) ^ ((fiEnable && (23 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_7_0 <=( _mesh_1_2_io_out_a_0) ^ ((fiEnable && (24 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_8_0 <=( io_in_a_2_0) ^ ((fiEnable && (25 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_9_0 <=( _mesh_2_0_io_out_a_0) ^ ((fiEnable && (26 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_10_0 <=( _mesh_2_1_io_out_a_0) ^ ((fiEnable && (27 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_11_0 <=( _mesh_2_2_io_out_a_0) ^ ((fiEnable && (28 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_12_0 <=( io_in_a_3_0) ^ ((fiEnable && (29 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_13_0 <=( _mesh_3_0_io_out_a_0) ^ ((fiEnable && (30 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_14_0 <=( _mesh_3_1_io_out_a_0) ^ ((fiEnable && (31 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_15_0 <=( _mesh_3_2_io_out_a_0) ^ ((fiEnable && (32 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		if (io_in_valid_0_0) begin
			b_0 <=( io_in_b_0_0) ^ ((fiEnable && (33 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_16_0 <=( io_in_d_0_0) ^ ((fiEnable && (34 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_0_io_in_control_0_shift_b <=( io_in_control_0_0_shift) ^ ((fiEnable && (35 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_0_io_in_control_0_dataflow_b <=( io_in_control_0_0_dataflow) ^ ((fiEnable && (36 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_0_io_in_control_0_propagate_b <=( io_in_control_0_0_propagate) ^ ((fiEnable && (37 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_0_io_out_valid_0) begin
			b_1_0 <=( _mesh_0_0_io_out_b_0) ^ ((fiEnable && (38 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_17_0 <=( _mesh_0_0_io_out_c_0) ^ ((fiEnable && (39 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_0_io_in_control_0_shift_b <=( _mesh_0_0_io_out_control_0_shift) ^ ((fiEnable && (40 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_0_io_in_control_0_dataflow_b <=( _mesh_0_0_io_out_control_0_dataflow) ^ ((fiEnable && (41 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_0_io_in_control_0_propagate_b <=( _mesh_0_0_io_out_control_0_propagate) ^ ((fiEnable && (42 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_0_io_out_valid_0) begin
			b_2_0 <=( _mesh_1_0_io_out_b_0) ^ ((fiEnable && (43 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_18_0 <=( _mesh_1_0_io_out_c_0) ^ ((fiEnable && (44 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_0_io_in_control_0_shift_b <=( _mesh_1_0_io_out_control_0_shift) ^ ((fiEnable && (45 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_0_io_in_control_0_dataflow_b <=( _mesh_1_0_io_out_control_0_dataflow) ^ ((fiEnable && (46 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_0_io_in_control_0_propagate_b <=( _mesh_1_0_io_out_control_0_propagate) ^ ((fiEnable && (47 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_0_io_out_valid_0) begin
			b_3_0 <=( _mesh_2_0_io_out_b_0) ^ ((fiEnable && (48 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_19_0 <=( _mesh_2_0_io_out_c_0) ^ ((fiEnable && (49 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_0_io_in_control_0_shift_b <=( _mesh_2_0_io_out_control_0_shift) ^ ((fiEnable && (50 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_0_io_in_control_0_dataflow_b <=( _mesh_2_0_io_out_control_0_dataflow) ^ ((fiEnable && (51 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_0_io_in_control_0_propagate_b <=( _mesh_2_0_io_out_control_0_propagate) ^ ((fiEnable && (52 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_1_0) begin
			b_4_0 <=( io_in_b_1_0) ^ ((fiEnable && (53 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_20_0 <=( io_in_d_1_0) ^ ((fiEnable && (54 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_1_io_in_control_0_shift_b <=( io_in_control_1_0_shift) ^ ((fiEnable && (55 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_1_io_in_control_0_dataflow_b <=( io_in_control_1_0_dataflow) ^ ((fiEnable && (56 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_1_io_in_control_0_propagate_b <=( io_in_control_1_0_propagate) ^ ((fiEnable && (57 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_1_io_out_valid_0) begin
			b_5_0 <=( _mesh_0_1_io_out_b_0) ^ ((fiEnable && (58 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_21_0 <=( _mesh_0_1_io_out_c_0) ^ ((fiEnable && (59 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_1_io_in_control_0_shift_b <=( _mesh_0_1_io_out_control_0_shift) ^ ((fiEnable && (60 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_1_io_in_control_0_dataflow_b <=( _mesh_0_1_io_out_control_0_dataflow) ^ ((fiEnable && (61 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_1_io_in_control_0_propagate_b <=( _mesh_0_1_io_out_control_0_propagate) ^ ((fiEnable && (62 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_1_io_out_valid_0) begin
			b_6_0 <=( _mesh_1_1_io_out_b_0) ^ ((fiEnable && (63 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_22_0 <=( _mesh_1_1_io_out_c_0) ^ ((fiEnable && (64 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_1_io_in_control_0_shift_b <=( _mesh_1_1_io_out_control_0_shift) ^ ((fiEnable && (65 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_1_io_in_control_0_dataflow_b <=( _mesh_1_1_io_out_control_0_dataflow) ^ ((fiEnable && (66 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_1_io_in_control_0_propagate_b <=( _mesh_1_1_io_out_control_0_propagate) ^ ((fiEnable && (67 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_1_io_out_valid_0) begin
			b_7_0 <=( _mesh_2_1_io_out_b_0) ^ ((fiEnable && (68 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_23_0 <=( _mesh_2_1_io_out_c_0) ^ ((fiEnable && (69 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_1_io_in_control_0_shift_b <=( _mesh_2_1_io_out_control_0_shift) ^ ((fiEnable && (70 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_1_io_in_control_0_dataflow_b <=( _mesh_2_1_io_out_control_0_dataflow) ^ ((fiEnable && (71 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_1_io_in_control_0_propagate_b <=( _mesh_2_1_io_out_control_0_propagate) ^ ((fiEnable && (72 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_2_0) begin
			b_8_0 <=( io_in_b_2_0) ^ ((fiEnable && (73 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_24_0 <=( io_in_d_2_0) ^ ((fiEnable && (74 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_2_io_in_control_0_shift_b <=( io_in_control_2_0_shift) ^ ((fiEnable && (75 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_2_io_in_control_0_dataflow_b <=( io_in_control_2_0_dataflow) ^ ((fiEnable && (76 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_2_io_in_control_0_propagate_b <=( io_in_control_2_0_propagate) ^ ((fiEnable && (77 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_2_io_out_valid_0) begin
			b_9_0 <=( _mesh_0_2_io_out_b_0) ^ ((fiEnable && (78 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_25_0 <=( _mesh_0_2_io_out_c_0) ^ ((fiEnable && (79 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_2_io_in_control_0_shift_b <=( _mesh_0_2_io_out_control_0_shift) ^ ((fiEnable && (80 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_2_io_in_control_0_dataflow_b <=( _mesh_0_2_io_out_control_0_dataflow) ^ ((fiEnable && (81 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_2_io_in_control_0_propagate_b <=( _mesh_0_2_io_out_control_0_propagate) ^ ((fiEnable && (82 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_2_io_out_valid_0) begin
			b_10_0 <=( _mesh_1_2_io_out_b_0) ^ ((fiEnable && (83 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_26_0 <=( _mesh_1_2_io_out_c_0) ^ ((fiEnable && (84 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_2_io_in_control_0_shift_b <=( _mesh_1_2_io_out_control_0_shift) ^ ((fiEnable && (85 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_2_io_in_control_0_dataflow_b <=( _mesh_1_2_io_out_control_0_dataflow) ^ ((fiEnable && (86 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_2_io_in_control_0_propagate_b <=( _mesh_1_2_io_out_control_0_propagate) ^ ((fiEnable && (87 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_2_io_out_valid_0) begin
			b_11_0 <=( _mesh_2_2_io_out_b_0) ^ ((fiEnable && (88 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_27_0 <=( _mesh_2_2_io_out_c_0) ^ ((fiEnable && (89 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_2_io_in_control_0_shift_b <=( _mesh_2_2_io_out_control_0_shift) ^ ((fiEnable && (90 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_2_io_in_control_0_dataflow_b <=( _mesh_2_2_io_out_control_0_dataflow) ^ ((fiEnable && (91 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_2_io_in_control_0_propagate_b <=( _mesh_2_2_io_out_control_0_propagate) ^ ((fiEnable && (92 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_3_0) begin
			b_12_0 <=( io_in_b_3_0) ^ ((fiEnable && (93 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_28_0 <=( io_in_d_3_0) ^ ((fiEnable && (94 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_3_io_in_control_0_shift_b <=( io_in_control_3_0_shift) ^ ((fiEnable && (95 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_3_io_in_control_0_dataflow_b <=( io_in_control_3_0_dataflow) ^ ((fiEnable && (96 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_3_io_in_control_0_propagate_b <=( io_in_control_3_0_propagate) ^ ((fiEnable && (97 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_3_io_out_valid_0) begin
			b_13_0 <=( _mesh_0_3_io_out_b_0) ^ ((fiEnable && (98 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_29_0 <=( _mesh_0_3_io_out_c_0) ^ ((fiEnable && (99 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_3_io_in_control_0_shift_b <=( _mesh_0_3_io_out_control_0_shift) ^ ((fiEnable && (100 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_3_io_in_control_0_dataflow_b <=( _mesh_0_3_io_out_control_0_dataflow) ^ ((fiEnable && (101 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_3_io_in_control_0_propagate_b <=( _mesh_0_3_io_out_control_0_propagate) ^ ((fiEnable && (102 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_3_io_out_valid_0) begin
			b_14_0 <=( _mesh_1_3_io_out_b_0) ^ ((fiEnable && (103 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_30_0 <=( _mesh_1_3_io_out_c_0) ^ ((fiEnable && (104 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_3_io_in_control_0_shift_b <=( _mesh_1_3_io_out_control_0_shift) ^ ((fiEnable && (105 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_3_io_in_control_0_dataflow_b <=( _mesh_1_3_io_out_control_0_dataflow) ^ ((fiEnable && (106 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_3_io_in_control_0_propagate_b <=( _mesh_1_3_io_out_control_0_propagate) ^ ((fiEnable && (107 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_3_io_out_valid_0) begin
			b_15_0 <=( _mesh_2_3_io_out_b_0) ^ ((fiEnable && (108 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_31_0 <=( _mesh_2_3_io_out_c_0) ^ ((fiEnable && (109 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_3_io_in_control_0_shift_b <=( _mesh_2_3_io_out_control_0_shift) ^ ((fiEnable && (110 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_3_io_in_control_0_dataflow_b <=( _mesh_2_3_io_out_control_0_dataflow) ^ ((fiEnable && (111 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_3_io_in_control_0_propagate_b <=( _mesh_2_3_io_out_control_0_propagate) ^ ((fiEnable && (112 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		r_16_0 <=( io_in_valid_0_0) ^ ((fiEnable && (113 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_17_0 <=( _mesh_0_0_io_out_valid_0) ^ ((fiEnable && (114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_18_0 <=( _mesh_1_0_io_out_valid_0) ^ ((fiEnable && (115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_19_0 <=( _mesh_2_0_io_out_valid_0) ^ ((fiEnable && (116 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_20_0 <=( io_in_valid_1_0) ^ ((fiEnable && (117 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_21_0 <=( _mesh_0_1_io_out_valid_0) ^ ((fiEnable && (118 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_22_0 <=( _mesh_1_1_io_out_valid_0) ^ ((fiEnable && (119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_23_0 <=( _mesh_2_1_io_out_valid_0) ^ ((fiEnable && (120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_24_0 <=( io_in_valid_2_0) ^ ((fiEnable && (121 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_25_0 <=( _mesh_0_2_io_out_valid_0) ^ ((fiEnable && (122 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_26_0 <=( _mesh_1_2_io_out_valid_0) ^ ((fiEnable && (123 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_27_0 <=( _mesh_2_2_io_out_valid_0) ^ ((fiEnable && (124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_28_0 <=( io_in_valid_3_0) ^ ((fiEnable && (125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_29_0 <=( _mesh_0_3_io_out_valid_0) ^ ((fiEnable && (126 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_30_0 <=( _mesh_1_3_io_out_valid_0) ^ ((fiEnable && (127 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_31_0 <=( _mesh_2_3_io_out_valid_0) ^ ((fiEnable && (128 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_32_0 <=( io_in_id_0_0) ^ ((fiEnable && (129 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_33_0 <=( _mesh_0_0_io_out_id_0) ^ ((fiEnable && (130 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_34_0 <=( _mesh_1_0_io_out_id_0) ^ ((fiEnable && (131 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_35_0 <=( _mesh_2_0_io_out_id_0) ^ ((fiEnable && (132 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_36_0 <=( io_in_id_1_0) ^ ((fiEnable && (133 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_37_0 <=( _mesh_0_1_io_out_id_0) ^ ((fiEnable && (134 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_38_0 <=( _mesh_1_1_io_out_id_0) ^ ((fiEnable && (135 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_39_0 <=( _mesh_2_1_io_out_id_0) ^ ((fiEnable && (136 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_40_0 <=( io_in_id_2_0) ^ ((fiEnable && (137 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_41_0 <=( _mesh_0_2_io_out_id_0) ^ ((fiEnable && (138 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_42_0 <=( _mesh_1_2_io_out_id_0) ^ ((fiEnable && (139 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_43_0 <=( _mesh_2_2_io_out_id_0) ^ ((fiEnable && (140 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_44_0 <=( io_in_id_3_0) ^ ((fiEnable && (141 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_45_0 <=( _mesh_0_3_io_out_id_0) ^ ((fiEnable && (142 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_46_0 <=( _mesh_1_3_io_out_id_0) ^ ((fiEnable && (143 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_47_0 <=( _mesh_2_3_io_out_id_0) ^ ((fiEnable && (144 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_48_0 <=( io_in_last_0_0) ^ ((fiEnable && (145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_49_0 <=( _mesh_0_0_io_out_last_0) ^ ((fiEnable && (146 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_50_0 <=( _mesh_1_0_io_out_last_0) ^ ((fiEnable && (147 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_51_0 <=( _mesh_2_0_io_out_last_0) ^ ((fiEnable && (148 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_52_0 <=( io_in_last_1_0) ^ ((fiEnable && (149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_53_0 <=( _mesh_0_1_io_out_last_0) ^ ((fiEnable && (150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_54_0 <=( _mesh_1_1_io_out_last_0) ^ ((fiEnable && (151 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_55_0 <=( _mesh_2_1_io_out_last_0) ^ ((fiEnable && (152 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_56_0 <=( io_in_last_2_0) ^ ((fiEnable && (153 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_57_0 <=( _mesh_0_2_io_out_last_0) ^ ((fiEnable && (154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_58_0 <=( _mesh_1_2_io_out_last_0) ^ ((fiEnable && (155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_59_0 <=( _mesh_2_2_io_out_last_0) ^ ((fiEnable && (156 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_60_0 <=( io_in_last_3_0) ^ ((fiEnable && (157 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_61_0 <=( _mesh_0_3_io_out_last_0) ^ ((fiEnable && (158 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_62_0 <=( _mesh_1_3_io_out_last_0) ^ ((fiEnable && (159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_63_0 <=( _mesh_2_3_io_out_last_0) ^ ((fiEnable && (160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_64_0 <=( _mesh_3_0_io_out_b_0) ^ ((fiEnable && (161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_65_0 <=( _mesh_3_0_io_out_c_0) ^ ((fiEnable && (162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_66_0 <=( _mesh_3_0_io_out_valid_0) ^ ((fiEnable && (163 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_67_0_dataflow <=( _mesh_3_0_io_out_control_0_dataflow) ^ ((fiEnable && (164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_68_0 <=( _mesh_3_0_io_out_id_0) ^ ((fiEnable && (165 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_69_0 <=( _mesh_3_0_io_out_last_0) ^ ((fiEnable && (166 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_70_0 <=( _mesh_3_1_io_out_b_0) ^ ((fiEnable && (167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_71_0 <=( _mesh_3_1_io_out_c_0) ^ ((fiEnable && (168 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_76_0 <=( _mesh_3_2_io_out_b_0) ^ ((fiEnable && (169 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_77_0 <=( _mesh_3_2_io_out_c_0) ^ ((fiEnable && (170 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_82_0 <=( _mesh_3_3_io_out_b_0) ^ ((fiEnable && (171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_83_0 <=( _mesh_3_3_io_out_c_0) ^ ((fiEnable && (172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	logic [31:0] _RANDOM_3;
	logic [31:0] _RANDOM_4;
	logic [31:0] _RANDOM_5;
	logic [31:0] _RANDOM_6;
	logic [31:0] _RANDOM_7;
	logic [31:0] _RANDOM_8;
	logic [31:0] _RANDOM_9;
	logic [31:0] _RANDOM_10;
	logic [31:0] _RANDOM_11;
	logic [31:0] _RANDOM_12;
	logic [31:0] _RANDOM_13;
	logic [31:0] _RANDOM_14;
	logic [31:0] _RANDOM_15;
	logic [31:0] _RANDOM_16;
	logic [31:0] _RANDOM_17;
	logic [31:0] _RANDOM_18;
	logic [31:0] _RANDOM_19;
	logic [31:0] _RANDOM_20;
	logic [31:0] _RANDOM_21;
	logic [31:0] _RANDOM_22;
	logic [31:0] _RANDOM_23;
	logic [31:0] _RANDOM_24;
	logic [31:0] _RANDOM_25;
	logic [31:0] _RANDOM_26;
	logic [31:0] _RANDOM_27;
	logic [31:0] _RANDOM_28;
	logic [31:0] _RANDOM_29;
	logic [31:0] _RANDOM_30;
	logic [31:0] _RANDOM_31;
	logic [31:0] _RANDOM_32;
	logic [31:0] _RANDOM_33;
	logic [31:0] _RANDOM_34;
	logic [31:0] _RANDOM_35;
	logic [31:0] _RANDOM_36;
	logic [31:0] _RANDOM_37;
	logic [31:0] _RANDOM_38;
	logic [31:0] _RANDOM_39;
	logic [31:0] _RANDOM_40;
	logic [31:0] _RANDOM_41;
	logic [31:0] _RANDOM_42;
	logic [31:0] _RANDOM_43;
	logic [31:0] _RANDOM_44;
	logic [31:0] _RANDOM_45;
	logic [31:0] _RANDOM_46;
	logic [31:0] _RANDOM_47;
	logic [31:0] _RANDOM_48;
	logic [31:0] _RANDOM_49;
	logic [31:0] _RANDOM_50;
	logic [31:0] _RANDOM_51;
	logic [31:0] _RANDOM_52;
	logic [31:0] _RANDOM_53;
	logic [31:0] _RANDOM_54;
	logic [31:0] _RANDOM_55;
	logic [31:0] _RANDOM_56;
	logic [31:0] _RANDOM_57;
	logic [31:0] _RANDOM_58;
	logic [31:0] _RANDOM_59;
	logic [31:0] _RANDOM_60;
	logic [31:0] _RANDOM_61;
	logic [31:0] _RANDOM_62;
	logic [31:0] _RANDOM_63;
	logic [31:0] _RANDOM_64;
	logic [31:0] _RANDOM_65;
	Tile mesh_0_0(
		.clock(clock),
		.io_in_a_0(r_0),
		.io_in_b_0(b_0),
		.io_in_d_0(b_16_0),
		.io_in_control_0_dataflow(mesh_0_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_0_io_in_control_0_shift_b),
		.io_in_id_0(r_32_0),
		.io_in_last_0(r_48_0),
		.io_in_valid_0(r_16_0),
		.io_out_a_0(_mesh_0_0_io_out_a_0),
		.io_out_c_0(_mesh_0_0_io_out_c_0),
		.io_out_b_0(_mesh_0_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_0_io_out_id_0),
		.io_out_last_0(_mesh_0_0_io_out_last_0),
		.io_out_valid_0(_mesh_0_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((187 == GlobalFiModInstNr[0]) || (187 == GlobalFiModInstNr[1]) || (187 == GlobalFiModInstNr[2]) || (187 == GlobalFiModInstNr[3]))));
	Tile mesh_0_1(
		.clock(clock),
		.io_in_a_0(r_1_0),
		.io_in_b_0(b_4_0),
		.io_in_d_0(b_20_0),
		.io_in_control_0_dataflow(mesh_0_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_1_io_in_control_0_shift_b),
		.io_in_id_0(r_36_0),
		.io_in_last_0(r_52_0),
		.io_in_valid_0(r_20_0),
		.io_out_a_0(_mesh_0_1_io_out_a_0),
		.io_out_c_0(_mesh_0_1_io_out_c_0),
		.io_out_b_0(_mesh_0_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_1_io_out_id_0),
		.io_out_last_0(_mesh_0_1_io_out_last_0),
		.io_out_valid_0(_mesh_0_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((188 == GlobalFiModInstNr[0]) || (188 == GlobalFiModInstNr[1]) || (188 == GlobalFiModInstNr[2]) || (188 == GlobalFiModInstNr[3]))));
	Tile mesh_0_2(
		.clock(clock),
		.io_in_a_0(r_2_0),
		.io_in_b_0(b_8_0),
		.io_in_d_0(b_24_0),
		.io_in_control_0_dataflow(mesh_0_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_2_io_in_control_0_shift_b),
		.io_in_id_0(r_40_0),
		.io_in_last_0(r_56_0),
		.io_in_valid_0(r_24_0),
		.io_out_a_0(_mesh_0_2_io_out_a_0),
		.io_out_c_0(_mesh_0_2_io_out_c_0),
		.io_out_b_0(_mesh_0_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_2_io_out_id_0),
		.io_out_last_0(_mesh_0_2_io_out_last_0),
		.io_out_valid_0(_mesh_0_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((189 == GlobalFiModInstNr[0]) || (189 == GlobalFiModInstNr[1]) || (189 == GlobalFiModInstNr[2]) || (189 == GlobalFiModInstNr[3]))));
	Tile mesh_0_3(
		.clock(clock),
		.io_in_a_0(r_3_0),
		.io_in_b_0(b_12_0),
		.io_in_d_0(b_28_0),
		.io_in_control_0_dataflow(mesh_0_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_3_io_in_control_0_shift_b),
		.io_in_id_0(r_44_0),
		.io_in_last_0(r_60_0),
		.io_in_valid_0(r_28_0),
		.io_out_a_0(_mesh_0_3_io_out_a_0),
		.io_out_c_0(_mesh_0_3_io_out_c_0),
		.io_out_b_0(_mesh_0_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_3_io_out_id_0),
		.io_out_last_0(_mesh_0_3_io_out_last_0),
		.io_out_valid_0(_mesh_0_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((190 == GlobalFiModInstNr[0]) || (190 == GlobalFiModInstNr[1]) || (190 == GlobalFiModInstNr[2]) || (190 == GlobalFiModInstNr[3]))));
	Tile mesh_1_0(
		.clock(clock),
		.io_in_a_0(r_4_0),
		.io_in_b_0(b_1_0),
		.io_in_d_0(b_17_0),
		.io_in_control_0_dataflow(mesh_1_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_0_io_in_control_0_shift_b),
		.io_in_id_0(r_33_0),
		.io_in_last_0(r_49_0),
		.io_in_valid_0(r_17_0),
		.io_out_a_0(_mesh_1_0_io_out_a_0),
		.io_out_c_0(_mesh_1_0_io_out_c_0),
		.io_out_b_0(_mesh_1_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_0_io_out_id_0),
		.io_out_last_0(_mesh_1_0_io_out_last_0),
		.io_out_valid_0(_mesh_1_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((191 == GlobalFiModInstNr[0]) || (191 == GlobalFiModInstNr[1]) || (191 == GlobalFiModInstNr[2]) || (191 == GlobalFiModInstNr[3]))));
	Tile mesh_1_1(
		.clock(clock),
		.io_in_a_0(r_5_0),
		.io_in_b_0(b_5_0),
		.io_in_d_0(b_21_0),
		.io_in_control_0_dataflow(mesh_1_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_1_io_in_control_0_shift_b),
		.io_in_id_0(r_37_0),
		.io_in_last_0(r_53_0),
		.io_in_valid_0(r_21_0),
		.io_out_a_0(_mesh_1_1_io_out_a_0),
		.io_out_c_0(_mesh_1_1_io_out_c_0),
		.io_out_b_0(_mesh_1_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_1_io_out_id_0),
		.io_out_last_0(_mesh_1_1_io_out_last_0),
		.io_out_valid_0(_mesh_1_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((192 == GlobalFiModInstNr[0]) || (192 == GlobalFiModInstNr[1]) || (192 == GlobalFiModInstNr[2]) || (192 == GlobalFiModInstNr[3]))));
	Tile mesh_1_2(
		.clock(clock),
		.io_in_a_0(r_6_0),
		.io_in_b_0(b_9_0),
		.io_in_d_0(b_25_0),
		.io_in_control_0_dataflow(mesh_1_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_2_io_in_control_0_shift_b),
		.io_in_id_0(r_41_0),
		.io_in_last_0(r_57_0),
		.io_in_valid_0(r_25_0),
		.io_out_a_0(_mesh_1_2_io_out_a_0),
		.io_out_c_0(_mesh_1_2_io_out_c_0),
		.io_out_b_0(_mesh_1_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_2_io_out_id_0),
		.io_out_last_0(_mesh_1_2_io_out_last_0),
		.io_out_valid_0(_mesh_1_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((193 == GlobalFiModInstNr[0]) || (193 == GlobalFiModInstNr[1]) || (193 == GlobalFiModInstNr[2]) || (193 == GlobalFiModInstNr[3]))));
	Tile mesh_1_3(
		.clock(clock),
		.io_in_a_0(r_7_0),
		.io_in_b_0(b_13_0),
		.io_in_d_0(b_29_0),
		.io_in_control_0_dataflow(mesh_1_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_3_io_in_control_0_shift_b),
		.io_in_id_0(r_45_0),
		.io_in_last_0(r_61_0),
		.io_in_valid_0(r_29_0),
		.io_out_a_0(_mesh_1_3_io_out_a_0),
		.io_out_c_0(_mesh_1_3_io_out_c_0),
		.io_out_b_0(_mesh_1_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_3_io_out_id_0),
		.io_out_last_0(_mesh_1_3_io_out_last_0),
		.io_out_valid_0(_mesh_1_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((194 == GlobalFiModInstNr[0]) || (194 == GlobalFiModInstNr[1]) || (194 == GlobalFiModInstNr[2]) || (194 == GlobalFiModInstNr[3]))));
	Tile mesh_2_0(
		.clock(clock),
		.io_in_a_0(r_8_0),
		.io_in_b_0(b_2_0),
		.io_in_d_0(b_18_0),
		.io_in_control_0_dataflow(mesh_2_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_0_io_in_control_0_shift_b),
		.io_in_id_0(r_34_0),
		.io_in_last_0(r_50_0),
		.io_in_valid_0(r_18_0),
		.io_out_a_0(_mesh_2_0_io_out_a_0),
		.io_out_c_0(_mesh_2_0_io_out_c_0),
		.io_out_b_0(_mesh_2_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_0_io_out_id_0),
		.io_out_last_0(_mesh_2_0_io_out_last_0),
		.io_out_valid_0(_mesh_2_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((195 == GlobalFiModInstNr[0]) || (195 == GlobalFiModInstNr[1]) || (195 == GlobalFiModInstNr[2]) || (195 == GlobalFiModInstNr[3]))));
	Tile mesh_2_1(
		.clock(clock),
		.io_in_a_0(r_9_0),
		.io_in_b_0(b_6_0),
		.io_in_d_0(b_22_0),
		.io_in_control_0_dataflow(mesh_2_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_1_io_in_control_0_shift_b),
		.io_in_id_0(r_38_0),
		.io_in_last_0(r_54_0),
		.io_in_valid_0(r_22_0),
		.io_out_a_0(_mesh_2_1_io_out_a_0),
		.io_out_c_0(_mesh_2_1_io_out_c_0),
		.io_out_b_0(_mesh_2_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_1_io_out_id_0),
		.io_out_last_0(_mesh_2_1_io_out_last_0),
		.io_out_valid_0(_mesh_2_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((196 == GlobalFiModInstNr[0]) || (196 == GlobalFiModInstNr[1]) || (196 == GlobalFiModInstNr[2]) || (196 == GlobalFiModInstNr[3]))));
	Tile mesh_2_2(
		.clock(clock),
		.io_in_a_0(r_10_0),
		.io_in_b_0(b_10_0),
		.io_in_d_0(b_26_0),
		.io_in_control_0_dataflow(mesh_2_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_2_io_in_control_0_shift_b),
		.io_in_id_0(r_42_0),
		.io_in_last_0(r_58_0),
		.io_in_valid_0(r_26_0),
		.io_out_a_0(_mesh_2_2_io_out_a_0),
		.io_out_c_0(_mesh_2_2_io_out_c_0),
		.io_out_b_0(_mesh_2_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_2_io_out_id_0),
		.io_out_last_0(_mesh_2_2_io_out_last_0),
		.io_out_valid_0(_mesh_2_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((197 == GlobalFiModInstNr[0]) || (197 == GlobalFiModInstNr[1]) || (197 == GlobalFiModInstNr[2]) || (197 == GlobalFiModInstNr[3]))));
	Tile mesh_2_3(
		.clock(clock),
		.io_in_a_0(r_11_0),
		.io_in_b_0(b_14_0),
		.io_in_d_0(b_30_0),
		.io_in_control_0_dataflow(mesh_2_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_3_io_in_control_0_shift_b),
		.io_in_id_0(r_46_0),
		.io_in_last_0(r_62_0),
		.io_in_valid_0(r_30_0),
		.io_out_a_0(_mesh_2_3_io_out_a_0),
		.io_out_c_0(_mesh_2_3_io_out_c_0),
		.io_out_b_0(_mesh_2_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_3_io_out_id_0),
		.io_out_last_0(_mesh_2_3_io_out_last_0),
		.io_out_valid_0(_mesh_2_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((198 == GlobalFiModInstNr[0]) || (198 == GlobalFiModInstNr[1]) || (198 == GlobalFiModInstNr[2]) || (198 == GlobalFiModInstNr[3]))));
	Tile mesh_3_0(
		.clock(clock),
		.io_in_a_0(r_12_0),
		.io_in_b_0(b_3_0),
		.io_in_d_0(b_19_0),
		.io_in_control_0_dataflow(mesh_3_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_0_io_in_control_0_shift_b),
		.io_in_id_0(r_35_0),
		.io_in_last_0(r_51_0),
		.io_in_valid_0(r_19_0),
		.io_out_a_0(_mesh_3_0_io_out_a_0),
		.io_out_c_0(_mesh_3_0_io_out_c_0),
		.io_out_b_0(_mesh_3_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_0_io_out_id_0),
		.io_out_last_0(_mesh_3_0_io_out_last_0),
		.io_out_valid_0(_mesh_3_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((199 == GlobalFiModInstNr[0]) || (199 == GlobalFiModInstNr[1]) || (199 == GlobalFiModInstNr[2]) || (199 == GlobalFiModInstNr[3]))));
	Tile mesh_3_1(
		.clock(clock),
		.io_in_a_0(r_13_0),
		.io_in_b_0(b_7_0),
		.io_in_d_0(b_23_0),
		.io_in_control_0_dataflow(mesh_3_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_1_io_in_control_0_shift_b),
		.io_in_id_0(r_39_0),
		.io_in_last_0(r_55_0),
		.io_in_valid_0(r_23_0),
		.io_out_a_0(_mesh_3_1_io_out_a_0),
		.io_out_c_0(_mesh_3_1_io_out_c_0),
		.io_out_b_0(_mesh_3_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_1_io_out_id_0),
		.io_out_last_0(_mesh_3_1_io_out_last_0),
		.io_out_valid_0(_mesh_3_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((200 == GlobalFiModInstNr[0]) || (200 == GlobalFiModInstNr[1]) || (200 == GlobalFiModInstNr[2]) || (200 == GlobalFiModInstNr[3]))));
	Tile mesh_3_2(
		.clock(clock),
		.io_in_a_0(r_14_0),
		.io_in_b_0(b_11_0),
		.io_in_d_0(b_27_0),
		.io_in_control_0_dataflow(mesh_3_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_2_io_in_control_0_shift_b),
		.io_in_id_0(r_43_0),
		.io_in_last_0(r_59_0),
		.io_in_valid_0(r_27_0),
		.io_out_a_0(_mesh_3_2_io_out_a_0),
		.io_out_c_0(_mesh_3_2_io_out_c_0),
		.io_out_b_0(_mesh_3_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_2_io_out_id_0),
		.io_out_last_0(_mesh_3_2_io_out_last_0),
		.io_out_valid_0(_mesh_3_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((201 == GlobalFiModInstNr[0]) || (201 == GlobalFiModInstNr[1]) || (201 == GlobalFiModInstNr[2]) || (201 == GlobalFiModInstNr[3]))));
	Tile mesh_3_3(
		.clock(clock),
		.io_in_a_0(r_15_0),
		.io_in_b_0(b_15_0),
		.io_in_d_0(b_31_0),
		.io_in_control_0_dataflow(mesh_3_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_3_io_in_control_0_shift_b),
		.io_in_id_0(r_47_0),
		.io_in_last_0(r_63_0),
		.io_in_valid_0(r_31_0),
		.io_out_a_0(_mesh_3_3_io_out_a_0),
		.io_out_c_0(_mesh_3_3_io_out_c_0),
		.io_out_b_0(_mesh_3_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_3_io_out_id_0),
		.io_out_last_0(_mesh_3_3_io_out_last_0),
		.io_out_valid_0(_mesh_3_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((202 == GlobalFiModInstNr[0]) || (202 == GlobalFiModInstNr[1]) || (202 == GlobalFiModInstNr[2]) || (202 == GlobalFiModInstNr[3]))));
	assign io_out_b_0_0 =( r_64_0) ^ ((fiEnable && (173 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_1_0 =( r_70_0) ^ ((fiEnable && (174 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_2_0 =( r_76_0) ^ ((fiEnable && (175 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_3_0 =( r_82_0) ^ ((fiEnable && (176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_0_0 =( r_65_0) ^ ((fiEnable && (177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_1_0 =( r_71_0) ^ ((fiEnable && (178 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_2_0 =( r_77_0) ^ ((fiEnable && (179 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_3_0 =( r_83_0) ^ ((fiEnable && (180 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_valid_0_0 =( r_66_0) ^ ((fiEnable && (181 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_0_0_dataflow =( r_67_0_dataflow) ^ ((fiEnable && (182 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_id_0_0 =( r_68_0) ^ ((fiEnable && (183 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last_0_0 =( r_69_0) ^ ((fiEnable && (184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
endmodule