module MacUnit (
	io_in_a,
	io_in_b,
	io_in_c,
	io_out_d
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_c;
	output logic [31:0] io_out_d;
	assign io_out_d =( (io_in_a * io_in_b) + io_in_c) ^ ((fiEnable && (2 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
endmodule
module PE_1024 (
	clock,
	io_in_a,
	io_in_b,
	io_in_d,
	io_in_control_dataflow,
	io_in_control_propagate,
	io_in_control_shift,
	io_in_id,
	io_in_last,
	io_in_valid,
	io_out_a,
	io_out_b,
	io_out_c,
	io_out_control_dataflow,
	io_out_control_propagate,
	io_out_control_shift,
	io_out_id,
	io_out_last,
	io_out_valid
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_d;
	input io_in_control_dataflow;
	input io_in_control_propagate;
	input [4:0] io_in_control_shift;
	input [2:0] io_in_id;
	input io_in_last;
	input io_in_valid;
	output logic [31:0] io_out_a;
	output logic [31:0] io_out_b;
	output logic [31:0] io_out_c;
	output logic io_out_control_dataflow;
	output logic io_out_control_propagate;
	output logic [4:0] io_out_control_shift;
	output logic [2:0] io_out_id;
	output logic io_out_last;
	output logic io_out_valid;
	wire [31:0] _mac_unit_io_out_d;
	reg [31:0] c1;
	reg [31:0] c2;
	reg last_s;
	wire [4:0] shift_offset = (last_s != io_in_control_propagate ? io_in_control_shift : 5'h00);
	wire [31:0] _GEN = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_3 = $signed($signed(c1) >>> _GEN);
	wire [31:0] _GEN_0 = {27'h0000000, shift_offset};
	wire [31:0] _io_out_c_T = $signed($signed(c1) >>> _GEN_0);
	wire [31:0] _GEN_1 = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_8 = $signed($signed(c2) >>> _GEN_1);
	wire [31:0] _io_out_c_T_11 = $signed($signed(c2) >>> _GEN_0);
	always @(posedge clock)
		if (io_in_valid) begin
			if (io_in_control_propagate) begin
				c1 <=( io_in_d) ^ ((fiEnable && (3 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( _mac_unit_io_out_d) ^ ((fiEnable && (4 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			end
			else begin
				c1 <=( _mac_unit_io_out_d) ^ ((fiEnable && (5 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( io_in_d) ^ ((fiEnable && (6 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			end
			last_s <=( io_in_control_propagate) ^ ((fiEnable && (7 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
		end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	MacUnit mac_unit(
		.io_in_a(io_in_a),
		.io_in_b(io_in_b),
		.io_in_c((io_in_control_propagate ? c2 : c1)),
		.io_out_d(_mac_unit_io_out_d)
	,
    .fiEnable(fiEnable && ((9369 == Mesh.GlobalFiModInstNr[0]) || (9369 == Mesh.GlobalFiModInstNr[1]) || (9369 == Mesh.GlobalFiModInstNr[2]) || (9369 == Mesh.GlobalFiModInstNr[3]))));
	assign io_out_a =( io_in_a) ^ ((fiEnable && (8 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b =( io_in_b) ^ ((fiEnable && (9 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c =( (io_in_control_propagate ? _io_out_c_T + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_3[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c1 & ((32'h00000001 << _GEN) - 32'h00000001)) | _io_out_c_T[0])} : _io_out_c_T_11 + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_8[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c2 & ((32'h00000001 << _GEN_1) - 32'h00000001)) | _io_out_c_T_11[0])})) ^ ((fiEnable && (10 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_control_dataflow =( io_in_control_dataflow) ^ ((fiEnable && (11 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_propagate =( io_in_control_propagate) ^ ((fiEnable && (12 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_shift =( io_in_control_shift) ^ ((fiEnable && (13 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[4:0] : {5{1'b0}});
	assign io_out_id =( io_in_id) ^ ((fiEnable && (14 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last =( io_in_last) ^ ((fiEnable && (15 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_valid =( io_in_valid) ^ ((fiEnable && (16 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
endmodule
module Tile (
	clock,
	io_in_a_0,
	io_in_b_0,
	io_in_d_0,
	io_in_control_0_dataflow,
	io_in_control_0_propagate,
	io_in_control_0_shift,
	io_in_id_0,
	io_in_last_0,
	io_in_valid_0,
	io_out_a_0,
	io_out_c_0,
	io_out_b_0,
	io_out_control_0_dataflow,
	io_out_control_0_propagate,
	io_out_control_0_shift,
	io_out_id_0,
	io_out_last_0,
	io_out_valid_0
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a_0;
	input [31:0] io_in_b_0;
	input [31:0] io_in_d_0;
	input io_in_control_0_dataflow;
	input io_in_control_0_propagate;
	input [4:0] io_in_control_0_shift;
	input [2:0] io_in_id_0;
	input io_in_last_0;
	input io_in_valid_0;
	output logic [31:0] io_out_a_0;
	output logic [31:0] io_out_c_0;
	output logic [31:0] io_out_b_0;
	output logic io_out_control_0_dataflow;
	output logic io_out_control_0_propagate;
	output logic [4:0] io_out_control_0_shift;
	output logic [2:0] io_out_id_0;
	output logic io_out_last_0;
	output logic io_out_valid_0;
	PE_1024 tile_0_0(
		.clock(clock),
		.io_in_a(io_in_a_0),
		.io_in_b(io_in_b_0),
		.io_in_d(io_in_d_0),
		.io_in_control_dataflow(io_in_control_0_dataflow),
		.io_in_control_propagate(io_in_control_0_propagate),
		.io_in_control_shift(io_in_control_0_shift),
		.io_in_id(io_in_id_0),
		.io_in_last(io_in_last_0),
		.io_in_valid(io_in_valid_0),
		.io_out_a(io_out_a_0),
		.io_out_b(io_out_b_0),
		.io_out_c(io_out_c_0),
		.io_out_control_dataflow(io_out_control_0_dataflow),
		.io_out_control_propagate(io_out_control_0_propagate),
		.io_out_control_shift(io_out_control_0_shift),
		.io_out_id(io_out_id_0),
		.io_out_last(io_out_last_0),
		.io_out_valid(io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9370 == Mesh.GlobalFiModInstNr[0]) || (9370 == Mesh.GlobalFiModInstNr[1]) || (9370 == Mesh.GlobalFiModInstNr[2]) || (9370 == Mesh.GlobalFiModInstNr[3]))));
endmodule
module Mesh (
	clock,
	io_in_a_0_0,
	io_in_a_1_0,
	io_in_a_2_0,
	io_in_a_3_0,
	io_in_a_4_0,
	io_in_a_5_0,
	io_in_a_6_0,
	io_in_a_7_0,
	io_in_a_8_0,
	io_in_a_9_0,
	io_in_a_10_0,
	io_in_a_11_0,
	io_in_a_12_0,
	io_in_a_13_0,
	io_in_a_14_0,
	io_in_a_15_0,
	io_in_a_16_0,
	io_in_a_17_0,
	io_in_a_18_0,
	io_in_a_19_0,
	io_in_a_20_0,
	io_in_a_21_0,
	io_in_a_22_0,
	io_in_a_23_0,
	io_in_a_24_0,
	io_in_a_25_0,
	io_in_a_26_0,
	io_in_a_27_0,
	io_in_a_28_0,
	io_in_a_29_0,
	io_in_a_30_0,
	io_in_a_31_0,
	io_in_b_0_0,
	io_in_b_1_0,
	io_in_b_2_0,
	io_in_b_3_0,
	io_in_b_4_0,
	io_in_b_5_0,
	io_in_b_6_0,
	io_in_b_7_0,
	io_in_b_8_0,
	io_in_b_9_0,
	io_in_b_10_0,
	io_in_b_11_0,
	io_in_b_12_0,
	io_in_b_13_0,
	io_in_b_14_0,
	io_in_b_15_0,
	io_in_b_16_0,
	io_in_b_17_0,
	io_in_b_18_0,
	io_in_b_19_0,
	io_in_b_20_0,
	io_in_b_21_0,
	io_in_b_22_0,
	io_in_b_23_0,
	io_in_b_24_0,
	io_in_b_25_0,
	io_in_b_26_0,
	io_in_b_27_0,
	io_in_b_28_0,
	io_in_b_29_0,
	io_in_b_30_0,
	io_in_b_31_0,
	io_in_d_0_0,
	io_in_d_1_0,
	io_in_d_2_0,
	io_in_d_3_0,
	io_in_d_4_0,
	io_in_d_5_0,
	io_in_d_6_0,
	io_in_d_7_0,
	io_in_d_8_0,
	io_in_d_9_0,
	io_in_d_10_0,
	io_in_d_11_0,
	io_in_d_12_0,
	io_in_d_13_0,
	io_in_d_14_0,
	io_in_d_15_0,
	io_in_d_16_0,
	io_in_d_17_0,
	io_in_d_18_0,
	io_in_d_19_0,
	io_in_d_20_0,
	io_in_d_21_0,
	io_in_d_22_0,
	io_in_d_23_0,
	io_in_d_24_0,
	io_in_d_25_0,
	io_in_d_26_0,
	io_in_d_27_0,
	io_in_d_28_0,
	io_in_d_29_0,
	io_in_d_30_0,
	io_in_d_31_0,
	io_in_control_0_0_dataflow,
	io_in_control_0_0_propagate,
	io_in_control_0_0_shift,
	io_in_control_1_0_dataflow,
	io_in_control_1_0_propagate,
	io_in_control_1_0_shift,
	io_in_control_2_0_dataflow,
	io_in_control_2_0_propagate,
	io_in_control_2_0_shift,
	io_in_control_3_0_dataflow,
	io_in_control_3_0_propagate,
	io_in_control_3_0_shift,
	io_in_control_4_0_dataflow,
	io_in_control_4_0_propagate,
	io_in_control_4_0_shift,
	io_in_control_5_0_dataflow,
	io_in_control_5_0_propagate,
	io_in_control_5_0_shift,
	io_in_control_6_0_dataflow,
	io_in_control_6_0_propagate,
	io_in_control_6_0_shift,
	io_in_control_7_0_dataflow,
	io_in_control_7_0_propagate,
	io_in_control_7_0_shift,
	io_in_control_8_0_dataflow,
	io_in_control_8_0_propagate,
	io_in_control_8_0_shift,
	io_in_control_9_0_dataflow,
	io_in_control_9_0_propagate,
	io_in_control_9_0_shift,
	io_in_control_10_0_dataflow,
	io_in_control_10_0_propagate,
	io_in_control_10_0_shift,
	io_in_control_11_0_dataflow,
	io_in_control_11_0_propagate,
	io_in_control_11_0_shift,
	io_in_control_12_0_dataflow,
	io_in_control_12_0_propagate,
	io_in_control_12_0_shift,
	io_in_control_13_0_dataflow,
	io_in_control_13_0_propagate,
	io_in_control_13_0_shift,
	io_in_control_14_0_dataflow,
	io_in_control_14_0_propagate,
	io_in_control_14_0_shift,
	io_in_control_15_0_dataflow,
	io_in_control_15_0_propagate,
	io_in_control_15_0_shift,
	io_in_control_16_0_dataflow,
	io_in_control_16_0_propagate,
	io_in_control_16_0_shift,
	io_in_control_17_0_dataflow,
	io_in_control_17_0_propagate,
	io_in_control_17_0_shift,
	io_in_control_18_0_dataflow,
	io_in_control_18_0_propagate,
	io_in_control_18_0_shift,
	io_in_control_19_0_dataflow,
	io_in_control_19_0_propagate,
	io_in_control_19_0_shift,
	io_in_control_20_0_dataflow,
	io_in_control_20_0_propagate,
	io_in_control_20_0_shift,
	io_in_control_21_0_dataflow,
	io_in_control_21_0_propagate,
	io_in_control_21_0_shift,
	io_in_control_22_0_dataflow,
	io_in_control_22_0_propagate,
	io_in_control_22_0_shift,
	io_in_control_23_0_dataflow,
	io_in_control_23_0_propagate,
	io_in_control_23_0_shift,
	io_in_control_24_0_dataflow,
	io_in_control_24_0_propagate,
	io_in_control_24_0_shift,
	io_in_control_25_0_dataflow,
	io_in_control_25_0_propagate,
	io_in_control_25_0_shift,
	io_in_control_26_0_dataflow,
	io_in_control_26_0_propagate,
	io_in_control_26_0_shift,
	io_in_control_27_0_dataflow,
	io_in_control_27_0_propagate,
	io_in_control_27_0_shift,
	io_in_control_28_0_dataflow,
	io_in_control_28_0_propagate,
	io_in_control_28_0_shift,
	io_in_control_29_0_dataflow,
	io_in_control_29_0_propagate,
	io_in_control_29_0_shift,
	io_in_control_30_0_dataflow,
	io_in_control_30_0_propagate,
	io_in_control_30_0_shift,
	io_in_control_31_0_dataflow,
	io_in_control_31_0_propagate,
	io_in_control_31_0_shift,
	io_in_id_0_0,
	io_in_id_1_0,
	io_in_id_2_0,
	io_in_id_3_0,
	io_in_id_4_0,
	io_in_id_5_0,
	io_in_id_6_0,
	io_in_id_7_0,
	io_in_id_8_0,
	io_in_id_9_0,
	io_in_id_10_0,
	io_in_id_11_0,
	io_in_id_12_0,
	io_in_id_13_0,
	io_in_id_14_0,
	io_in_id_15_0,
	io_in_id_16_0,
	io_in_id_17_0,
	io_in_id_18_0,
	io_in_id_19_0,
	io_in_id_20_0,
	io_in_id_21_0,
	io_in_id_22_0,
	io_in_id_23_0,
	io_in_id_24_0,
	io_in_id_25_0,
	io_in_id_26_0,
	io_in_id_27_0,
	io_in_id_28_0,
	io_in_id_29_0,
	io_in_id_30_0,
	io_in_id_31_0,
	io_in_last_0_0,
	io_in_last_1_0,
	io_in_last_2_0,
	io_in_last_3_0,
	io_in_last_4_0,
	io_in_last_5_0,
	io_in_last_6_0,
	io_in_last_7_0,
	io_in_last_8_0,
	io_in_last_9_0,
	io_in_last_10_0,
	io_in_last_11_0,
	io_in_last_12_0,
	io_in_last_13_0,
	io_in_last_14_0,
	io_in_last_15_0,
	io_in_last_16_0,
	io_in_last_17_0,
	io_in_last_18_0,
	io_in_last_19_0,
	io_in_last_20_0,
	io_in_last_21_0,
	io_in_last_22_0,
	io_in_last_23_0,
	io_in_last_24_0,
	io_in_last_25_0,
	io_in_last_26_0,
	io_in_last_27_0,
	io_in_last_28_0,
	io_in_last_29_0,
	io_in_last_30_0,
	io_in_last_31_0,
	io_in_valid_0_0,
	io_in_valid_1_0,
	io_in_valid_2_0,
	io_in_valid_3_0,
	io_in_valid_4_0,
	io_in_valid_5_0,
	io_in_valid_6_0,
	io_in_valid_7_0,
	io_in_valid_8_0,
	io_in_valid_9_0,
	io_in_valid_10_0,
	io_in_valid_11_0,
	io_in_valid_12_0,
	io_in_valid_13_0,
	io_in_valid_14_0,
	io_in_valid_15_0,
	io_in_valid_16_0,
	io_in_valid_17_0,
	io_in_valid_18_0,
	io_in_valid_19_0,
	io_in_valid_20_0,
	io_in_valid_21_0,
	io_in_valid_22_0,
	io_in_valid_23_0,
	io_in_valid_24_0,
	io_in_valid_25_0,
	io_in_valid_26_0,
	io_in_valid_27_0,
	io_in_valid_28_0,
	io_in_valid_29_0,
	io_in_valid_30_0,
	io_in_valid_31_0,
	io_out_b_0_0,
	io_out_b_1_0,
	io_out_b_2_0,
	io_out_b_3_0,
	io_out_b_4_0,
	io_out_b_5_0,
	io_out_b_6_0,
	io_out_b_7_0,
	io_out_b_8_0,
	io_out_b_9_0,
	io_out_b_10_0,
	io_out_b_11_0,
	io_out_b_12_0,
	io_out_b_13_0,
	io_out_b_14_0,
	io_out_b_15_0,
	io_out_b_16_0,
	io_out_b_17_0,
	io_out_b_18_0,
	io_out_b_19_0,
	io_out_b_20_0,
	io_out_b_21_0,
	io_out_b_22_0,
	io_out_b_23_0,
	io_out_b_24_0,
	io_out_b_25_0,
	io_out_b_26_0,
	io_out_b_27_0,
	io_out_b_28_0,
	io_out_b_29_0,
	io_out_b_30_0,
	io_out_b_31_0,
	io_out_c_0_0,
	io_out_c_1_0,
	io_out_c_2_0,
	io_out_c_3_0,
	io_out_c_4_0,
	io_out_c_5_0,
	io_out_c_6_0,
	io_out_c_7_0,
	io_out_c_8_0,
	io_out_c_9_0,
	io_out_c_10_0,
	io_out_c_11_0,
	io_out_c_12_0,
	io_out_c_13_0,
	io_out_c_14_0,
	io_out_c_15_0,
	io_out_c_16_0,
	io_out_c_17_0,
	io_out_c_18_0,
	io_out_c_19_0,
	io_out_c_20_0,
	io_out_c_21_0,
	io_out_c_22_0,
	io_out_c_23_0,
	io_out_c_24_0,
	io_out_c_25_0,
	io_out_c_26_0,
	io_out_c_27_0,
	io_out_c_28_0,
	io_out_c_29_0,
	io_out_c_30_0,
	io_out_c_31_0,
	io_out_valid_0_0,
	io_out_control_0_0_dataflow,
	io_out_id_0_0,
	io_out_last_0_0
, GlobalFiSignal, GlobalFiNumber, GlobalFiModInstNr);
input GlobalFiSignal;
wire [31:0] GlobalFiSignal;
input GlobalFiNumber;
wire [31:0] GlobalFiNumber;
input GlobalFiModInstNr;
wire [15:0] GlobalFiModInstNr[4];
wire fiEnable;
assign fiEnable = (1 == GlobalFiModInstNr[0]) || (1 == GlobalFiModInstNr[1]) || (1 == GlobalFiModInstNr[2]) || (1 == GlobalFiModInstNr[3]);

	input clock;
	input [31:0] io_in_a_0_0;
	input [31:0] io_in_a_1_0;
	input [31:0] io_in_a_2_0;
	input [31:0] io_in_a_3_0;
	input [31:0] io_in_a_4_0;
	input [31:0] io_in_a_5_0;
	input [31:0] io_in_a_6_0;
	input [31:0] io_in_a_7_0;
	input [31:0] io_in_a_8_0;
	input [31:0] io_in_a_9_0;
	input [31:0] io_in_a_10_0;
	input [31:0] io_in_a_11_0;
	input [31:0] io_in_a_12_0;
	input [31:0] io_in_a_13_0;
	input [31:0] io_in_a_14_0;
	input [31:0] io_in_a_15_0;
	input [31:0] io_in_a_16_0;
	input [31:0] io_in_a_17_0;
	input [31:0] io_in_a_18_0;
	input [31:0] io_in_a_19_0;
	input [31:0] io_in_a_20_0;
	input [31:0] io_in_a_21_0;
	input [31:0] io_in_a_22_0;
	input [31:0] io_in_a_23_0;
	input [31:0] io_in_a_24_0;
	input [31:0] io_in_a_25_0;
	input [31:0] io_in_a_26_0;
	input [31:0] io_in_a_27_0;
	input [31:0] io_in_a_28_0;
	input [31:0] io_in_a_29_0;
	input [31:0] io_in_a_30_0;
	input [31:0] io_in_a_31_0;
	input [31:0] io_in_b_0_0;
	input [31:0] io_in_b_1_0;
	input [31:0] io_in_b_2_0;
	input [31:0] io_in_b_3_0;
	input [31:0] io_in_b_4_0;
	input [31:0] io_in_b_5_0;
	input [31:0] io_in_b_6_0;
	input [31:0] io_in_b_7_0;
	input [31:0] io_in_b_8_0;
	input [31:0] io_in_b_9_0;
	input [31:0] io_in_b_10_0;
	input [31:0] io_in_b_11_0;
	input [31:0] io_in_b_12_0;
	input [31:0] io_in_b_13_0;
	input [31:0] io_in_b_14_0;
	input [31:0] io_in_b_15_0;
	input [31:0] io_in_b_16_0;
	input [31:0] io_in_b_17_0;
	input [31:0] io_in_b_18_0;
	input [31:0] io_in_b_19_0;
	input [31:0] io_in_b_20_0;
	input [31:0] io_in_b_21_0;
	input [31:0] io_in_b_22_0;
	input [31:0] io_in_b_23_0;
	input [31:0] io_in_b_24_0;
	input [31:0] io_in_b_25_0;
	input [31:0] io_in_b_26_0;
	input [31:0] io_in_b_27_0;
	input [31:0] io_in_b_28_0;
	input [31:0] io_in_b_29_0;
	input [31:0] io_in_b_30_0;
	input [31:0] io_in_b_31_0;
	input [31:0] io_in_d_0_0;
	input [31:0] io_in_d_1_0;
	input [31:0] io_in_d_2_0;
	input [31:0] io_in_d_3_0;
	input [31:0] io_in_d_4_0;
	input [31:0] io_in_d_5_0;
	input [31:0] io_in_d_6_0;
	input [31:0] io_in_d_7_0;
	input [31:0] io_in_d_8_0;
	input [31:0] io_in_d_9_0;
	input [31:0] io_in_d_10_0;
	input [31:0] io_in_d_11_0;
	input [31:0] io_in_d_12_0;
	input [31:0] io_in_d_13_0;
	input [31:0] io_in_d_14_0;
	input [31:0] io_in_d_15_0;
	input [31:0] io_in_d_16_0;
	input [31:0] io_in_d_17_0;
	input [31:0] io_in_d_18_0;
	input [31:0] io_in_d_19_0;
	input [31:0] io_in_d_20_0;
	input [31:0] io_in_d_21_0;
	input [31:0] io_in_d_22_0;
	input [31:0] io_in_d_23_0;
	input [31:0] io_in_d_24_0;
	input [31:0] io_in_d_25_0;
	input [31:0] io_in_d_26_0;
	input [31:0] io_in_d_27_0;
	input [31:0] io_in_d_28_0;
	input [31:0] io_in_d_29_0;
	input [31:0] io_in_d_30_0;
	input [31:0] io_in_d_31_0;
	input io_in_control_0_0_dataflow;
	input io_in_control_0_0_propagate;
	input [4:0] io_in_control_0_0_shift;
	input io_in_control_1_0_dataflow;
	input io_in_control_1_0_propagate;
	input [4:0] io_in_control_1_0_shift;
	input io_in_control_2_0_dataflow;
	input io_in_control_2_0_propagate;
	input [4:0] io_in_control_2_0_shift;
	input io_in_control_3_0_dataflow;
	input io_in_control_3_0_propagate;
	input [4:0] io_in_control_3_0_shift;
	input io_in_control_4_0_dataflow;
	input io_in_control_4_0_propagate;
	input [4:0] io_in_control_4_0_shift;
	input io_in_control_5_0_dataflow;
	input io_in_control_5_0_propagate;
	input [4:0] io_in_control_5_0_shift;
	input io_in_control_6_0_dataflow;
	input io_in_control_6_0_propagate;
	input [4:0] io_in_control_6_0_shift;
	input io_in_control_7_0_dataflow;
	input io_in_control_7_0_propagate;
	input [4:0] io_in_control_7_0_shift;
	input io_in_control_8_0_dataflow;
	input io_in_control_8_0_propagate;
	input [4:0] io_in_control_8_0_shift;
	input io_in_control_9_0_dataflow;
	input io_in_control_9_0_propagate;
	input [4:0] io_in_control_9_0_shift;
	input io_in_control_10_0_dataflow;
	input io_in_control_10_0_propagate;
	input [4:0] io_in_control_10_0_shift;
	input io_in_control_11_0_dataflow;
	input io_in_control_11_0_propagate;
	input [4:0] io_in_control_11_0_shift;
	input io_in_control_12_0_dataflow;
	input io_in_control_12_0_propagate;
	input [4:0] io_in_control_12_0_shift;
	input io_in_control_13_0_dataflow;
	input io_in_control_13_0_propagate;
	input [4:0] io_in_control_13_0_shift;
	input io_in_control_14_0_dataflow;
	input io_in_control_14_0_propagate;
	input [4:0] io_in_control_14_0_shift;
	input io_in_control_15_0_dataflow;
	input io_in_control_15_0_propagate;
	input [4:0] io_in_control_15_0_shift;
	input io_in_control_16_0_dataflow;
	input io_in_control_16_0_propagate;
	input [4:0] io_in_control_16_0_shift;
	input io_in_control_17_0_dataflow;
	input io_in_control_17_0_propagate;
	input [4:0] io_in_control_17_0_shift;
	input io_in_control_18_0_dataflow;
	input io_in_control_18_0_propagate;
	input [4:0] io_in_control_18_0_shift;
	input io_in_control_19_0_dataflow;
	input io_in_control_19_0_propagate;
	input [4:0] io_in_control_19_0_shift;
	input io_in_control_20_0_dataflow;
	input io_in_control_20_0_propagate;
	input [4:0] io_in_control_20_0_shift;
	input io_in_control_21_0_dataflow;
	input io_in_control_21_0_propagate;
	input [4:0] io_in_control_21_0_shift;
	input io_in_control_22_0_dataflow;
	input io_in_control_22_0_propagate;
	input [4:0] io_in_control_22_0_shift;
	input io_in_control_23_0_dataflow;
	input io_in_control_23_0_propagate;
	input [4:0] io_in_control_23_0_shift;
	input io_in_control_24_0_dataflow;
	input io_in_control_24_0_propagate;
	input [4:0] io_in_control_24_0_shift;
	input io_in_control_25_0_dataflow;
	input io_in_control_25_0_propagate;
	input [4:0] io_in_control_25_0_shift;
	input io_in_control_26_0_dataflow;
	input io_in_control_26_0_propagate;
	input [4:0] io_in_control_26_0_shift;
	input io_in_control_27_0_dataflow;
	input io_in_control_27_0_propagate;
	input [4:0] io_in_control_27_0_shift;
	input io_in_control_28_0_dataflow;
	input io_in_control_28_0_propagate;
	input [4:0] io_in_control_28_0_shift;
	input io_in_control_29_0_dataflow;
	input io_in_control_29_0_propagate;
	input [4:0] io_in_control_29_0_shift;
	input io_in_control_30_0_dataflow;
	input io_in_control_30_0_propagate;
	input [4:0] io_in_control_30_0_shift;
	input io_in_control_31_0_dataflow;
	input io_in_control_31_0_propagate;
	input [4:0] io_in_control_31_0_shift;
	input [2:0] io_in_id_0_0;
	input [2:0] io_in_id_1_0;
	input [2:0] io_in_id_2_0;
	input [2:0] io_in_id_3_0;
	input [2:0] io_in_id_4_0;
	input [2:0] io_in_id_5_0;
	input [2:0] io_in_id_6_0;
	input [2:0] io_in_id_7_0;
	input [2:0] io_in_id_8_0;
	input [2:0] io_in_id_9_0;
	input [2:0] io_in_id_10_0;
	input [2:0] io_in_id_11_0;
	input [2:0] io_in_id_12_0;
	input [2:0] io_in_id_13_0;
	input [2:0] io_in_id_14_0;
	input [2:0] io_in_id_15_0;
	input [2:0] io_in_id_16_0;
	input [2:0] io_in_id_17_0;
	input [2:0] io_in_id_18_0;
	input [2:0] io_in_id_19_0;
	input [2:0] io_in_id_20_0;
	input [2:0] io_in_id_21_0;
	input [2:0] io_in_id_22_0;
	input [2:0] io_in_id_23_0;
	input [2:0] io_in_id_24_0;
	input [2:0] io_in_id_25_0;
	input [2:0] io_in_id_26_0;
	input [2:0] io_in_id_27_0;
	input [2:0] io_in_id_28_0;
	input [2:0] io_in_id_29_0;
	input [2:0] io_in_id_30_0;
	input [2:0] io_in_id_31_0;
	input io_in_last_0_0;
	input io_in_last_1_0;
	input io_in_last_2_0;
	input io_in_last_3_0;
	input io_in_last_4_0;
	input io_in_last_5_0;
	input io_in_last_6_0;
	input io_in_last_7_0;
	input io_in_last_8_0;
	input io_in_last_9_0;
	input io_in_last_10_0;
	input io_in_last_11_0;
	input io_in_last_12_0;
	input io_in_last_13_0;
	input io_in_last_14_0;
	input io_in_last_15_0;
	input io_in_last_16_0;
	input io_in_last_17_0;
	input io_in_last_18_0;
	input io_in_last_19_0;
	input io_in_last_20_0;
	input io_in_last_21_0;
	input io_in_last_22_0;
	input io_in_last_23_0;
	input io_in_last_24_0;
	input io_in_last_25_0;
	input io_in_last_26_0;
	input io_in_last_27_0;
	input io_in_last_28_0;
	input io_in_last_29_0;
	input io_in_last_30_0;
	input io_in_last_31_0;
	input io_in_valid_0_0;
	input io_in_valid_1_0;
	input io_in_valid_2_0;
	input io_in_valid_3_0;
	input io_in_valid_4_0;
	input io_in_valid_5_0;
	input io_in_valid_6_0;
	input io_in_valid_7_0;
	input io_in_valid_8_0;
	input io_in_valid_9_0;
	input io_in_valid_10_0;
	input io_in_valid_11_0;
	input io_in_valid_12_0;
	input io_in_valid_13_0;
	input io_in_valid_14_0;
	input io_in_valid_15_0;
	input io_in_valid_16_0;
	input io_in_valid_17_0;
	input io_in_valid_18_0;
	input io_in_valid_19_0;
	input io_in_valid_20_0;
	input io_in_valid_21_0;
	input io_in_valid_22_0;
	input io_in_valid_23_0;
	input io_in_valid_24_0;
	input io_in_valid_25_0;
	input io_in_valid_26_0;
	input io_in_valid_27_0;
	input io_in_valid_28_0;
	input io_in_valid_29_0;
	input io_in_valid_30_0;
	input io_in_valid_31_0;
	output logic [31:0] io_out_b_0_0;
	output logic [31:0] io_out_b_1_0;
	output logic [31:0] io_out_b_2_0;
	output logic [31:0] io_out_b_3_0;
	output logic [31:0] io_out_b_4_0;
	output logic [31:0] io_out_b_5_0;
	output logic [31:0] io_out_b_6_0;
	output logic [31:0] io_out_b_7_0;
	output logic [31:0] io_out_b_8_0;
	output logic [31:0] io_out_b_9_0;
	output logic [31:0] io_out_b_10_0;
	output logic [31:0] io_out_b_11_0;
	output logic [31:0] io_out_b_12_0;
	output logic [31:0] io_out_b_13_0;
	output logic [31:0] io_out_b_14_0;
	output logic [31:0] io_out_b_15_0;
	output logic [31:0] io_out_b_16_0;
	output logic [31:0] io_out_b_17_0;
	output logic [31:0] io_out_b_18_0;
	output logic [31:0] io_out_b_19_0;
	output logic [31:0] io_out_b_20_0;
	output logic [31:0] io_out_b_21_0;
	output logic [31:0] io_out_b_22_0;
	output logic [31:0] io_out_b_23_0;
	output logic [31:0] io_out_b_24_0;
	output logic [31:0] io_out_b_25_0;
	output logic [31:0] io_out_b_26_0;
	output logic [31:0] io_out_b_27_0;
	output logic [31:0] io_out_b_28_0;
	output logic [31:0] io_out_b_29_0;
	output logic [31:0] io_out_b_30_0;
	output logic [31:0] io_out_b_31_0;
	output logic [31:0] io_out_c_0_0;
	output logic [31:0] io_out_c_1_0;
	output logic [31:0] io_out_c_2_0;
	output logic [31:0] io_out_c_3_0;
	output logic [31:0] io_out_c_4_0;
	output logic [31:0] io_out_c_5_0;
	output logic [31:0] io_out_c_6_0;
	output logic [31:0] io_out_c_7_0;
	output logic [31:0] io_out_c_8_0;
	output logic [31:0] io_out_c_9_0;
	output logic [31:0] io_out_c_10_0;
	output logic [31:0] io_out_c_11_0;
	output logic [31:0] io_out_c_12_0;
	output logic [31:0] io_out_c_13_0;
	output logic [31:0] io_out_c_14_0;
	output logic [31:0] io_out_c_15_0;
	output logic [31:0] io_out_c_16_0;
	output logic [31:0] io_out_c_17_0;
	output logic [31:0] io_out_c_18_0;
	output logic [31:0] io_out_c_19_0;
	output logic [31:0] io_out_c_20_0;
	output logic [31:0] io_out_c_21_0;
	output logic [31:0] io_out_c_22_0;
	output logic [31:0] io_out_c_23_0;
	output logic [31:0] io_out_c_24_0;
	output logic [31:0] io_out_c_25_0;
	output logic [31:0] io_out_c_26_0;
	output logic [31:0] io_out_c_27_0;
	output logic [31:0] io_out_c_28_0;
	output logic [31:0] io_out_c_29_0;
	output logic [31:0] io_out_c_30_0;
	output logic [31:0] io_out_c_31_0;
	output logic io_out_valid_0_0;
	output logic io_out_control_0_0_dataflow;
	output logic [2:0] io_out_id_0_0;
	output logic io_out_last_0_0;
	wire [31:0] _mesh_31_31_io_out_a_0;
	wire [31:0] _mesh_31_31_io_out_c_0;
	wire [31:0] _mesh_31_31_io_out_b_0;
	wire _mesh_31_31_io_out_control_0_dataflow;
	wire _mesh_31_31_io_out_control_0_propagate;
	wire [4:0] _mesh_31_31_io_out_control_0_shift;
	wire [2:0] _mesh_31_31_io_out_id_0;
	wire _mesh_31_31_io_out_last_0;
	wire _mesh_31_31_io_out_valid_0;
	wire [31:0] _mesh_31_30_io_out_a_0;
	wire [31:0] _mesh_31_30_io_out_c_0;
	wire [31:0] _mesh_31_30_io_out_b_0;
	wire _mesh_31_30_io_out_control_0_dataflow;
	wire _mesh_31_30_io_out_control_0_propagate;
	wire [4:0] _mesh_31_30_io_out_control_0_shift;
	wire [2:0] _mesh_31_30_io_out_id_0;
	wire _mesh_31_30_io_out_last_0;
	wire _mesh_31_30_io_out_valid_0;
	wire [31:0] _mesh_31_29_io_out_a_0;
	wire [31:0] _mesh_31_29_io_out_c_0;
	wire [31:0] _mesh_31_29_io_out_b_0;
	wire _mesh_31_29_io_out_control_0_dataflow;
	wire _mesh_31_29_io_out_control_0_propagate;
	wire [4:0] _mesh_31_29_io_out_control_0_shift;
	wire [2:0] _mesh_31_29_io_out_id_0;
	wire _mesh_31_29_io_out_last_0;
	wire _mesh_31_29_io_out_valid_0;
	wire [31:0] _mesh_31_28_io_out_a_0;
	wire [31:0] _mesh_31_28_io_out_c_0;
	wire [31:0] _mesh_31_28_io_out_b_0;
	wire _mesh_31_28_io_out_control_0_dataflow;
	wire _mesh_31_28_io_out_control_0_propagate;
	wire [4:0] _mesh_31_28_io_out_control_0_shift;
	wire [2:0] _mesh_31_28_io_out_id_0;
	wire _mesh_31_28_io_out_last_0;
	wire _mesh_31_28_io_out_valid_0;
	wire [31:0] _mesh_31_27_io_out_a_0;
	wire [31:0] _mesh_31_27_io_out_c_0;
	wire [31:0] _mesh_31_27_io_out_b_0;
	wire _mesh_31_27_io_out_control_0_dataflow;
	wire _mesh_31_27_io_out_control_0_propagate;
	wire [4:0] _mesh_31_27_io_out_control_0_shift;
	wire [2:0] _mesh_31_27_io_out_id_0;
	wire _mesh_31_27_io_out_last_0;
	wire _mesh_31_27_io_out_valid_0;
	wire [31:0] _mesh_31_26_io_out_a_0;
	wire [31:0] _mesh_31_26_io_out_c_0;
	wire [31:0] _mesh_31_26_io_out_b_0;
	wire _mesh_31_26_io_out_control_0_dataflow;
	wire _mesh_31_26_io_out_control_0_propagate;
	wire [4:0] _mesh_31_26_io_out_control_0_shift;
	wire [2:0] _mesh_31_26_io_out_id_0;
	wire _mesh_31_26_io_out_last_0;
	wire _mesh_31_26_io_out_valid_0;
	wire [31:0] _mesh_31_25_io_out_a_0;
	wire [31:0] _mesh_31_25_io_out_c_0;
	wire [31:0] _mesh_31_25_io_out_b_0;
	wire _mesh_31_25_io_out_control_0_dataflow;
	wire _mesh_31_25_io_out_control_0_propagate;
	wire [4:0] _mesh_31_25_io_out_control_0_shift;
	wire [2:0] _mesh_31_25_io_out_id_0;
	wire _mesh_31_25_io_out_last_0;
	wire _mesh_31_25_io_out_valid_0;
	wire [31:0] _mesh_31_24_io_out_a_0;
	wire [31:0] _mesh_31_24_io_out_c_0;
	wire [31:0] _mesh_31_24_io_out_b_0;
	wire _mesh_31_24_io_out_control_0_dataflow;
	wire _mesh_31_24_io_out_control_0_propagate;
	wire [4:0] _mesh_31_24_io_out_control_0_shift;
	wire [2:0] _mesh_31_24_io_out_id_0;
	wire _mesh_31_24_io_out_last_0;
	wire _mesh_31_24_io_out_valid_0;
	wire [31:0] _mesh_31_23_io_out_a_0;
	wire [31:0] _mesh_31_23_io_out_c_0;
	wire [31:0] _mesh_31_23_io_out_b_0;
	wire _mesh_31_23_io_out_control_0_dataflow;
	wire _mesh_31_23_io_out_control_0_propagate;
	wire [4:0] _mesh_31_23_io_out_control_0_shift;
	wire [2:0] _mesh_31_23_io_out_id_0;
	wire _mesh_31_23_io_out_last_0;
	wire _mesh_31_23_io_out_valid_0;
	wire [31:0] _mesh_31_22_io_out_a_0;
	wire [31:0] _mesh_31_22_io_out_c_0;
	wire [31:0] _mesh_31_22_io_out_b_0;
	wire _mesh_31_22_io_out_control_0_dataflow;
	wire _mesh_31_22_io_out_control_0_propagate;
	wire [4:0] _mesh_31_22_io_out_control_0_shift;
	wire [2:0] _mesh_31_22_io_out_id_0;
	wire _mesh_31_22_io_out_last_0;
	wire _mesh_31_22_io_out_valid_0;
	wire [31:0] _mesh_31_21_io_out_a_0;
	wire [31:0] _mesh_31_21_io_out_c_0;
	wire [31:0] _mesh_31_21_io_out_b_0;
	wire _mesh_31_21_io_out_control_0_dataflow;
	wire _mesh_31_21_io_out_control_0_propagate;
	wire [4:0] _mesh_31_21_io_out_control_0_shift;
	wire [2:0] _mesh_31_21_io_out_id_0;
	wire _mesh_31_21_io_out_last_0;
	wire _mesh_31_21_io_out_valid_0;
	wire [31:0] _mesh_31_20_io_out_a_0;
	wire [31:0] _mesh_31_20_io_out_c_0;
	wire [31:0] _mesh_31_20_io_out_b_0;
	wire _mesh_31_20_io_out_control_0_dataflow;
	wire _mesh_31_20_io_out_control_0_propagate;
	wire [4:0] _mesh_31_20_io_out_control_0_shift;
	wire [2:0] _mesh_31_20_io_out_id_0;
	wire _mesh_31_20_io_out_last_0;
	wire _mesh_31_20_io_out_valid_0;
	wire [31:0] _mesh_31_19_io_out_a_0;
	wire [31:0] _mesh_31_19_io_out_c_0;
	wire [31:0] _mesh_31_19_io_out_b_0;
	wire _mesh_31_19_io_out_control_0_dataflow;
	wire _mesh_31_19_io_out_control_0_propagate;
	wire [4:0] _mesh_31_19_io_out_control_0_shift;
	wire [2:0] _mesh_31_19_io_out_id_0;
	wire _mesh_31_19_io_out_last_0;
	wire _mesh_31_19_io_out_valid_0;
	wire [31:0] _mesh_31_18_io_out_a_0;
	wire [31:0] _mesh_31_18_io_out_c_0;
	wire [31:0] _mesh_31_18_io_out_b_0;
	wire _mesh_31_18_io_out_control_0_dataflow;
	wire _mesh_31_18_io_out_control_0_propagate;
	wire [4:0] _mesh_31_18_io_out_control_0_shift;
	wire [2:0] _mesh_31_18_io_out_id_0;
	wire _mesh_31_18_io_out_last_0;
	wire _mesh_31_18_io_out_valid_0;
	wire [31:0] _mesh_31_17_io_out_a_0;
	wire [31:0] _mesh_31_17_io_out_c_0;
	wire [31:0] _mesh_31_17_io_out_b_0;
	wire _mesh_31_17_io_out_control_0_dataflow;
	wire _mesh_31_17_io_out_control_0_propagate;
	wire [4:0] _mesh_31_17_io_out_control_0_shift;
	wire [2:0] _mesh_31_17_io_out_id_0;
	wire _mesh_31_17_io_out_last_0;
	wire _mesh_31_17_io_out_valid_0;
	wire [31:0] _mesh_31_16_io_out_a_0;
	wire [31:0] _mesh_31_16_io_out_c_0;
	wire [31:0] _mesh_31_16_io_out_b_0;
	wire _mesh_31_16_io_out_control_0_dataflow;
	wire _mesh_31_16_io_out_control_0_propagate;
	wire [4:0] _mesh_31_16_io_out_control_0_shift;
	wire [2:0] _mesh_31_16_io_out_id_0;
	wire _mesh_31_16_io_out_last_0;
	wire _mesh_31_16_io_out_valid_0;
	wire [31:0] _mesh_31_15_io_out_a_0;
	wire [31:0] _mesh_31_15_io_out_c_0;
	wire [31:0] _mesh_31_15_io_out_b_0;
	wire _mesh_31_15_io_out_control_0_dataflow;
	wire _mesh_31_15_io_out_control_0_propagate;
	wire [4:0] _mesh_31_15_io_out_control_0_shift;
	wire [2:0] _mesh_31_15_io_out_id_0;
	wire _mesh_31_15_io_out_last_0;
	wire _mesh_31_15_io_out_valid_0;
	wire [31:0] _mesh_31_14_io_out_a_0;
	wire [31:0] _mesh_31_14_io_out_c_0;
	wire [31:0] _mesh_31_14_io_out_b_0;
	wire _mesh_31_14_io_out_control_0_dataflow;
	wire _mesh_31_14_io_out_control_0_propagate;
	wire [4:0] _mesh_31_14_io_out_control_0_shift;
	wire [2:0] _mesh_31_14_io_out_id_0;
	wire _mesh_31_14_io_out_last_0;
	wire _mesh_31_14_io_out_valid_0;
	wire [31:0] _mesh_31_13_io_out_a_0;
	wire [31:0] _mesh_31_13_io_out_c_0;
	wire [31:0] _mesh_31_13_io_out_b_0;
	wire _mesh_31_13_io_out_control_0_dataflow;
	wire _mesh_31_13_io_out_control_0_propagate;
	wire [4:0] _mesh_31_13_io_out_control_0_shift;
	wire [2:0] _mesh_31_13_io_out_id_0;
	wire _mesh_31_13_io_out_last_0;
	wire _mesh_31_13_io_out_valid_0;
	wire [31:0] _mesh_31_12_io_out_a_0;
	wire [31:0] _mesh_31_12_io_out_c_0;
	wire [31:0] _mesh_31_12_io_out_b_0;
	wire _mesh_31_12_io_out_control_0_dataflow;
	wire _mesh_31_12_io_out_control_0_propagate;
	wire [4:0] _mesh_31_12_io_out_control_0_shift;
	wire [2:0] _mesh_31_12_io_out_id_0;
	wire _mesh_31_12_io_out_last_0;
	wire _mesh_31_12_io_out_valid_0;
	wire [31:0] _mesh_31_11_io_out_a_0;
	wire [31:0] _mesh_31_11_io_out_c_0;
	wire [31:0] _mesh_31_11_io_out_b_0;
	wire _mesh_31_11_io_out_control_0_dataflow;
	wire _mesh_31_11_io_out_control_0_propagate;
	wire [4:0] _mesh_31_11_io_out_control_0_shift;
	wire [2:0] _mesh_31_11_io_out_id_0;
	wire _mesh_31_11_io_out_last_0;
	wire _mesh_31_11_io_out_valid_0;
	wire [31:0] _mesh_31_10_io_out_a_0;
	wire [31:0] _mesh_31_10_io_out_c_0;
	wire [31:0] _mesh_31_10_io_out_b_0;
	wire _mesh_31_10_io_out_control_0_dataflow;
	wire _mesh_31_10_io_out_control_0_propagate;
	wire [4:0] _mesh_31_10_io_out_control_0_shift;
	wire [2:0] _mesh_31_10_io_out_id_0;
	wire _mesh_31_10_io_out_last_0;
	wire _mesh_31_10_io_out_valid_0;
	wire [31:0] _mesh_31_9_io_out_a_0;
	wire [31:0] _mesh_31_9_io_out_c_0;
	wire [31:0] _mesh_31_9_io_out_b_0;
	wire _mesh_31_9_io_out_control_0_dataflow;
	wire _mesh_31_9_io_out_control_0_propagate;
	wire [4:0] _mesh_31_9_io_out_control_0_shift;
	wire [2:0] _mesh_31_9_io_out_id_0;
	wire _mesh_31_9_io_out_last_0;
	wire _mesh_31_9_io_out_valid_0;
	wire [31:0] _mesh_31_8_io_out_a_0;
	wire [31:0] _mesh_31_8_io_out_c_0;
	wire [31:0] _mesh_31_8_io_out_b_0;
	wire _mesh_31_8_io_out_control_0_dataflow;
	wire _mesh_31_8_io_out_control_0_propagate;
	wire [4:0] _mesh_31_8_io_out_control_0_shift;
	wire [2:0] _mesh_31_8_io_out_id_0;
	wire _mesh_31_8_io_out_last_0;
	wire _mesh_31_8_io_out_valid_0;
	wire [31:0] _mesh_31_7_io_out_a_0;
	wire [31:0] _mesh_31_7_io_out_c_0;
	wire [31:0] _mesh_31_7_io_out_b_0;
	wire _mesh_31_7_io_out_control_0_dataflow;
	wire _mesh_31_7_io_out_control_0_propagate;
	wire [4:0] _mesh_31_7_io_out_control_0_shift;
	wire [2:0] _mesh_31_7_io_out_id_0;
	wire _mesh_31_7_io_out_last_0;
	wire _mesh_31_7_io_out_valid_0;
	wire [31:0] _mesh_31_6_io_out_a_0;
	wire [31:0] _mesh_31_6_io_out_c_0;
	wire [31:0] _mesh_31_6_io_out_b_0;
	wire _mesh_31_6_io_out_control_0_dataflow;
	wire _mesh_31_6_io_out_control_0_propagate;
	wire [4:0] _mesh_31_6_io_out_control_0_shift;
	wire [2:0] _mesh_31_6_io_out_id_0;
	wire _mesh_31_6_io_out_last_0;
	wire _mesh_31_6_io_out_valid_0;
	wire [31:0] _mesh_31_5_io_out_a_0;
	wire [31:0] _mesh_31_5_io_out_c_0;
	wire [31:0] _mesh_31_5_io_out_b_0;
	wire _mesh_31_5_io_out_control_0_dataflow;
	wire _mesh_31_5_io_out_control_0_propagate;
	wire [4:0] _mesh_31_5_io_out_control_0_shift;
	wire [2:0] _mesh_31_5_io_out_id_0;
	wire _mesh_31_5_io_out_last_0;
	wire _mesh_31_5_io_out_valid_0;
	wire [31:0] _mesh_31_4_io_out_a_0;
	wire [31:0] _mesh_31_4_io_out_c_0;
	wire [31:0] _mesh_31_4_io_out_b_0;
	wire _mesh_31_4_io_out_control_0_dataflow;
	wire _mesh_31_4_io_out_control_0_propagate;
	wire [4:0] _mesh_31_4_io_out_control_0_shift;
	wire [2:0] _mesh_31_4_io_out_id_0;
	wire _mesh_31_4_io_out_last_0;
	wire _mesh_31_4_io_out_valid_0;
	wire [31:0] _mesh_31_3_io_out_a_0;
	wire [31:0] _mesh_31_3_io_out_c_0;
	wire [31:0] _mesh_31_3_io_out_b_0;
	wire _mesh_31_3_io_out_control_0_dataflow;
	wire _mesh_31_3_io_out_control_0_propagate;
	wire [4:0] _mesh_31_3_io_out_control_0_shift;
	wire [2:0] _mesh_31_3_io_out_id_0;
	wire _mesh_31_3_io_out_last_0;
	wire _mesh_31_3_io_out_valid_0;
	wire [31:0] _mesh_31_2_io_out_a_0;
	wire [31:0] _mesh_31_2_io_out_c_0;
	wire [31:0] _mesh_31_2_io_out_b_0;
	wire _mesh_31_2_io_out_control_0_dataflow;
	wire _mesh_31_2_io_out_control_0_propagate;
	wire [4:0] _mesh_31_2_io_out_control_0_shift;
	wire [2:0] _mesh_31_2_io_out_id_0;
	wire _mesh_31_2_io_out_last_0;
	wire _mesh_31_2_io_out_valid_0;
	wire [31:0] _mesh_31_1_io_out_a_0;
	wire [31:0] _mesh_31_1_io_out_c_0;
	wire [31:0] _mesh_31_1_io_out_b_0;
	wire _mesh_31_1_io_out_control_0_dataflow;
	wire _mesh_31_1_io_out_control_0_propagate;
	wire [4:0] _mesh_31_1_io_out_control_0_shift;
	wire [2:0] _mesh_31_1_io_out_id_0;
	wire _mesh_31_1_io_out_last_0;
	wire _mesh_31_1_io_out_valid_0;
	wire [31:0] _mesh_31_0_io_out_a_0;
	wire [31:0] _mesh_31_0_io_out_c_0;
	wire [31:0] _mesh_31_0_io_out_b_0;
	wire _mesh_31_0_io_out_control_0_dataflow;
	wire _mesh_31_0_io_out_control_0_propagate;
	wire [4:0] _mesh_31_0_io_out_control_0_shift;
	wire [2:0] _mesh_31_0_io_out_id_0;
	wire _mesh_31_0_io_out_last_0;
	wire _mesh_31_0_io_out_valid_0;
	wire [31:0] _mesh_30_31_io_out_a_0;
	wire [31:0] _mesh_30_31_io_out_c_0;
	wire [31:0] _mesh_30_31_io_out_b_0;
	wire _mesh_30_31_io_out_control_0_dataflow;
	wire _mesh_30_31_io_out_control_0_propagate;
	wire [4:0] _mesh_30_31_io_out_control_0_shift;
	wire [2:0] _mesh_30_31_io_out_id_0;
	wire _mesh_30_31_io_out_last_0;
	wire _mesh_30_31_io_out_valid_0;
	wire [31:0] _mesh_30_30_io_out_a_0;
	wire [31:0] _mesh_30_30_io_out_c_0;
	wire [31:0] _mesh_30_30_io_out_b_0;
	wire _mesh_30_30_io_out_control_0_dataflow;
	wire _mesh_30_30_io_out_control_0_propagate;
	wire [4:0] _mesh_30_30_io_out_control_0_shift;
	wire [2:0] _mesh_30_30_io_out_id_0;
	wire _mesh_30_30_io_out_last_0;
	wire _mesh_30_30_io_out_valid_0;
	wire [31:0] _mesh_30_29_io_out_a_0;
	wire [31:0] _mesh_30_29_io_out_c_0;
	wire [31:0] _mesh_30_29_io_out_b_0;
	wire _mesh_30_29_io_out_control_0_dataflow;
	wire _mesh_30_29_io_out_control_0_propagate;
	wire [4:0] _mesh_30_29_io_out_control_0_shift;
	wire [2:0] _mesh_30_29_io_out_id_0;
	wire _mesh_30_29_io_out_last_0;
	wire _mesh_30_29_io_out_valid_0;
	wire [31:0] _mesh_30_28_io_out_a_0;
	wire [31:0] _mesh_30_28_io_out_c_0;
	wire [31:0] _mesh_30_28_io_out_b_0;
	wire _mesh_30_28_io_out_control_0_dataflow;
	wire _mesh_30_28_io_out_control_0_propagate;
	wire [4:0] _mesh_30_28_io_out_control_0_shift;
	wire [2:0] _mesh_30_28_io_out_id_0;
	wire _mesh_30_28_io_out_last_0;
	wire _mesh_30_28_io_out_valid_0;
	wire [31:0] _mesh_30_27_io_out_a_0;
	wire [31:0] _mesh_30_27_io_out_c_0;
	wire [31:0] _mesh_30_27_io_out_b_0;
	wire _mesh_30_27_io_out_control_0_dataflow;
	wire _mesh_30_27_io_out_control_0_propagate;
	wire [4:0] _mesh_30_27_io_out_control_0_shift;
	wire [2:0] _mesh_30_27_io_out_id_0;
	wire _mesh_30_27_io_out_last_0;
	wire _mesh_30_27_io_out_valid_0;
	wire [31:0] _mesh_30_26_io_out_a_0;
	wire [31:0] _mesh_30_26_io_out_c_0;
	wire [31:0] _mesh_30_26_io_out_b_0;
	wire _mesh_30_26_io_out_control_0_dataflow;
	wire _mesh_30_26_io_out_control_0_propagate;
	wire [4:0] _mesh_30_26_io_out_control_0_shift;
	wire [2:0] _mesh_30_26_io_out_id_0;
	wire _mesh_30_26_io_out_last_0;
	wire _mesh_30_26_io_out_valid_0;
	wire [31:0] _mesh_30_25_io_out_a_0;
	wire [31:0] _mesh_30_25_io_out_c_0;
	wire [31:0] _mesh_30_25_io_out_b_0;
	wire _mesh_30_25_io_out_control_0_dataflow;
	wire _mesh_30_25_io_out_control_0_propagate;
	wire [4:0] _mesh_30_25_io_out_control_0_shift;
	wire [2:0] _mesh_30_25_io_out_id_0;
	wire _mesh_30_25_io_out_last_0;
	wire _mesh_30_25_io_out_valid_0;
	wire [31:0] _mesh_30_24_io_out_a_0;
	wire [31:0] _mesh_30_24_io_out_c_0;
	wire [31:0] _mesh_30_24_io_out_b_0;
	wire _mesh_30_24_io_out_control_0_dataflow;
	wire _mesh_30_24_io_out_control_0_propagate;
	wire [4:0] _mesh_30_24_io_out_control_0_shift;
	wire [2:0] _mesh_30_24_io_out_id_0;
	wire _mesh_30_24_io_out_last_0;
	wire _mesh_30_24_io_out_valid_0;
	wire [31:0] _mesh_30_23_io_out_a_0;
	wire [31:0] _mesh_30_23_io_out_c_0;
	wire [31:0] _mesh_30_23_io_out_b_0;
	wire _mesh_30_23_io_out_control_0_dataflow;
	wire _mesh_30_23_io_out_control_0_propagate;
	wire [4:0] _mesh_30_23_io_out_control_0_shift;
	wire [2:0] _mesh_30_23_io_out_id_0;
	wire _mesh_30_23_io_out_last_0;
	wire _mesh_30_23_io_out_valid_0;
	wire [31:0] _mesh_30_22_io_out_a_0;
	wire [31:0] _mesh_30_22_io_out_c_0;
	wire [31:0] _mesh_30_22_io_out_b_0;
	wire _mesh_30_22_io_out_control_0_dataflow;
	wire _mesh_30_22_io_out_control_0_propagate;
	wire [4:0] _mesh_30_22_io_out_control_0_shift;
	wire [2:0] _mesh_30_22_io_out_id_0;
	wire _mesh_30_22_io_out_last_0;
	wire _mesh_30_22_io_out_valid_0;
	wire [31:0] _mesh_30_21_io_out_a_0;
	wire [31:0] _mesh_30_21_io_out_c_0;
	wire [31:0] _mesh_30_21_io_out_b_0;
	wire _mesh_30_21_io_out_control_0_dataflow;
	wire _mesh_30_21_io_out_control_0_propagate;
	wire [4:0] _mesh_30_21_io_out_control_0_shift;
	wire [2:0] _mesh_30_21_io_out_id_0;
	wire _mesh_30_21_io_out_last_0;
	wire _mesh_30_21_io_out_valid_0;
	wire [31:0] _mesh_30_20_io_out_a_0;
	wire [31:0] _mesh_30_20_io_out_c_0;
	wire [31:0] _mesh_30_20_io_out_b_0;
	wire _mesh_30_20_io_out_control_0_dataflow;
	wire _mesh_30_20_io_out_control_0_propagate;
	wire [4:0] _mesh_30_20_io_out_control_0_shift;
	wire [2:0] _mesh_30_20_io_out_id_0;
	wire _mesh_30_20_io_out_last_0;
	wire _mesh_30_20_io_out_valid_0;
	wire [31:0] _mesh_30_19_io_out_a_0;
	wire [31:0] _mesh_30_19_io_out_c_0;
	wire [31:0] _mesh_30_19_io_out_b_0;
	wire _mesh_30_19_io_out_control_0_dataflow;
	wire _mesh_30_19_io_out_control_0_propagate;
	wire [4:0] _mesh_30_19_io_out_control_0_shift;
	wire [2:0] _mesh_30_19_io_out_id_0;
	wire _mesh_30_19_io_out_last_0;
	wire _mesh_30_19_io_out_valid_0;
	wire [31:0] _mesh_30_18_io_out_a_0;
	wire [31:0] _mesh_30_18_io_out_c_0;
	wire [31:0] _mesh_30_18_io_out_b_0;
	wire _mesh_30_18_io_out_control_0_dataflow;
	wire _mesh_30_18_io_out_control_0_propagate;
	wire [4:0] _mesh_30_18_io_out_control_0_shift;
	wire [2:0] _mesh_30_18_io_out_id_0;
	wire _mesh_30_18_io_out_last_0;
	wire _mesh_30_18_io_out_valid_0;
	wire [31:0] _mesh_30_17_io_out_a_0;
	wire [31:0] _mesh_30_17_io_out_c_0;
	wire [31:0] _mesh_30_17_io_out_b_0;
	wire _mesh_30_17_io_out_control_0_dataflow;
	wire _mesh_30_17_io_out_control_0_propagate;
	wire [4:0] _mesh_30_17_io_out_control_0_shift;
	wire [2:0] _mesh_30_17_io_out_id_0;
	wire _mesh_30_17_io_out_last_0;
	wire _mesh_30_17_io_out_valid_0;
	wire [31:0] _mesh_30_16_io_out_a_0;
	wire [31:0] _mesh_30_16_io_out_c_0;
	wire [31:0] _mesh_30_16_io_out_b_0;
	wire _mesh_30_16_io_out_control_0_dataflow;
	wire _mesh_30_16_io_out_control_0_propagate;
	wire [4:0] _mesh_30_16_io_out_control_0_shift;
	wire [2:0] _mesh_30_16_io_out_id_0;
	wire _mesh_30_16_io_out_last_0;
	wire _mesh_30_16_io_out_valid_0;
	wire [31:0] _mesh_30_15_io_out_a_0;
	wire [31:0] _mesh_30_15_io_out_c_0;
	wire [31:0] _mesh_30_15_io_out_b_0;
	wire _mesh_30_15_io_out_control_0_dataflow;
	wire _mesh_30_15_io_out_control_0_propagate;
	wire [4:0] _mesh_30_15_io_out_control_0_shift;
	wire [2:0] _mesh_30_15_io_out_id_0;
	wire _mesh_30_15_io_out_last_0;
	wire _mesh_30_15_io_out_valid_0;
	wire [31:0] _mesh_30_14_io_out_a_0;
	wire [31:0] _mesh_30_14_io_out_c_0;
	wire [31:0] _mesh_30_14_io_out_b_0;
	wire _mesh_30_14_io_out_control_0_dataflow;
	wire _mesh_30_14_io_out_control_0_propagate;
	wire [4:0] _mesh_30_14_io_out_control_0_shift;
	wire [2:0] _mesh_30_14_io_out_id_0;
	wire _mesh_30_14_io_out_last_0;
	wire _mesh_30_14_io_out_valid_0;
	wire [31:0] _mesh_30_13_io_out_a_0;
	wire [31:0] _mesh_30_13_io_out_c_0;
	wire [31:0] _mesh_30_13_io_out_b_0;
	wire _mesh_30_13_io_out_control_0_dataflow;
	wire _mesh_30_13_io_out_control_0_propagate;
	wire [4:0] _mesh_30_13_io_out_control_0_shift;
	wire [2:0] _mesh_30_13_io_out_id_0;
	wire _mesh_30_13_io_out_last_0;
	wire _mesh_30_13_io_out_valid_0;
	wire [31:0] _mesh_30_12_io_out_a_0;
	wire [31:0] _mesh_30_12_io_out_c_0;
	wire [31:0] _mesh_30_12_io_out_b_0;
	wire _mesh_30_12_io_out_control_0_dataflow;
	wire _mesh_30_12_io_out_control_0_propagate;
	wire [4:0] _mesh_30_12_io_out_control_0_shift;
	wire [2:0] _mesh_30_12_io_out_id_0;
	wire _mesh_30_12_io_out_last_0;
	wire _mesh_30_12_io_out_valid_0;
	wire [31:0] _mesh_30_11_io_out_a_0;
	wire [31:0] _mesh_30_11_io_out_c_0;
	wire [31:0] _mesh_30_11_io_out_b_0;
	wire _mesh_30_11_io_out_control_0_dataflow;
	wire _mesh_30_11_io_out_control_0_propagate;
	wire [4:0] _mesh_30_11_io_out_control_0_shift;
	wire [2:0] _mesh_30_11_io_out_id_0;
	wire _mesh_30_11_io_out_last_0;
	wire _mesh_30_11_io_out_valid_0;
	wire [31:0] _mesh_30_10_io_out_a_0;
	wire [31:0] _mesh_30_10_io_out_c_0;
	wire [31:0] _mesh_30_10_io_out_b_0;
	wire _mesh_30_10_io_out_control_0_dataflow;
	wire _mesh_30_10_io_out_control_0_propagate;
	wire [4:0] _mesh_30_10_io_out_control_0_shift;
	wire [2:0] _mesh_30_10_io_out_id_0;
	wire _mesh_30_10_io_out_last_0;
	wire _mesh_30_10_io_out_valid_0;
	wire [31:0] _mesh_30_9_io_out_a_0;
	wire [31:0] _mesh_30_9_io_out_c_0;
	wire [31:0] _mesh_30_9_io_out_b_0;
	wire _mesh_30_9_io_out_control_0_dataflow;
	wire _mesh_30_9_io_out_control_0_propagate;
	wire [4:0] _mesh_30_9_io_out_control_0_shift;
	wire [2:0] _mesh_30_9_io_out_id_0;
	wire _mesh_30_9_io_out_last_0;
	wire _mesh_30_9_io_out_valid_0;
	wire [31:0] _mesh_30_8_io_out_a_0;
	wire [31:0] _mesh_30_8_io_out_c_0;
	wire [31:0] _mesh_30_8_io_out_b_0;
	wire _mesh_30_8_io_out_control_0_dataflow;
	wire _mesh_30_8_io_out_control_0_propagate;
	wire [4:0] _mesh_30_8_io_out_control_0_shift;
	wire [2:0] _mesh_30_8_io_out_id_0;
	wire _mesh_30_8_io_out_last_0;
	wire _mesh_30_8_io_out_valid_0;
	wire [31:0] _mesh_30_7_io_out_a_0;
	wire [31:0] _mesh_30_7_io_out_c_0;
	wire [31:0] _mesh_30_7_io_out_b_0;
	wire _mesh_30_7_io_out_control_0_dataflow;
	wire _mesh_30_7_io_out_control_0_propagate;
	wire [4:0] _mesh_30_7_io_out_control_0_shift;
	wire [2:0] _mesh_30_7_io_out_id_0;
	wire _mesh_30_7_io_out_last_0;
	wire _mesh_30_7_io_out_valid_0;
	wire [31:0] _mesh_30_6_io_out_a_0;
	wire [31:0] _mesh_30_6_io_out_c_0;
	wire [31:0] _mesh_30_6_io_out_b_0;
	wire _mesh_30_6_io_out_control_0_dataflow;
	wire _mesh_30_6_io_out_control_0_propagate;
	wire [4:0] _mesh_30_6_io_out_control_0_shift;
	wire [2:0] _mesh_30_6_io_out_id_0;
	wire _mesh_30_6_io_out_last_0;
	wire _mesh_30_6_io_out_valid_0;
	wire [31:0] _mesh_30_5_io_out_a_0;
	wire [31:0] _mesh_30_5_io_out_c_0;
	wire [31:0] _mesh_30_5_io_out_b_0;
	wire _mesh_30_5_io_out_control_0_dataflow;
	wire _mesh_30_5_io_out_control_0_propagate;
	wire [4:0] _mesh_30_5_io_out_control_0_shift;
	wire [2:0] _mesh_30_5_io_out_id_0;
	wire _mesh_30_5_io_out_last_0;
	wire _mesh_30_5_io_out_valid_0;
	wire [31:0] _mesh_30_4_io_out_a_0;
	wire [31:0] _mesh_30_4_io_out_c_0;
	wire [31:0] _mesh_30_4_io_out_b_0;
	wire _mesh_30_4_io_out_control_0_dataflow;
	wire _mesh_30_4_io_out_control_0_propagate;
	wire [4:0] _mesh_30_4_io_out_control_0_shift;
	wire [2:0] _mesh_30_4_io_out_id_0;
	wire _mesh_30_4_io_out_last_0;
	wire _mesh_30_4_io_out_valid_0;
	wire [31:0] _mesh_30_3_io_out_a_0;
	wire [31:0] _mesh_30_3_io_out_c_0;
	wire [31:0] _mesh_30_3_io_out_b_0;
	wire _mesh_30_3_io_out_control_0_dataflow;
	wire _mesh_30_3_io_out_control_0_propagate;
	wire [4:0] _mesh_30_3_io_out_control_0_shift;
	wire [2:0] _mesh_30_3_io_out_id_0;
	wire _mesh_30_3_io_out_last_0;
	wire _mesh_30_3_io_out_valid_0;
	wire [31:0] _mesh_30_2_io_out_a_0;
	wire [31:0] _mesh_30_2_io_out_c_0;
	wire [31:0] _mesh_30_2_io_out_b_0;
	wire _mesh_30_2_io_out_control_0_dataflow;
	wire _mesh_30_2_io_out_control_0_propagate;
	wire [4:0] _mesh_30_2_io_out_control_0_shift;
	wire [2:0] _mesh_30_2_io_out_id_0;
	wire _mesh_30_2_io_out_last_0;
	wire _mesh_30_2_io_out_valid_0;
	wire [31:0] _mesh_30_1_io_out_a_0;
	wire [31:0] _mesh_30_1_io_out_c_0;
	wire [31:0] _mesh_30_1_io_out_b_0;
	wire _mesh_30_1_io_out_control_0_dataflow;
	wire _mesh_30_1_io_out_control_0_propagate;
	wire [4:0] _mesh_30_1_io_out_control_0_shift;
	wire [2:0] _mesh_30_1_io_out_id_0;
	wire _mesh_30_1_io_out_last_0;
	wire _mesh_30_1_io_out_valid_0;
	wire [31:0] _mesh_30_0_io_out_a_0;
	wire [31:0] _mesh_30_0_io_out_c_0;
	wire [31:0] _mesh_30_0_io_out_b_0;
	wire _mesh_30_0_io_out_control_0_dataflow;
	wire _mesh_30_0_io_out_control_0_propagate;
	wire [4:0] _mesh_30_0_io_out_control_0_shift;
	wire [2:0] _mesh_30_0_io_out_id_0;
	wire _mesh_30_0_io_out_last_0;
	wire _mesh_30_0_io_out_valid_0;
	wire [31:0] _mesh_29_31_io_out_a_0;
	wire [31:0] _mesh_29_31_io_out_c_0;
	wire [31:0] _mesh_29_31_io_out_b_0;
	wire _mesh_29_31_io_out_control_0_dataflow;
	wire _mesh_29_31_io_out_control_0_propagate;
	wire [4:0] _mesh_29_31_io_out_control_0_shift;
	wire [2:0] _mesh_29_31_io_out_id_0;
	wire _mesh_29_31_io_out_last_0;
	wire _mesh_29_31_io_out_valid_0;
	wire [31:0] _mesh_29_30_io_out_a_0;
	wire [31:0] _mesh_29_30_io_out_c_0;
	wire [31:0] _mesh_29_30_io_out_b_0;
	wire _mesh_29_30_io_out_control_0_dataflow;
	wire _mesh_29_30_io_out_control_0_propagate;
	wire [4:0] _mesh_29_30_io_out_control_0_shift;
	wire [2:0] _mesh_29_30_io_out_id_0;
	wire _mesh_29_30_io_out_last_0;
	wire _mesh_29_30_io_out_valid_0;
	wire [31:0] _mesh_29_29_io_out_a_0;
	wire [31:0] _mesh_29_29_io_out_c_0;
	wire [31:0] _mesh_29_29_io_out_b_0;
	wire _mesh_29_29_io_out_control_0_dataflow;
	wire _mesh_29_29_io_out_control_0_propagate;
	wire [4:0] _mesh_29_29_io_out_control_0_shift;
	wire [2:0] _mesh_29_29_io_out_id_0;
	wire _mesh_29_29_io_out_last_0;
	wire _mesh_29_29_io_out_valid_0;
	wire [31:0] _mesh_29_28_io_out_a_0;
	wire [31:0] _mesh_29_28_io_out_c_0;
	wire [31:0] _mesh_29_28_io_out_b_0;
	wire _mesh_29_28_io_out_control_0_dataflow;
	wire _mesh_29_28_io_out_control_0_propagate;
	wire [4:0] _mesh_29_28_io_out_control_0_shift;
	wire [2:0] _mesh_29_28_io_out_id_0;
	wire _mesh_29_28_io_out_last_0;
	wire _mesh_29_28_io_out_valid_0;
	wire [31:0] _mesh_29_27_io_out_a_0;
	wire [31:0] _mesh_29_27_io_out_c_0;
	wire [31:0] _mesh_29_27_io_out_b_0;
	wire _mesh_29_27_io_out_control_0_dataflow;
	wire _mesh_29_27_io_out_control_0_propagate;
	wire [4:0] _mesh_29_27_io_out_control_0_shift;
	wire [2:0] _mesh_29_27_io_out_id_0;
	wire _mesh_29_27_io_out_last_0;
	wire _mesh_29_27_io_out_valid_0;
	wire [31:0] _mesh_29_26_io_out_a_0;
	wire [31:0] _mesh_29_26_io_out_c_0;
	wire [31:0] _mesh_29_26_io_out_b_0;
	wire _mesh_29_26_io_out_control_0_dataflow;
	wire _mesh_29_26_io_out_control_0_propagate;
	wire [4:0] _mesh_29_26_io_out_control_0_shift;
	wire [2:0] _mesh_29_26_io_out_id_0;
	wire _mesh_29_26_io_out_last_0;
	wire _mesh_29_26_io_out_valid_0;
	wire [31:0] _mesh_29_25_io_out_a_0;
	wire [31:0] _mesh_29_25_io_out_c_0;
	wire [31:0] _mesh_29_25_io_out_b_0;
	wire _mesh_29_25_io_out_control_0_dataflow;
	wire _mesh_29_25_io_out_control_0_propagate;
	wire [4:0] _mesh_29_25_io_out_control_0_shift;
	wire [2:0] _mesh_29_25_io_out_id_0;
	wire _mesh_29_25_io_out_last_0;
	wire _mesh_29_25_io_out_valid_0;
	wire [31:0] _mesh_29_24_io_out_a_0;
	wire [31:0] _mesh_29_24_io_out_c_0;
	wire [31:0] _mesh_29_24_io_out_b_0;
	wire _mesh_29_24_io_out_control_0_dataflow;
	wire _mesh_29_24_io_out_control_0_propagate;
	wire [4:0] _mesh_29_24_io_out_control_0_shift;
	wire [2:0] _mesh_29_24_io_out_id_0;
	wire _mesh_29_24_io_out_last_0;
	wire _mesh_29_24_io_out_valid_0;
	wire [31:0] _mesh_29_23_io_out_a_0;
	wire [31:0] _mesh_29_23_io_out_c_0;
	wire [31:0] _mesh_29_23_io_out_b_0;
	wire _mesh_29_23_io_out_control_0_dataflow;
	wire _mesh_29_23_io_out_control_0_propagate;
	wire [4:0] _mesh_29_23_io_out_control_0_shift;
	wire [2:0] _mesh_29_23_io_out_id_0;
	wire _mesh_29_23_io_out_last_0;
	wire _mesh_29_23_io_out_valid_0;
	wire [31:0] _mesh_29_22_io_out_a_0;
	wire [31:0] _mesh_29_22_io_out_c_0;
	wire [31:0] _mesh_29_22_io_out_b_0;
	wire _mesh_29_22_io_out_control_0_dataflow;
	wire _mesh_29_22_io_out_control_0_propagate;
	wire [4:0] _mesh_29_22_io_out_control_0_shift;
	wire [2:0] _mesh_29_22_io_out_id_0;
	wire _mesh_29_22_io_out_last_0;
	wire _mesh_29_22_io_out_valid_0;
	wire [31:0] _mesh_29_21_io_out_a_0;
	wire [31:0] _mesh_29_21_io_out_c_0;
	wire [31:0] _mesh_29_21_io_out_b_0;
	wire _mesh_29_21_io_out_control_0_dataflow;
	wire _mesh_29_21_io_out_control_0_propagate;
	wire [4:0] _mesh_29_21_io_out_control_0_shift;
	wire [2:0] _mesh_29_21_io_out_id_0;
	wire _mesh_29_21_io_out_last_0;
	wire _mesh_29_21_io_out_valid_0;
	wire [31:0] _mesh_29_20_io_out_a_0;
	wire [31:0] _mesh_29_20_io_out_c_0;
	wire [31:0] _mesh_29_20_io_out_b_0;
	wire _mesh_29_20_io_out_control_0_dataflow;
	wire _mesh_29_20_io_out_control_0_propagate;
	wire [4:0] _mesh_29_20_io_out_control_0_shift;
	wire [2:0] _mesh_29_20_io_out_id_0;
	wire _mesh_29_20_io_out_last_0;
	wire _mesh_29_20_io_out_valid_0;
	wire [31:0] _mesh_29_19_io_out_a_0;
	wire [31:0] _mesh_29_19_io_out_c_0;
	wire [31:0] _mesh_29_19_io_out_b_0;
	wire _mesh_29_19_io_out_control_0_dataflow;
	wire _mesh_29_19_io_out_control_0_propagate;
	wire [4:0] _mesh_29_19_io_out_control_0_shift;
	wire [2:0] _mesh_29_19_io_out_id_0;
	wire _mesh_29_19_io_out_last_0;
	wire _mesh_29_19_io_out_valid_0;
	wire [31:0] _mesh_29_18_io_out_a_0;
	wire [31:0] _mesh_29_18_io_out_c_0;
	wire [31:0] _mesh_29_18_io_out_b_0;
	wire _mesh_29_18_io_out_control_0_dataflow;
	wire _mesh_29_18_io_out_control_0_propagate;
	wire [4:0] _mesh_29_18_io_out_control_0_shift;
	wire [2:0] _mesh_29_18_io_out_id_0;
	wire _mesh_29_18_io_out_last_0;
	wire _mesh_29_18_io_out_valid_0;
	wire [31:0] _mesh_29_17_io_out_a_0;
	wire [31:0] _mesh_29_17_io_out_c_0;
	wire [31:0] _mesh_29_17_io_out_b_0;
	wire _mesh_29_17_io_out_control_0_dataflow;
	wire _mesh_29_17_io_out_control_0_propagate;
	wire [4:0] _mesh_29_17_io_out_control_0_shift;
	wire [2:0] _mesh_29_17_io_out_id_0;
	wire _mesh_29_17_io_out_last_0;
	wire _mesh_29_17_io_out_valid_0;
	wire [31:0] _mesh_29_16_io_out_a_0;
	wire [31:0] _mesh_29_16_io_out_c_0;
	wire [31:0] _mesh_29_16_io_out_b_0;
	wire _mesh_29_16_io_out_control_0_dataflow;
	wire _mesh_29_16_io_out_control_0_propagate;
	wire [4:0] _mesh_29_16_io_out_control_0_shift;
	wire [2:0] _mesh_29_16_io_out_id_0;
	wire _mesh_29_16_io_out_last_0;
	wire _mesh_29_16_io_out_valid_0;
	wire [31:0] _mesh_29_15_io_out_a_0;
	wire [31:0] _mesh_29_15_io_out_c_0;
	wire [31:0] _mesh_29_15_io_out_b_0;
	wire _mesh_29_15_io_out_control_0_dataflow;
	wire _mesh_29_15_io_out_control_0_propagate;
	wire [4:0] _mesh_29_15_io_out_control_0_shift;
	wire [2:0] _mesh_29_15_io_out_id_0;
	wire _mesh_29_15_io_out_last_0;
	wire _mesh_29_15_io_out_valid_0;
	wire [31:0] _mesh_29_14_io_out_a_0;
	wire [31:0] _mesh_29_14_io_out_c_0;
	wire [31:0] _mesh_29_14_io_out_b_0;
	wire _mesh_29_14_io_out_control_0_dataflow;
	wire _mesh_29_14_io_out_control_0_propagate;
	wire [4:0] _mesh_29_14_io_out_control_0_shift;
	wire [2:0] _mesh_29_14_io_out_id_0;
	wire _mesh_29_14_io_out_last_0;
	wire _mesh_29_14_io_out_valid_0;
	wire [31:0] _mesh_29_13_io_out_a_0;
	wire [31:0] _mesh_29_13_io_out_c_0;
	wire [31:0] _mesh_29_13_io_out_b_0;
	wire _mesh_29_13_io_out_control_0_dataflow;
	wire _mesh_29_13_io_out_control_0_propagate;
	wire [4:0] _mesh_29_13_io_out_control_0_shift;
	wire [2:0] _mesh_29_13_io_out_id_0;
	wire _mesh_29_13_io_out_last_0;
	wire _mesh_29_13_io_out_valid_0;
	wire [31:0] _mesh_29_12_io_out_a_0;
	wire [31:0] _mesh_29_12_io_out_c_0;
	wire [31:0] _mesh_29_12_io_out_b_0;
	wire _mesh_29_12_io_out_control_0_dataflow;
	wire _mesh_29_12_io_out_control_0_propagate;
	wire [4:0] _mesh_29_12_io_out_control_0_shift;
	wire [2:0] _mesh_29_12_io_out_id_0;
	wire _mesh_29_12_io_out_last_0;
	wire _mesh_29_12_io_out_valid_0;
	wire [31:0] _mesh_29_11_io_out_a_0;
	wire [31:0] _mesh_29_11_io_out_c_0;
	wire [31:0] _mesh_29_11_io_out_b_0;
	wire _mesh_29_11_io_out_control_0_dataflow;
	wire _mesh_29_11_io_out_control_0_propagate;
	wire [4:0] _mesh_29_11_io_out_control_0_shift;
	wire [2:0] _mesh_29_11_io_out_id_0;
	wire _mesh_29_11_io_out_last_0;
	wire _mesh_29_11_io_out_valid_0;
	wire [31:0] _mesh_29_10_io_out_a_0;
	wire [31:0] _mesh_29_10_io_out_c_0;
	wire [31:0] _mesh_29_10_io_out_b_0;
	wire _mesh_29_10_io_out_control_0_dataflow;
	wire _mesh_29_10_io_out_control_0_propagate;
	wire [4:0] _mesh_29_10_io_out_control_0_shift;
	wire [2:0] _mesh_29_10_io_out_id_0;
	wire _mesh_29_10_io_out_last_0;
	wire _mesh_29_10_io_out_valid_0;
	wire [31:0] _mesh_29_9_io_out_a_0;
	wire [31:0] _mesh_29_9_io_out_c_0;
	wire [31:0] _mesh_29_9_io_out_b_0;
	wire _mesh_29_9_io_out_control_0_dataflow;
	wire _mesh_29_9_io_out_control_0_propagate;
	wire [4:0] _mesh_29_9_io_out_control_0_shift;
	wire [2:0] _mesh_29_9_io_out_id_0;
	wire _mesh_29_9_io_out_last_0;
	wire _mesh_29_9_io_out_valid_0;
	wire [31:0] _mesh_29_8_io_out_a_0;
	wire [31:0] _mesh_29_8_io_out_c_0;
	wire [31:0] _mesh_29_8_io_out_b_0;
	wire _mesh_29_8_io_out_control_0_dataflow;
	wire _mesh_29_8_io_out_control_0_propagate;
	wire [4:0] _mesh_29_8_io_out_control_0_shift;
	wire [2:0] _mesh_29_8_io_out_id_0;
	wire _mesh_29_8_io_out_last_0;
	wire _mesh_29_8_io_out_valid_0;
	wire [31:0] _mesh_29_7_io_out_a_0;
	wire [31:0] _mesh_29_7_io_out_c_0;
	wire [31:0] _mesh_29_7_io_out_b_0;
	wire _mesh_29_7_io_out_control_0_dataflow;
	wire _mesh_29_7_io_out_control_0_propagate;
	wire [4:0] _mesh_29_7_io_out_control_0_shift;
	wire [2:0] _mesh_29_7_io_out_id_0;
	wire _mesh_29_7_io_out_last_0;
	wire _mesh_29_7_io_out_valid_0;
	wire [31:0] _mesh_29_6_io_out_a_0;
	wire [31:0] _mesh_29_6_io_out_c_0;
	wire [31:0] _mesh_29_6_io_out_b_0;
	wire _mesh_29_6_io_out_control_0_dataflow;
	wire _mesh_29_6_io_out_control_0_propagate;
	wire [4:0] _mesh_29_6_io_out_control_0_shift;
	wire [2:0] _mesh_29_6_io_out_id_0;
	wire _mesh_29_6_io_out_last_0;
	wire _mesh_29_6_io_out_valid_0;
	wire [31:0] _mesh_29_5_io_out_a_0;
	wire [31:0] _mesh_29_5_io_out_c_0;
	wire [31:0] _mesh_29_5_io_out_b_0;
	wire _mesh_29_5_io_out_control_0_dataflow;
	wire _mesh_29_5_io_out_control_0_propagate;
	wire [4:0] _mesh_29_5_io_out_control_0_shift;
	wire [2:0] _mesh_29_5_io_out_id_0;
	wire _mesh_29_5_io_out_last_0;
	wire _mesh_29_5_io_out_valid_0;
	wire [31:0] _mesh_29_4_io_out_a_0;
	wire [31:0] _mesh_29_4_io_out_c_0;
	wire [31:0] _mesh_29_4_io_out_b_0;
	wire _mesh_29_4_io_out_control_0_dataflow;
	wire _mesh_29_4_io_out_control_0_propagate;
	wire [4:0] _mesh_29_4_io_out_control_0_shift;
	wire [2:0] _mesh_29_4_io_out_id_0;
	wire _mesh_29_4_io_out_last_0;
	wire _mesh_29_4_io_out_valid_0;
	wire [31:0] _mesh_29_3_io_out_a_0;
	wire [31:0] _mesh_29_3_io_out_c_0;
	wire [31:0] _mesh_29_3_io_out_b_0;
	wire _mesh_29_3_io_out_control_0_dataflow;
	wire _mesh_29_3_io_out_control_0_propagate;
	wire [4:0] _mesh_29_3_io_out_control_0_shift;
	wire [2:0] _mesh_29_3_io_out_id_0;
	wire _mesh_29_3_io_out_last_0;
	wire _mesh_29_3_io_out_valid_0;
	wire [31:0] _mesh_29_2_io_out_a_0;
	wire [31:0] _mesh_29_2_io_out_c_0;
	wire [31:0] _mesh_29_2_io_out_b_0;
	wire _mesh_29_2_io_out_control_0_dataflow;
	wire _mesh_29_2_io_out_control_0_propagate;
	wire [4:0] _mesh_29_2_io_out_control_0_shift;
	wire [2:0] _mesh_29_2_io_out_id_0;
	wire _mesh_29_2_io_out_last_0;
	wire _mesh_29_2_io_out_valid_0;
	wire [31:0] _mesh_29_1_io_out_a_0;
	wire [31:0] _mesh_29_1_io_out_c_0;
	wire [31:0] _mesh_29_1_io_out_b_0;
	wire _mesh_29_1_io_out_control_0_dataflow;
	wire _mesh_29_1_io_out_control_0_propagate;
	wire [4:0] _mesh_29_1_io_out_control_0_shift;
	wire [2:0] _mesh_29_1_io_out_id_0;
	wire _mesh_29_1_io_out_last_0;
	wire _mesh_29_1_io_out_valid_0;
	wire [31:0] _mesh_29_0_io_out_a_0;
	wire [31:0] _mesh_29_0_io_out_c_0;
	wire [31:0] _mesh_29_0_io_out_b_0;
	wire _mesh_29_0_io_out_control_0_dataflow;
	wire _mesh_29_0_io_out_control_0_propagate;
	wire [4:0] _mesh_29_0_io_out_control_0_shift;
	wire [2:0] _mesh_29_0_io_out_id_0;
	wire _mesh_29_0_io_out_last_0;
	wire _mesh_29_0_io_out_valid_0;
	wire [31:0] _mesh_28_31_io_out_a_0;
	wire [31:0] _mesh_28_31_io_out_c_0;
	wire [31:0] _mesh_28_31_io_out_b_0;
	wire _mesh_28_31_io_out_control_0_dataflow;
	wire _mesh_28_31_io_out_control_0_propagate;
	wire [4:0] _mesh_28_31_io_out_control_0_shift;
	wire [2:0] _mesh_28_31_io_out_id_0;
	wire _mesh_28_31_io_out_last_0;
	wire _mesh_28_31_io_out_valid_0;
	wire [31:0] _mesh_28_30_io_out_a_0;
	wire [31:0] _mesh_28_30_io_out_c_0;
	wire [31:0] _mesh_28_30_io_out_b_0;
	wire _mesh_28_30_io_out_control_0_dataflow;
	wire _mesh_28_30_io_out_control_0_propagate;
	wire [4:0] _mesh_28_30_io_out_control_0_shift;
	wire [2:0] _mesh_28_30_io_out_id_0;
	wire _mesh_28_30_io_out_last_0;
	wire _mesh_28_30_io_out_valid_0;
	wire [31:0] _mesh_28_29_io_out_a_0;
	wire [31:0] _mesh_28_29_io_out_c_0;
	wire [31:0] _mesh_28_29_io_out_b_0;
	wire _mesh_28_29_io_out_control_0_dataflow;
	wire _mesh_28_29_io_out_control_0_propagate;
	wire [4:0] _mesh_28_29_io_out_control_0_shift;
	wire [2:0] _mesh_28_29_io_out_id_0;
	wire _mesh_28_29_io_out_last_0;
	wire _mesh_28_29_io_out_valid_0;
	wire [31:0] _mesh_28_28_io_out_a_0;
	wire [31:0] _mesh_28_28_io_out_c_0;
	wire [31:0] _mesh_28_28_io_out_b_0;
	wire _mesh_28_28_io_out_control_0_dataflow;
	wire _mesh_28_28_io_out_control_0_propagate;
	wire [4:0] _mesh_28_28_io_out_control_0_shift;
	wire [2:0] _mesh_28_28_io_out_id_0;
	wire _mesh_28_28_io_out_last_0;
	wire _mesh_28_28_io_out_valid_0;
	wire [31:0] _mesh_28_27_io_out_a_0;
	wire [31:0] _mesh_28_27_io_out_c_0;
	wire [31:0] _mesh_28_27_io_out_b_0;
	wire _mesh_28_27_io_out_control_0_dataflow;
	wire _mesh_28_27_io_out_control_0_propagate;
	wire [4:0] _mesh_28_27_io_out_control_0_shift;
	wire [2:0] _mesh_28_27_io_out_id_0;
	wire _mesh_28_27_io_out_last_0;
	wire _mesh_28_27_io_out_valid_0;
	wire [31:0] _mesh_28_26_io_out_a_0;
	wire [31:0] _mesh_28_26_io_out_c_0;
	wire [31:0] _mesh_28_26_io_out_b_0;
	wire _mesh_28_26_io_out_control_0_dataflow;
	wire _mesh_28_26_io_out_control_0_propagate;
	wire [4:0] _mesh_28_26_io_out_control_0_shift;
	wire [2:0] _mesh_28_26_io_out_id_0;
	wire _mesh_28_26_io_out_last_0;
	wire _mesh_28_26_io_out_valid_0;
	wire [31:0] _mesh_28_25_io_out_a_0;
	wire [31:0] _mesh_28_25_io_out_c_0;
	wire [31:0] _mesh_28_25_io_out_b_0;
	wire _mesh_28_25_io_out_control_0_dataflow;
	wire _mesh_28_25_io_out_control_0_propagate;
	wire [4:0] _mesh_28_25_io_out_control_0_shift;
	wire [2:0] _mesh_28_25_io_out_id_0;
	wire _mesh_28_25_io_out_last_0;
	wire _mesh_28_25_io_out_valid_0;
	wire [31:0] _mesh_28_24_io_out_a_0;
	wire [31:0] _mesh_28_24_io_out_c_0;
	wire [31:0] _mesh_28_24_io_out_b_0;
	wire _mesh_28_24_io_out_control_0_dataflow;
	wire _mesh_28_24_io_out_control_0_propagate;
	wire [4:0] _mesh_28_24_io_out_control_0_shift;
	wire [2:0] _mesh_28_24_io_out_id_0;
	wire _mesh_28_24_io_out_last_0;
	wire _mesh_28_24_io_out_valid_0;
	wire [31:0] _mesh_28_23_io_out_a_0;
	wire [31:0] _mesh_28_23_io_out_c_0;
	wire [31:0] _mesh_28_23_io_out_b_0;
	wire _mesh_28_23_io_out_control_0_dataflow;
	wire _mesh_28_23_io_out_control_0_propagate;
	wire [4:0] _mesh_28_23_io_out_control_0_shift;
	wire [2:0] _mesh_28_23_io_out_id_0;
	wire _mesh_28_23_io_out_last_0;
	wire _mesh_28_23_io_out_valid_0;
	wire [31:0] _mesh_28_22_io_out_a_0;
	wire [31:0] _mesh_28_22_io_out_c_0;
	wire [31:0] _mesh_28_22_io_out_b_0;
	wire _mesh_28_22_io_out_control_0_dataflow;
	wire _mesh_28_22_io_out_control_0_propagate;
	wire [4:0] _mesh_28_22_io_out_control_0_shift;
	wire [2:0] _mesh_28_22_io_out_id_0;
	wire _mesh_28_22_io_out_last_0;
	wire _mesh_28_22_io_out_valid_0;
	wire [31:0] _mesh_28_21_io_out_a_0;
	wire [31:0] _mesh_28_21_io_out_c_0;
	wire [31:0] _mesh_28_21_io_out_b_0;
	wire _mesh_28_21_io_out_control_0_dataflow;
	wire _mesh_28_21_io_out_control_0_propagate;
	wire [4:0] _mesh_28_21_io_out_control_0_shift;
	wire [2:0] _mesh_28_21_io_out_id_0;
	wire _mesh_28_21_io_out_last_0;
	wire _mesh_28_21_io_out_valid_0;
	wire [31:0] _mesh_28_20_io_out_a_0;
	wire [31:0] _mesh_28_20_io_out_c_0;
	wire [31:0] _mesh_28_20_io_out_b_0;
	wire _mesh_28_20_io_out_control_0_dataflow;
	wire _mesh_28_20_io_out_control_0_propagate;
	wire [4:0] _mesh_28_20_io_out_control_0_shift;
	wire [2:0] _mesh_28_20_io_out_id_0;
	wire _mesh_28_20_io_out_last_0;
	wire _mesh_28_20_io_out_valid_0;
	wire [31:0] _mesh_28_19_io_out_a_0;
	wire [31:0] _mesh_28_19_io_out_c_0;
	wire [31:0] _mesh_28_19_io_out_b_0;
	wire _mesh_28_19_io_out_control_0_dataflow;
	wire _mesh_28_19_io_out_control_0_propagate;
	wire [4:0] _mesh_28_19_io_out_control_0_shift;
	wire [2:0] _mesh_28_19_io_out_id_0;
	wire _mesh_28_19_io_out_last_0;
	wire _mesh_28_19_io_out_valid_0;
	wire [31:0] _mesh_28_18_io_out_a_0;
	wire [31:0] _mesh_28_18_io_out_c_0;
	wire [31:0] _mesh_28_18_io_out_b_0;
	wire _mesh_28_18_io_out_control_0_dataflow;
	wire _mesh_28_18_io_out_control_0_propagate;
	wire [4:0] _mesh_28_18_io_out_control_0_shift;
	wire [2:0] _mesh_28_18_io_out_id_0;
	wire _mesh_28_18_io_out_last_0;
	wire _mesh_28_18_io_out_valid_0;
	wire [31:0] _mesh_28_17_io_out_a_0;
	wire [31:0] _mesh_28_17_io_out_c_0;
	wire [31:0] _mesh_28_17_io_out_b_0;
	wire _mesh_28_17_io_out_control_0_dataflow;
	wire _mesh_28_17_io_out_control_0_propagate;
	wire [4:0] _mesh_28_17_io_out_control_0_shift;
	wire [2:0] _mesh_28_17_io_out_id_0;
	wire _mesh_28_17_io_out_last_0;
	wire _mesh_28_17_io_out_valid_0;
	wire [31:0] _mesh_28_16_io_out_a_0;
	wire [31:0] _mesh_28_16_io_out_c_0;
	wire [31:0] _mesh_28_16_io_out_b_0;
	wire _mesh_28_16_io_out_control_0_dataflow;
	wire _mesh_28_16_io_out_control_0_propagate;
	wire [4:0] _mesh_28_16_io_out_control_0_shift;
	wire [2:0] _mesh_28_16_io_out_id_0;
	wire _mesh_28_16_io_out_last_0;
	wire _mesh_28_16_io_out_valid_0;
	wire [31:0] _mesh_28_15_io_out_a_0;
	wire [31:0] _mesh_28_15_io_out_c_0;
	wire [31:0] _mesh_28_15_io_out_b_0;
	wire _mesh_28_15_io_out_control_0_dataflow;
	wire _mesh_28_15_io_out_control_0_propagate;
	wire [4:0] _mesh_28_15_io_out_control_0_shift;
	wire [2:0] _mesh_28_15_io_out_id_0;
	wire _mesh_28_15_io_out_last_0;
	wire _mesh_28_15_io_out_valid_0;
	wire [31:0] _mesh_28_14_io_out_a_0;
	wire [31:0] _mesh_28_14_io_out_c_0;
	wire [31:0] _mesh_28_14_io_out_b_0;
	wire _mesh_28_14_io_out_control_0_dataflow;
	wire _mesh_28_14_io_out_control_0_propagate;
	wire [4:0] _mesh_28_14_io_out_control_0_shift;
	wire [2:0] _mesh_28_14_io_out_id_0;
	wire _mesh_28_14_io_out_last_0;
	wire _mesh_28_14_io_out_valid_0;
	wire [31:0] _mesh_28_13_io_out_a_0;
	wire [31:0] _mesh_28_13_io_out_c_0;
	wire [31:0] _mesh_28_13_io_out_b_0;
	wire _mesh_28_13_io_out_control_0_dataflow;
	wire _mesh_28_13_io_out_control_0_propagate;
	wire [4:0] _mesh_28_13_io_out_control_0_shift;
	wire [2:0] _mesh_28_13_io_out_id_0;
	wire _mesh_28_13_io_out_last_0;
	wire _mesh_28_13_io_out_valid_0;
	wire [31:0] _mesh_28_12_io_out_a_0;
	wire [31:0] _mesh_28_12_io_out_c_0;
	wire [31:0] _mesh_28_12_io_out_b_0;
	wire _mesh_28_12_io_out_control_0_dataflow;
	wire _mesh_28_12_io_out_control_0_propagate;
	wire [4:0] _mesh_28_12_io_out_control_0_shift;
	wire [2:0] _mesh_28_12_io_out_id_0;
	wire _mesh_28_12_io_out_last_0;
	wire _mesh_28_12_io_out_valid_0;
	wire [31:0] _mesh_28_11_io_out_a_0;
	wire [31:0] _mesh_28_11_io_out_c_0;
	wire [31:0] _mesh_28_11_io_out_b_0;
	wire _mesh_28_11_io_out_control_0_dataflow;
	wire _mesh_28_11_io_out_control_0_propagate;
	wire [4:0] _mesh_28_11_io_out_control_0_shift;
	wire [2:0] _mesh_28_11_io_out_id_0;
	wire _mesh_28_11_io_out_last_0;
	wire _mesh_28_11_io_out_valid_0;
	wire [31:0] _mesh_28_10_io_out_a_0;
	wire [31:0] _mesh_28_10_io_out_c_0;
	wire [31:0] _mesh_28_10_io_out_b_0;
	wire _mesh_28_10_io_out_control_0_dataflow;
	wire _mesh_28_10_io_out_control_0_propagate;
	wire [4:0] _mesh_28_10_io_out_control_0_shift;
	wire [2:0] _mesh_28_10_io_out_id_0;
	wire _mesh_28_10_io_out_last_0;
	wire _mesh_28_10_io_out_valid_0;
	wire [31:0] _mesh_28_9_io_out_a_0;
	wire [31:0] _mesh_28_9_io_out_c_0;
	wire [31:0] _mesh_28_9_io_out_b_0;
	wire _mesh_28_9_io_out_control_0_dataflow;
	wire _mesh_28_9_io_out_control_0_propagate;
	wire [4:0] _mesh_28_9_io_out_control_0_shift;
	wire [2:0] _mesh_28_9_io_out_id_0;
	wire _mesh_28_9_io_out_last_0;
	wire _mesh_28_9_io_out_valid_0;
	wire [31:0] _mesh_28_8_io_out_a_0;
	wire [31:0] _mesh_28_8_io_out_c_0;
	wire [31:0] _mesh_28_8_io_out_b_0;
	wire _mesh_28_8_io_out_control_0_dataflow;
	wire _mesh_28_8_io_out_control_0_propagate;
	wire [4:0] _mesh_28_8_io_out_control_0_shift;
	wire [2:0] _mesh_28_8_io_out_id_0;
	wire _mesh_28_8_io_out_last_0;
	wire _mesh_28_8_io_out_valid_0;
	wire [31:0] _mesh_28_7_io_out_a_0;
	wire [31:0] _mesh_28_7_io_out_c_0;
	wire [31:0] _mesh_28_7_io_out_b_0;
	wire _mesh_28_7_io_out_control_0_dataflow;
	wire _mesh_28_7_io_out_control_0_propagate;
	wire [4:0] _mesh_28_7_io_out_control_0_shift;
	wire [2:0] _mesh_28_7_io_out_id_0;
	wire _mesh_28_7_io_out_last_0;
	wire _mesh_28_7_io_out_valid_0;
	wire [31:0] _mesh_28_6_io_out_a_0;
	wire [31:0] _mesh_28_6_io_out_c_0;
	wire [31:0] _mesh_28_6_io_out_b_0;
	wire _mesh_28_6_io_out_control_0_dataflow;
	wire _mesh_28_6_io_out_control_0_propagate;
	wire [4:0] _mesh_28_6_io_out_control_0_shift;
	wire [2:0] _mesh_28_6_io_out_id_0;
	wire _mesh_28_6_io_out_last_0;
	wire _mesh_28_6_io_out_valid_0;
	wire [31:0] _mesh_28_5_io_out_a_0;
	wire [31:0] _mesh_28_5_io_out_c_0;
	wire [31:0] _mesh_28_5_io_out_b_0;
	wire _mesh_28_5_io_out_control_0_dataflow;
	wire _mesh_28_5_io_out_control_0_propagate;
	wire [4:0] _mesh_28_5_io_out_control_0_shift;
	wire [2:0] _mesh_28_5_io_out_id_0;
	wire _mesh_28_5_io_out_last_0;
	wire _mesh_28_5_io_out_valid_0;
	wire [31:0] _mesh_28_4_io_out_a_0;
	wire [31:0] _mesh_28_4_io_out_c_0;
	wire [31:0] _mesh_28_4_io_out_b_0;
	wire _mesh_28_4_io_out_control_0_dataflow;
	wire _mesh_28_4_io_out_control_0_propagate;
	wire [4:0] _mesh_28_4_io_out_control_0_shift;
	wire [2:0] _mesh_28_4_io_out_id_0;
	wire _mesh_28_4_io_out_last_0;
	wire _mesh_28_4_io_out_valid_0;
	wire [31:0] _mesh_28_3_io_out_a_0;
	wire [31:0] _mesh_28_3_io_out_c_0;
	wire [31:0] _mesh_28_3_io_out_b_0;
	wire _mesh_28_3_io_out_control_0_dataflow;
	wire _mesh_28_3_io_out_control_0_propagate;
	wire [4:0] _mesh_28_3_io_out_control_0_shift;
	wire [2:0] _mesh_28_3_io_out_id_0;
	wire _mesh_28_3_io_out_last_0;
	wire _mesh_28_3_io_out_valid_0;
	wire [31:0] _mesh_28_2_io_out_a_0;
	wire [31:0] _mesh_28_2_io_out_c_0;
	wire [31:0] _mesh_28_2_io_out_b_0;
	wire _mesh_28_2_io_out_control_0_dataflow;
	wire _mesh_28_2_io_out_control_0_propagate;
	wire [4:0] _mesh_28_2_io_out_control_0_shift;
	wire [2:0] _mesh_28_2_io_out_id_0;
	wire _mesh_28_2_io_out_last_0;
	wire _mesh_28_2_io_out_valid_0;
	wire [31:0] _mesh_28_1_io_out_a_0;
	wire [31:0] _mesh_28_1_io_out_c_0;
	wire [31:0] _mesh_28_1_io_out_b_0;
	wire _mesh_28_1_io_out_control_0_dataflow;
	wire _mesh_28_1_io_out_control_0_propagate;
	wire [4:0] _mesh_28_1_io_out_control_0_shift;
	wire [2:0] _mesh_28_1_io_out_id_0;
	wire _mesh_28_1_io_out_last_0;
	wire _mesh_28_1_io_out_valid_0;
	wire [31:0] _mesh_28_0_io_out_a_0;
	wire [31:0] _mesh_28_0_io_out_c_0;
	wire [31:0] _mesh_28_0_io_out_b_0;
	wire _mesh_28_0_io_out_control_0_dataflow;
	wire _mesh_28_0_io_out_control_0_propagate;
	wire [4:0] _mesh_28_0_io_out_control_0_shift;
	wire [2:0] _mesh_28_0_io_out_id_0;
	wire _mesh_28_0_io_out_last_0;
	wire _mesh_28_0_io_out_valid_0;
	wire [31:0] _mesh_27_31_io_out_a_0;
	wire [31:0] _mesh_27_31_io_out_c_0;
	wire [31:0] _mesh_27_31_io_out_b_0;
	wire _mesh_27_31_io_out_control_0_dataflow;
	wire _mesh_27_31_io_out_control_0_propagate;
	wire [4:0] _mesh_27_31_io_out_control_0_shift;
	wire [2:0] _mesh_27_31_io_out_id_0;
	wire _mesh_27_31_io_out_last_0;
	wire _mesh_27_31_io_out_valid_0;
	wire [31:0] _mesh_27_30_io_out_a_0;
	wire [31:0] _mesh_27_30_io_out_c_0;
	wire [31:0] _mesh_27_30_io_out_b_0;
	wire _mesh_27_30_io_out_control_0_dataflow;
	wire _mesh_27_30_io_out_control_0_propagate;
	wire [4:0] _mesh_27_30_io_out_control_0_shift;
	wire [2:0] _mesh_27_30_io_out_id_0;
	wire _mesh_27_30_io_out_last_0;
	wire _mesh_27_30_io_out_valid_0;
	wire [31:0] _mesh_27_29_io_out_a_0;
	wire [31:0] _mesh_27_29_io_out_c_0;
	wire [31:0] _mesh_27_29_io_out_b_0;
	wire _mesh_27_29_io_out_control_0_dataflow;
	wire _mesh_27_29_io_out_control_0_propagate;
	wire [4:0] _mesh_27_29_io_out_control_0_shift;
	wire [2:0] _mesh_27_29_io_out_id_0;
	wire _mesh_27_29_io_out_last_0;
	wire _mesh_27_29_io_out_valid_0;
	wire [31:0] _mesh_27_28_io_out_a_0;
	wire [31:0] _mesh_27_28_io_out_c_0;
	wire [31:0] _mesh_27_28_io_out_b_0;
	wire _mesh_27_28_io_out_control_0_dataflow;
	wire _mesh_27_28_io_out_control_0_propagate;
	wire [4:0] _mesh_27_28_io_out_control_0_shift;
	wire [2:0] _mesh_27_28_io_out_id_0;
	wire _mesh_27_28_io_out_last_0;
	wire _mesh_27_28_io_out_valid_0;
	wire [31:0] _mesh_27_27_io_out_a_0;
	wire [31:0] _mesh_27_27_io_out_c_0;
	wire [31:0] _mesh_27_27_io_out_b_0;
	wire _mesh_27_27_io_out_control_0_dataflow;
	wire _mesh_27_27_io_out_control_0_propagate;
	wire [4:0] _mesh_27_27_io_out_control_0_shift;
	wire [2:0] _mesh_27_27_io_out_id_0;
	wire _mesh_27_27_io_out_last_0;
	wire _mesh_27_27_io_out_valid_0;
	wire [31:0] _mesh_27_26_io_out_a_0;
	wire [31:0] _mesh_27_26_io_out_c_0;
	wire [31:0] _mesh_27_26_io_out_b_0;
	wire _mesh_27_26_io_out_control_0_dataflow;
	wire _mesh_27_26_io_out_control_0_propagate;
	wire [4:0] _mesh_27_26_io_out_control_0_shift;
	wire [2:0] _mesh_27_26_io_out_id_0;
	wire _mesh_27_26_io_out_last_0;
	wire _mesh_27_26_io_out_valid_0;
	wire [31:0] _mesh_27_25_io_out_a_0;
	wire [31:0] _mesh_27_25_io_out_c_0;
	wire [31:0] _mesh_27_25_io_out_b_0;
	wire _mesh_27_25_io_out_control_0_dataflow;
	wire _mesh_27_25_io_out_control_0_propagate;
	wire [4:0] _mesh_27_25_io_out_control_0_shift;
	wire [2:0] _mesh_27_25_io_out_id_0;
	wire _mesh_27_25_io_out_last_0;
	wire _mesh_27_25_io_out_valid_0;
	wire [31:0] _mesh_27_24_io_out_a_0;
	wire [31:0] _mesh_27_24_io_out_c_0;
	wire [31:0] _mesh_27_24_io_out_b_0;
	wire _mesh_27_24_io_out_control_0_dataflow;
	wire _mesh_27_24_io_out_control_0_propagate;
	wire [4:0] _mesh_27_24_io_out_control_0_shift;
	wire [2:0] _mesh_27_24_io_out_id_0;
	wire _mesh_27_24_io_out_last_0;
	wire _mesh_27_24_io_out_valid_0;
	wire [31:0] _mesh_27_23_io_out_a_0;
	wire [31:0] _mesh_27_23_io_out_c_0;
	wire [31:0] _mesh_27_23_io_out_b_0;
	wire _mesh_27_23_io_out_control_0_dataflow;
	wire _mesh_27_23_io_out_control_0_propagate;
	wire [4:0] _mesh_27_23_io_out_control_0_shift;
	wire [2:0] _mesh_27_23_io_out_id_0;
	wire _mesh_27_23_io_out_last_0;
	wire _mesh_27_23_io_out_valid_0;
	wire [31:0] _mesh_27_22_io_out_a_0;
	wire [31:0] _mesh_27_22_io_out_c_0;
	wire [31:0] _mesh_27_22_io_out_b_0;
	wire _mesh_27_22_io_out_control_0_dataflow;
	wire _mesh_27_22_io_out_control_0_propagate;
	wire [4:0] _mesh_27_22_io_out_control_0_shift;
	wire [2:0] _mesh_27_22_io_out_id_0;
	wire _mesh_27_22_io_out_last_0;
	wire _mesh_27_22_io_out_valid_0;
	wire [31:0] _mesh_27_21_io_out_a_0;
	wire [31:0] _mesh_27_21_io_out_c_0;
	wire [31:0] _mesh_27_21_io_out_b_0;
	wire _mesh_27_21_io_out_control_0_dataflow;
	wire _mesh_27_21_io_out_control_0_propagate;
	wire [4:0] _mesh_27_21_io_out_control_0_shift;
	wire [2:0] _mesh_27_21_io_out_id_0;
	wire _mesh_27_21_io_out_last_0;
	wire _mesh_27_21_io_out_valid_0;
	wire [31:0] _mesh_27_20_io_out_a_0;
	wire [31:0] _mesh_27_20_io_out_c_0;
	wire [31:0] _mesh_27_20_io_out_b_0;
	wire _mesh_27_20_io_out_control_0_dataflow;
	wire _mesh_27_20_io_out_control_0_propagate;
	wire [4:0] _mesh_27_20_io_out_control_0_shift;
	wire [2:0] _mesh_27_20_io_out_id_0;
	wire _mesh_27_20_io_out_last_0;
	wire _mesh_27_20_io_out_valid_0;
	wire [31:0] _mesh_27_19_io_out_a_0;
	wire [31:0] _mesh_27_19_io_out_c_0;
	wire [31:0] _mesh_27_19_io_out_b_0;
	wire _mesh_27_19_io_out_control_0_dataflow;
	wire _mesh_27_19_io_out_control_0_propagate;
	wire [4:0] _mesh_27_19_io_out_control_0_shift;
	wire [2:0] _mesh_27_19_io_out_id_0;
	wire _mesh_27_19_io_out_last_0;
	wire _mesh_27_19_io_out_valid_0;
	wire [31:0] _mesh_27_18_io_out_a_0;
	wire [31:0] _mesh_27_18_io_out_c_0;
	wire [31:0] _mesh_27_18_io_out_b_0;
	wire _mesh_27_18_io_out_control_0_dataflow;
	wire _mesh_27_18_io_out_control_0_propagate;
	wire [4:0] _mesh_27_18_io_out_control_0_shift;
	wire [2:0] _mesh_27_18_io_out_id_0;
	wire _mesh_27_18_io_out_last_0;
	wire _mesh_27_18_io_out_valid_0;
	wire [31:0] _mesh_27_17_io_out_a_0;
	wire [31:0] _mesh_27_17_io_out_c_0;
	wire [31:0] _mesh_27_17_io_out_b_0;
	wire _mesh_27_17_io_out_control_0_dataflow;
	wire _mesh_27_17_io_out_control_0_propagate;
	wire [4:0] _mesh_27_17_io_out_control_0_shift;
	wire [2:0] _mesh_27_17_io_out_id_0;
	wire _mesh_27_17_io_out_last_0;
	wire _mesh_27_17_io_out_valid_0;
	wire [31:0] _mesh_27_16_io_out_a_0;
	wire [31:0] _mesh_27_16_io_out_c_0;
	wire [31:0] _mesh_27_16_io_out_b_0;
	wire _mesh_27_16_io_out_control_0_dataflow;
	wire _mesh_27_16_io_out_control_0_propagate;
	wire [4:0] _mesh_27_16_io_out_control_0_shift;
	wire [2:0] _mesh_27_16_io_out_id_0;
	wire _mesh_27_16_io_out_last_0;
	wire _mesh_27_16_io_out_valid_0;
	wire [31:0] _mesh_27_15_io_out_a_0;
	wire [31:0] _mesh_27_15_io_out_c_0;
	wire [31:0] _mesh_27_15_io_out_b_0;
	wire _mesh_27_15_io_out_control_0_dataflow;
	wire _mesh_27_15_io_out_control_0_propagate;
	wire [4:0] _mesh_27_15_io_out_control_0_shift;
	wire [2:0] _mesh_27_15_io_out_id_0;
	wire _mesh_27_15_io_out_last_0;
	wire _mesh_27_15_io_out_valid_0;
	wire [31:0] _mesh_27_14_io_out_a_0;
	wire [31:0] _mesh_27_14_io_out_c_0;
	wire [31:0] _mesh_27_14_io_out_b_0;
	wire _mesh_27_14_io_out_control_0_dataflow;
	wire _mesh_27_14_io_out_control_0_propagate;
	wire [4:0] _mesh_27_14_io_out_control_0_shift;
	wire [2:0] _mesh_27_14_io_out_id_0;
	wire _mesh_27_14_io_out_last_0;
	wire _mesh_27_14_io_out_valid_0;
	wire [31:0] _mesh_27_13_io_out_a_0;
	wire [31:0] _mesh_27_13_io_out_c_0;
	wire [31:0] _mesh_27_13_io_out_b_0;
	wire _mesh_27_13_io_out_control_0_dataflow;
	wire _mesh_27_13_io_out_control_0_propagate;
	wire [4:0] _mesh_27_13_io_out_control_0_shift;
	wire [2:0] _mesh_27_13_io_out_id_0;
	wire _mesh_27_13_io_out_last_0;
	wire _mesh_27_13_io_out_valid_0;
	wire [31:0] _mesh_27_12_io_out_a_0;
	wire [31:0] _mesh_27_12_io_out_c_0;
	wire [31:0] _mesh_27_12_io_out_b_0;
	wire _mesh_27_12_io_out_control_0_dataflow;
	wire _mesh_27_12_io_out_control_0_propagate;
	wire [4:0] _mesh_27_12_io_out_control_0_shift;
	wire [2:0] _mesh_27_12_io_out_id_0;
	wire _mesh_27_12_io_out_last_0;
	wire _mesh_27_12_io_out_valid_0;
	wire [31:0] _mesh_27_11_io_out_a_0;
	wire [31:0] _mesh_27_11_io_out_c_0;
	wire [31:0] _mesh_27_11_io_out_b_0;
	wire _mesh_27_11_io_out_control_0_dataflow;
	wire _mesh_27_11_io_out_control_0_propagate;
	wire [4:0] _mesh_27_11_io_out_control_0_shift;
	wire [2:0] _mesh_27_11_io_out_id_0;
	wire _mesh_27_11_io_out_last_0;
	wire _mesh_27_11_io_out_valid_0;
	wire [31:0] _mesh_27_10_io_out_a_0;
	wire [31:0] _mesh_27_10_io_out_c_0;
	wire [31:0] _mesh_27_10_io_out_b_0;
	wire _mesh_27_10_io_out_control_0_dataflow;
	wire _mesh_27_10_io_out_control_0_propagate;
	wire [4:0] _mesh_27_10_io_out_control_0_shift;
	wire [2:0] _mesh_27_10_io_out_id_0;
	wire _mesh_27_10_io_out_last_0;
	wire _mesh_27_10_io_out_valid_0;
	wire [31:0] _mesh_27_9_io_out_a_0;
	wire [31:0] _mesh_27_9_io_out_c_0;
	wire [31:0] _mesh_27_9_io_out_b_0;
	wire _mesh_27_9_io_out_control_0_dataflow;
	wire _mesh_27_9_io_out_control_0_propagate;
	wire [4:0] _mesh_27_9_io_out_control_0_shift;
	wire [2:0] _mesh_27_9_io_out_id_0;
	wire _mesh_27_9_io_out_last_0;
	wire _mesh_27_9_io_out_valid_0;
	wire [31:0] _mesh_27_8_io_out_a_0;
	wire [31:0] _mesh_27_8_io_out_c_0;
	wire [31:0] _mesh_27_8_io_out_b_0;
	wire _mesh_27_8_io_out_control_0_dataflow;
	wire _mesh_27_8_io_out_control_0_propagate;
	wire [4:0] _mesh_27_8_io_out_control_0_shift;
	wire [2:0] _mesh_27_8_io_out_id_0;
	wire _mesh_27_8_io_out_last_0;
	wire _mesh_27_8_io_out_valid_0;
	wire [31:0] _mesh_27_7_io_out_a_0;
	wire [31:0] _mesh_27_7_io_out_c_0;
	wire [31:0] _mesh_27_7_io_out_b_0;
	wire _mesh_27_7_io_out_control_0_dataflow;
	wire _mesh_27_7_io_out_control_0_propagate;
	wire [4:0] _mesh_27_7_io_out_control_0_shift;
	wire [2:0] _mesh_27_7_io_out_id_0;
	wire _mesh_27_7_io_out_last_0;
	wire _mesh_27_7_io_out_valid_0;
	wire [31:0] _mesh_27_6_io_out_a_0;
	wire [31:0] _mesh_27_6_io_out_c_0;
	wire [31:0] _mesh_27_6_io_out_b_0;
	wire _mesh_27_6_io_out_control_0_dataflow;
	wire _mesh_27_6_io_out_control_0_propagate;
	wire [4:0] _mesh_27_6_io_out_control_0_shift;
	wire [2:0] _mesh_27_6_io_out_id_0;
	wire _mesh_27_6_io_out_last_0;
	wire _mesh_27_6_io_out_valid_0;
	wire [31:0] _mesh_27_5_io_out_a_0;
	wire [31:0] _mesh_27_5_io_out_c_0;
	wire [31:0] _mesh_27_5_io_out_b_0;
	wire _mesh_27_5_io_out_control_0_dataflow;
	wire _mesh_27_5_io_out_control_0_propagate;
	wire [4:0] _mesh_27_5_io_out_control_0_shift;
	wire [2:0] _mesh_27_5_io_out_id_0;
	wire _mesh_27_5_io_out_last_0;
	wire _mesh_27_5_io_out_valid_0;
	wire [31:0] _mesh_27_4_io_out_a_0;
	wire [31:0] _mesh_27_4_io_out_c_0;
	wire [31:0] _mesh_27_4_io_out_b_0;
	wire _mesh_27_4_io_out_control_0_dataflow;
	wire _mesh_27_4_io_out_control_0_propagate;
	wire [4:0] _mesh_27_4_io_out_control_0_shift;
	wire [2:0] _mesh_27_4_io_out_id_0;
	wire _mesh_27_4_io_out_last_0;
	wire _mesh_27_4_io_out_valid_0;
	wire [31:0] _mesh_27_3_io_out_a_0;
	wire [31:0] _mesh_27_3_io_out_c_0;
	wire [31:0] _mesh_27_3_io_out_b_0;
	wire _mesh_27_3_io_out_control_0_dataflow;
	wire _mesh_27_3_io_out_control_0_propagate;
	wire [4:0] _mesh_27_3_io_out_control_0_shift;
	wire [2:0] _mesh_27_3_io_out_id_0;
	wire _mesh_27_3_io_out_last_0;
	wire _mesh_27_3_io_out_valid_0;
	wire [31:0] _mesh_27_2_io_out_a_0;
	wire [31:0] _mesh_27_2_io_out_c_0;
	wire [31:0] _mesh_27_2_io_out_b_0;
	wire _mesh_27_2_io_out_control_0_dataflow;
	wire _mesh_27_2_io_out_control_0_propagate;
	wire [4:0] _mesh_27_2_io_out_control_0_shift;
	wire [2:0] _mesh_27_2_io_out_id_0;
	wire _mesh_27_2_io_out_last_0;
	wire _mesh_27_2_io_out_valid_0;
	wire [31:0] _mesh_27_1_io_out_a_0;
	wire [31:0] _mesh_27_1_io_out_c_0;
	wire [31:0] _mesh_27_1_io_out_b_0;
	wire _mesh_27_1_io_out_control_0_dataflow;
	wire _mesh_27_1_io_out_control_0_propagate;
	wire [4:0] _mesh_27_1_io_out_control_0_shift;
	wire [2:0] _mesh_27_1_io_out_id_0;
	wire _mesh_27_1_io_out_last_0;
	wire _mesh_27_1_io_out_valid_0;
	wire [31:0] _mesh_27_0_io_out_a_0;
	wire [31:0] _mesh_27_0_io_out_c_0;
	wire [31:0] _mesh_27_0_io_out_b_0;
	wire _mesh_27_0_io_out_control_0_dataflow;
	wire _mesh_27_0_io_out_control_0_propagate;
	wire [4:0] _mesh_27_0_io_out_control_0_shift;
	wire [2:0] _mesh_27_0_io_out_id_0;
	wire _mesh_27_0_io_out_last_0;
	wire _mesh_27_0_io_out_valid_0;
	wire [31:0] _mesh_26_31_io_out_a_0;
	wire [31:0] _mesh_26_31_io_out_c_0;
	wire [31:0] _mesh_26_31_io_out_b_0;
	wire _mesh_26_31_io_out_control_0_dataflow;
	wire _mesh_26_31_io_out_control_0_propagate;
	wire [4:0] _mesh_26_31_io_out_control_0_shift;
	wire [2:0] _mesh_26_31_io_out_id_0;
	wire _mesh_26_31_io_out_last_0;
	wire _mesh_26_31_io_out_valid_0;
	wire [31:0] _mesh_26_30_io_out_a_0;
	wire [31:0] _mesh_26_30_io_out_c_0;
	wire [31:0] _mesh_26_30_io_out_b_0;
	wire _mesh_26_30_io_out_control_0_dataflow;
	wire _mesh_26_30_io_out_control_0_propagate;
	wire [4:0] _mesh_26_30_io_out_control_0_shift;
	wire [2:0] _mesh_26_30_io_out_id_0;
	wire _mesh_26_30_io_out_last_0;
	wire _mesh_26_30_io_out_valid_0;
	wire [31:0] _mesh_26_29_io_out_a_0;
	wire [31:0] _mesh_26_29_io_out_c_0;
	wire [31:0] _mesh_26_29_io_out_b_0;
	wire _mesh_26_29_io_out_control_0_dataflow;
	wire _mesh_26_29_io_out_control_0_propagate;
	wire [4:0] _mesh_26_29_io_out_control_0_shift;
	wire [2:0] _mesh_26_29_io_out_id_0;
	wire _mesh_26_29_io_out_last_0;
	wire _mesh_26_29_io_out_valid_0;
	wire [31:0] _mesh_26_28_io_out_a_0;
	wire [31:0] _mesh_26_28_io_out_c_0;
	wire [31:0] _mesh_26_28_io_out_b_0;
	wire _mesh_26_28_io_out_control_0_dataflow;
	wire _mesh_26_28_io_out_control_0_propagate;
	wire [4:0] _mesh_26_28_io_out_control_0_shift;
	wire [2:0] _mesh_26_28_io_out_id_0;
	wire _mesh_26_28_io_out_last_0;
	wire _mesh_26_28_io_out_valid_0;
	wire [31:0] _mesh_26_27_io_out_a_0;
	wire [31:0] _mesh_26_27_io_out_c_0;
	wire [31:0] _mesh_26_27_io_out_b_0;
	wire _mesh_26_27_io_out_control_0_dataflow;
	wire _mesh_26_27_io_out_control_0_propagate;
	wire [4:0] _mesh_26_27_io_out_control_0_shift;
	wire [2:0] _mesh_26_27_io_out_id_0;
	wire _mesh_26_27_io_out_last_0;
	wire _mesh_26_27_io_out_valid_0;
	wire [31:0] _mesh_26_26_io_out_a_0;
	wire [31:0] _mesh_26_26_io_out_c_0;
	wire [31:0] _mesh_26_26_io_out_b_0;
	wire _mesh_26_26_io_out_control_0_dataflow;
	wire _mesh_26_26_io_out_control_0_propagate;
	wire [4:0] _mesh_26_26_io_out_control_0_shift;
	wire [2:0] _mesh_26_26_io_out_id_0;
	wire _mesh_26_26_io_out_last_0;
	wire _mesh_26_26_io_out_valid_0;
	wire [31:0] _mesh_26_25_io_out_a_0;
	wire [31:0] _mesh_26_25_io_out_c_0;
	wire [31:0] _mesh_26_25_io_out_b_0;
	wire _mesh_26_25_io_out_control_0_dataflow;
	wire _mesh_26_25_io_out_control_0_propagate;
	wire [4:0] _mesh_26_25_io_out_control_0_shift;
	wire [2:0] _mesh_26_25_io_out_id_0;
	wire _mesh_26_25_io_out_last_0;
	wire _mesh_26_25_io_out_valid_0;
	wire [31:0] _mesh_26_24_io_out_a_0;
	wire [31:0] _mesh_26_24_io_out_c_0;
	wire [31:0] _mesh_26_24_io_out_b_0;
	wire _mesh_26_24_io_out_control_0_dataflow;
	wire _mesh_26_24_io_out_control_0_propagate;
	wire [4:0] _mesh_26_24_io_out_control_0_shift;
	wire [2:0] _mesh_26_24_io_out_id_0;
	wire _mesh_26_24_io_out_last_0;
	wire _mesh_26_24_io_out_valid_0;
	wire [31:0] _mesh_26_23_io_out_a_0;
	wire [31:0] _mesh_26_23_io_out_c_0;
	wire [31:0] _mesh_26_23_io_out_b_0;
	wire _mesh_26_23_io_out_control_0_dataflow;
	wire _mesh_26_23_io_out_control_0_propagate;
	wire [4:0] _mesh_26_23_io_out_control_0_shift;
	wire [2:0] _mesh_26_23_io_out_id_0;
	wire _mesh_26_23_io_out_last_0;
	wire _mesh_26_23_io_out_valid_0;
	wire [31:0] _mesh_26_22_io_out_a_0;
	wire [31:0] _mesh_26_22_io_out_c_0;
	wire [31:0] _mesh_26_22_io_out_b_0;
	wire _mesh_26_22_io_out_control_0_dataflow;
	wire _mesh_26_22_io_out_control_0_propagate;
	wire [4:0] _mesh_26_22_io_out_control_0_shift;
	wire [2:0] _mesh_26_22_io_out_id_0;
	wire _mesh_26_22_io_out_last_0;
	wire _mesh_26_22_io_out_valid_0;
	wire [31:0] _mesh_26_21_io_out_a_0;
	wire [31:0] _mesh_26_21_io_out_c_0;
	wire [31:0] _mesh_26_21_io_out_b_0;
	wire _mesh_26_21_io_out_control_0_dataflow;
	wire _mesh_26_21_io_out_control_0_propagate;
	wire [4:0] _mesh_26_21_io_out_control_0_shift;
	wire [2:0] _mesh_26_21_io_out_id_0;
	wire _mesh_26_21_io_out_last_0;
	wire _mesh_26_21_io_out_valid_0;
	wire [31:0] _mesh_26_20_io_out_a_0;
	wire [31:0] _mesh_26_20_io_out_c_0;
	wire [31:0] _mesh_26_20_io_out_b_0;
	wire _mesh_26_20_io_out_control_0_dataflow;
	wire _mesh_26_20_io_out_control_0_propagate;
	wire [4:0] _mesh_26_20_io_out_control_0_shift;
	wire [2:0] _mesh_26_20_io_out_id_0;
	wire _mesh_26_20_io_out_last_0;
	wire _mesh_26_20_io_out_valid_0;
	wire [31:0] _mesh_26_19_io_out_a_0;
	wire [31:0] _mesh_26_19_io_out_c_0;
	wire [31:0] _mesh_26_19_io_out_b_0;
	wire _mesh_26_19_io_out_control_0_dataflow;
	wire _mesh_26_19_io_out_control_0_propagate;
	wire [4:0] _mesh_26_19_io_out_control_0_shift;
	wire [2:0] _mesh_26_19_io_out_id_0;
	wire _mesh_26_19_io_out_last_0;
	wire _mesh_26_19_io_out_valid_0;
	wire [31:0] _mesh_26_18_io_out_a_0;
	wire [31:0] _mesh_26_18_io_out_c_0;
	wire [31:0] _mesh_26_18_io_out_b_0;
	wire _mesh_26_18_io_out_control_0_dataflow;
	wire _mesh_26_18_io_out_control_0_propagate;
	wire [4:0] _mesh_26_18_io_out_control_0_shift;
	wire [2:0] _mesh_26_18_io_out_id_0;
	wire _mesh_26_18_io_out_last_0;
	wire _mesh_26_18_io_out_valid_0;
	wire [31:0] _mesh_26_17_io_out_a_0;
	wire [31:0] _mesh_26_17_io_out_c_0;
	wire [31:0] _mesh_26_17_io_out_b_0;
	wire _mesh_26_17_io_out_control_0_dataflow;
	wire _mesh_26_17_io_out_control_0_propagate;
	wire [4:0] _mesh_26_17_io_out_control_0_shift;
	wire [2:0] _mesh_26_17_io_out_id_0;
	wire _mesh_26_17_io_out_last_0;
	wire _mesh_26_17_io_out_valid_0;
	wire [31:0] _mesh_26_16_io_out_a_0;
	wire [31:0] _mesh_26_16_io_out_c_0;
	wire [31:0] _mesh_26_16_io_out_b_0;
	wire _mesh_26_16_io_out_control_0_dataflow;
	wire _mesh_26_16_io_out_control_0_propagate;
	wire [4:0] _mesh_26_16_io_out_control_0_shift;
	wire [2:0] _mesh_26_16_io_out_id_0;
	wire _mesh_26_16_io_out_last_0;
	wire _mesh_26_16_io_out_valid_0;
	wire [31:0] _mesh_26_15_io_out_a_0;
	wire [31:0] _mesh_26_15_io_out_c_0;
	wire [31:0] _mesh_26_15_io_out_b_0;
	wire _mesh_26_15_io_out_control_0_dataflow;
	wire _mesh_26_15_io_out_control_0_propagate;
	wire [4:0] _mesh_26_15_io_out_control_0_shift;
	wire [2:0] _mesh_26_15_io_out_id_0;
	wire _mesh_26_15_io_out_last_0;
	wire _mesh_26_15_io_out_valid_0;
	wire [31:0] _mesh_26_14_io_out_a_0;
	wire [31:0] _mesh_26_14_io_out_c_0;
	wire [31:0] _mesh_26_14_io_out_b_0;
	wire _mesh_26_14_io_out_control_0_dataflow;
	wire _mesh_26_14_io_out_control_0_propagate;
	wire [4:0] _mesh_26_14_io_out_control_0_shift;
	wire [2:0] _mesh_26_14_io_out_id_0;
	wire _mesh_26_14_io_out_last_0;
	wire _mesh_26_14_io_out_valid_0;
	wire [31:0] _mesh_26_13_io_out_a_0;
	wire [31:0] _mesh_26_13_io_out_c_0;
	wire [31:0] _mesh_26_13_io_out_b_0;
	wire _mesh_26_13_io_out_control_0_dataflow;
	wire _mesh_26_13_io_out_control_0_propagate;
	wire [4:0] _mesh_26_13_io_out_control_0_shift;
	wire [2:0] _mesh_26_13_io_out_id_0;
	wire _mesh_26_13_io_out_last_0;
	wire _mesh_26_13_io_out_valid_0;
	wire [31:0] _mesh_26_12_io_out_a_0;
	wire [31:0] _mesh_26_12_io_out_c_0;
	wire [31:0] _mesh_26_12_io_out_b_0;
	wire _mesh_26_12_io_out_control_0_dataflow;
	wire _mesh_26_12_io_out_control_0_propagate;
	wire [4:0] _mesh_26_12_io_out_control_0_shift;
	wire [2:0] _mesh_26_12_io_out_id_0;
	wire _mesh_26_12_io_out_last_0;
	wire _mesh_26_12_io_out_valid_0;
	wire [31:0] _mesh_26_11_io_out_a_0;
	wire [31:0] _mesh_26_11_io_out_c_0;
	wire [31:0] _mesh_26_11_io_out_b_0;
	wire _mesh_26_11_io_out_control_0_dataflow;
	wire _mesh_26_11_io_out_control_0_propagate;
	wire [4:0] _mesh_26_11_io_out_control_0_shift;
	wire [2:0] _mesh_26_11_io_out_id_0;
	wire _mesh_26_11_io_out_last_0;
	wire _mesh_26_11_io_out_valid_0;
	wire [31:0] _mesh_26_10_io_out_a_0;
	wire [31:0] _mesh_26_10_io_out_c_0;
	wire [31:0] _mesh_26_10_io_out_b_0;
	wire _mesh_26_10_io_out_control_0_dataflow;
	wire _mesh_26_10_io_out_control_0_propagate;
	wire [4:0] _mesh_26_10_io_out_control_0_shift;
	wire [2:0] _mesh_26_10_io_out_id_0;
	wire _mesh_26_10_io_out_last_0;
	wire _mesh_26_10_io_out_valid_0;
	wire [31:0] _mesh_26_9_io_out_a_0;
	wire [31:0] _mesh_26_9_io_out_c_0;
	wire [31:0] _mesh_26_9_io_out_b_0;
	wire _mesh_26_9_io_out_control_0_dataflow;
	wire _mesh_26_9_io_out_control_0_propagate;
	wire [4:0] _mesh_26_9_io_out_control_0_shift;
	wire [2:0] _mesh_26_9_io_out_id_0;
	wire _mesh_26_9_io_out_last_0;
	wire _mesh_26_9_io_out_valid_0;
	wire [31:0] _mesh_26_8_io_out_a_0;
	wire [31:0] _mesh_26_8_io_out_c_0;
	wire [31:0] _mesh_26_8_io_out_b_0;
	wire _mesh_26_8_io_out_control_0_dataflow;
	wire _mesh_26_8_io_out_control_0_propagate;
	wire [4:0] _mesh_26_8_io_out_control_0_shift;
	wire [2:0] _mesh_26_8_io_out_id_0;
	wire _mesh_26_8_io_out_last_0;
	wire _mesh_26_8_io_out_valid_0;
	wire [31:0] _mesh_26_7_io_out_a_0;
	wire [31:0] _mesh_26_7_io_out_c_0;
	wire [31:0] _mesh_26_7_io_out_b_0;
	wire _mesh_26_7_io_out_control_0_dataflow;
	wire _mesh_26_7_io_out_control_0_propagate;
	wire [4:0] _mesh_26_7_io_out_control_0_shift;
	wire [2:0] _mesh_26_7_io_out_id_0;
	wire _mesh_26_7_io_out_last_0;
	wire _mesh_26_7_io_out_valid_0;
	wire [31:0] _mesh_26_6_io_out_a_0;
	wire [31:0] _mesh_26_6_io_out_c_0;
	wire [31:0] _mesh_26_6_io_out_b_0;
	wire _mesh_26_6_io_out_control_0_dataflow;
	wire _mesh_26_6_io_out_control_0_propagate;
	wire [4:0] _mesh_26_6_io_out_control_0_shift;
	wire [2:0] _mesh_26_6_io_out_id_0;
	wire _mesh_26_6_io_out_last_0;
	wire _mesh_26_6_io_out_valid_0;
	wire [31:0] _mesh_26_5_io_out_a_0;
	wire [31:0] _mesh_26_5_io_out_c_0;
	wire [31:0] _mesh_26_5_io_out_b_0;
	wire _mesh_26_5_io_out_control_0_dataflow;
	wire _mesh_26_5_io_out_control_0_propagate;
	wire [4:0] _mesh_26_5_io_out_control_0_shift;
	wire [2:0] _mesh_26_5_io_out_id_0;
	wire _mesh_26_5_io_out_last_0;
	wire _mesh_26_5_io_out_valid_0;
	wire [31:0] _mesh_26_4_io_out_a_0;
	wire [31:0] _mesh_26_4_io_out_c_0;
	wire [31:0] _mesh_26_4_io_out_b_0;
	wire _mesh_26_4_io_out_control_0_dataflow;
	wire _mesh_26_4_io_out_control_0_propagate;
	wire [4:0] _mesh_26_4_io_out_control_0_shift;
	wire [2:0] _mesh_26_4_io_out_id_0;
	wire _mesh_26_4_io_out_last_0;
	wire _mesh_26_4_io_out_valid_0;
	wire [31:0] _mesh_26_3_io_out_a_0;
	wire [31:0] _mesh_26_3_io_out_c_0;
	wire [31:0] _mesh_26_3_io_out_b_0;
	wire _mesh_26_3_io_out_control_0_dataflow;
	wire _mesh_26_3_io_out_control_0_propagate;
	wire [4:0] _mesh_26_3_io_out_control_0_shift;
	wire [2:0] _mesh_26_3_io_out_id_0;
	wire _mesh_26_3_io_out_last_0;
	wire _mesh_26_3_io_out_valid_0;
	wire [31:0] _mesh_26_2_io_out_a_0;
	wire [31:0] _mesh_26_2_io_out_c_0;
	wire [31:0] _mesh_26_2_io_out_b_0;
	wire _mesh_26_2_io_out_control_0_dataflow;
	wire _mesh_26_2_io_out_control_0_propagate;
	wire [4:0] _mesh_26_2_io_out_control_0_shift;
	wire [2:0] _mesh_26_2_io_out_id_0;
	wire _mesh_26_2_io_out_last_0;
	wire _mesh_26_2_io_out_valid_0;
	wire [31:0] _mesh_26_1_io_out_a_0;
	wire [31:0] _mesh_26_1_io_out_c_0;
	wire [31:0] _mesh_26_1_io_out_b_0;
	wire _mesh_26_1_io_out_control_0_dataflow;
	wire _mesh_26_1_io_out_control_0_propagate;
	wire [4:0] _mesh_26_1_io_out_control_0_shift;
	wire [2:0] _mesh_26_1_io_out_id_0;
	wire _mesh_26_1_io_out_last_0;
	wire _mesh_26_1_io_out_valid_0;
	wire [31:0] _mesh_26_0_io_out_a_0;
	wire [31:0] _mesh_26_0_io_out_c_0;
	wire [31:0] _mesh_26_0_io_out_b_0;
	wire _mesh_26_0_io_out_control_0_dataflow;
	wire _mesh_26_0_io_out_control_0_propagate;
	wire [4:0] _mesh_26_0_io_out_control_0_shift;
	wire [2:0] _mesh_26_0_io_out_id_0;
	wire _mesh_26_0_io_out_last_0;
	wire _mesh_26_0_io_out_valid_0;
	wire [31:0] _mesh_25_31_io_out_a_0;
	wire [31:0] _mesh_25_31_io_out_c_0;
	wire [31:0] _mesh_25_31_io_out_b_0;
	wire _mesh_25_31_io_out_control_0_dataflow;
	wire _mesh_25_31_io_out_control_0_propagate;
	wire [4:0] _mesh_25_31_io_out_control_0_shift;
	wire [2:0] _mesh_25_31_io_out_id_0;
	wire _mesh_25_31_io_out_last_0;
	wire _mesh_25_31_io_out_valid_0;
	wire [31:0] _mesh_25_30_io_out_a_0;
	wire [31:0] _mesh_25_30_io_out_c_0;
	wire [31:0] _mesh_25_30_io_out_b_0;
	wire _mesh_25_30_io_out_control_0_dataflow;
	wire _mesh_25_30_io_out_control_0_propagate;
	wire [4:0] _mesh_25_30_io_out_control_0_shift;
	wire [2:0] _mesh_25_30_io_out_id_0;
	wire _mesh_25_30_io_out_last_0;
	wire _mesh_25_30_io_out_valid_0;
	wire [31:0] _mesh_25_29_io_out_a_0;
	wire [31:0] _mesh_25_29_io_out_c_0;
	wire [31:0] _mesh_25_29_io_out_b_0;
	wire _mesh_25_29_io_out_control_0_dataflow;
	wire _mesh_25_29_io_out_control_0_propagate;
	wire [4:0] _mesh_25_29_io_out_control_0_shift;
	wire [2:0] _mesh_25_29_io_out_id_0;
	wire _mesh_25_29_io_out_last_0;
	wire _mesh_25_29_io_out_valid_0;
	wire [31:0] _mesh_25_28_io_out_a_0;
	wire [31:0] _mesh_25_28_io_out_c_0;
	wire [31:0] _mesh_25_28_io_out_b_0;
	wire _mesh_25_28_io_out_control_0_dataflow;
	wire _mesh_25_28_io_out_control_0_propagate;
	wire [4:0] _mesh_25_28_io_out_control_0_shift;
	wire [2:0] _mesh_25_28_io_out_id_0;
	wire _mesh_25_28_io_out_last_0;
	wire _mesh_25_28_io_out_valid_0;
	wire [31:0] _mesh_25_27_io_out_a_0;
	wire [31:0] _mesh_25_27_io_out_c_0;
	wire [31:0] _mesh_25_27_io_out_b_0;
	wire _mesh_25_27_io_out_control_0_dataflow;
	wire _mesh_25_27_io_out_control_0_propagate;
	wire [4:0] _mesh_25_27_io_out_control_0_shift;
	wire [2:0] _mesh_25_27_io_out_id_0;
	wire _mesh_25_27_io_out_last_0;
	wire _mesh_25_27_io_out_valid_0;
	wire [31:0] _mesh_25_26_io_out_a_0;
	wire [31:0] _mesh_25_26_io_out_c_0;
	wire [31:0] _mesh_25_26_io_out_b_0;
	wire _mesh_25_26_io_out_control_0_dataflow;
	wire _mesh_25_26_io_out_control_0_propagate;
	wire [4:0] _mesh_25_26_io_out_control_0_shift;
	wire [2:0] _mesh_25_26_io_out_id_0;
	wire _mesh_25_26_io_out_last_0;
	wire _mesh_25_26_io_out_valid_0;
	wire [31:0] _mesh_25_25_io_out_a_0;
	wire [31:0] _mesh_25_25_io_out_c_0;
	wire [31:0] _mesh_25_25_io_out_b_0;
	wire _mesh_25_25_io_out_control_0_dataflow;
	wire _mesh_25_25_io_out_control_0_propagate;
	wire [4:0] _mesh_25_25_io_out_control_0_shift;
	wire [2:0] _mesh_25_25_io_out_id_0;
	wire _mesh_25_25_io_out_last_0;
	wire _mesh_25_25_io_out_valid_0;
	wire [31:0] _mesh_25_24_io_out_a_0;
	wire [31:0] _mesh_25_24_io_out_c_0;
	wire [31:0] _mesh_25_24_io_out_b_0;
	wire _mesh_25_24_io_out_control_0_dataflow;
	wire _mesh_25_24_io_out_control_0_propagate;
	wire [4:0] _mesh_25_24_io_out_control_0_shift;
	wire [2:0] _mesh_25_24_io_out_id_0;
	wire _mesh_25_24_io_out_last_0;
	wire _mesh_25_24_io_out_valid_0;
	wire [31:0] _mesh_25_23_io_out_a_0;
	wire [31:0] _mesh_25_23_io_out_c_0;
	wire [31:0] _mesh_25_23_io_out_b_0;
	wire _mesh_25_23_io_out_control_0_dataflow;
	wire _mesh_25_23_io_out_control_0_propagate;
	wire [4:0] _mesh_25_23_io_out_control_0_shift;
	wire [2:0] _mesh_25_23_io_out_id_0;
	wire _mesh_25_23_io_out_last_0;
	wire _mesh_25_23_io_out_valid_0;
	wire [31:0] _mesh_25_22_io_out_a_0;
	wire [31:0] _mesh_25_22_io_out_c_0;
	wire [31:0] _mesh_25_22_io_out_b_0;
	wire _mesh_25_22_io_out_control_0_dataflow;
	wire _mesh_25_22_io_out_control_0_propagate;
	wire [4:0] _mesh_25_22_io_out_control_0_shift;
	wire [2:0] _mesh_25_22_io_out_id_0;
	wire _mesh_25_22_io_out_last_0;
	wire _mesh_25_22_io_out_valid_0;
	wire [31:0] _mesh_25_21_io_out_a_0;
	wire [31:0] _mesh_25_21_io_out_c_0;
	wire [31:0] _mesh_25_21_io_out_b_0;
	wire _mesh_25_21_io_out_control_0_dataflow;
	wire _mesh_25_21_io_out_control_0_propagate;
	wire [4:0] _mesh_25_21_io_out_control_0_shift;
	wire [2:0] _mesh_25_21_io_out_id_0;
	wire _mesh_25_21_io_out_last_0;
	wire _mesh_25_21_io_out_valid_0;
	wire [31:0] _mesh_25_20_io_out_a_0;
	wire [31:0] _mesh_25_20_io_out_c_0;
	wire [31:0] _mesh_25_20_io_out_b_0;
	wire _mesh_25_20_io_out_control_0_dataflow;
	wire _mesh_25_20_io_out_control_0_propagate;
	wire [4:0] _mesh_25_20_io_out_control_0_shift;
	wire [2:0] _mesh_25_20_io_out_id_0;
	wire _mesh_25_20_io_out_last_0;
	wire _mesh_25_20_io_out_valid_0;
	wire [31:0] _mesh_25_19_io_out_a_0;
	wire [31:0] _mesh_25_19_io_out_c_0;
	wire [31:0] _mesh_25_19_io_out_b_0;
	wire _mesh_25_19_io_out_control_0_dataflow;
	wire _mesh_25_19_io_out_control_0_propagate;
	wire [4:0] _mesh_25_19_io_out_control_0_shift;
	wire [2:0] _mesh_25_19_io_out_id_0;
	wire _mesh_25_19_io_out_last_0;
	wire _mesh_25_19_io_out_valid_0;
	wire [31:0] _mesh_25_18_io_out_a_0;
	wire [31:0] _mesh_25_18_io_out_c_0;
	wire [31:0] _mesh_25_18_io_out_b_0;
	wire _mesh_25_18_io_out_control_0_dataflow;
	wire _mesh_25_18_io_out_control_0_propagate;
	wire [4:0] _mesh_25_18_io_out_control_0_shift;
	wire [2:0] _mesh_25_18_io_out_id_0;
	wire _mesh_25_18_io_out_last_0;
	wire _mesh_25_18_io_out_valid_0;
	wire [31:0] _mesh_25_17_io_out_a_0;
	wire [31:0] _mesh_25_17_io_out_c_0;
	wire [31:0] _mesh_25_17_io_out_b_0;
	wire _mesh_25_17_io_out_control_0_dataflow;
	wire _mesh_25_17_io_out_control_0_propagate;
	wire [4:0] _mesh_25_17_io_out_control_0_shift;
	wire [2:0] _mesh_25_17_io_out_id_0;
	wire _mesh_25_17_io_out_last_0;
	wire _mesh_25_17_io_out_valid_0;
	wire [31:0] _mesh_25_16_io_out_a_0;
	wire [31:0] _mesh_25_16_io_out_c_0;
	wire [31:0] _mesh_25_16_io_out_b_0;
	wire _mesh_25_16_io_out_control_0_dataflow;
	wire _mesh_25_16_io_out_control_0_propagate;
	wire [4:0] _mesh_25_16_io_out_control_0_shift;
	wire [2:0] _mesh_25_16_io_out_id_0;
	wire _mesh_25_16_io_out_last_0;
	wire _mesh_25_16_io_out_valid_0;
	wire [31:0] _mesh_25_15_io_out_a_0;
	wire [31:0] _mesh_25_15_io_out_c_0;
	wire [31:0] _mesh_25_15_io_out_b_0;
	wire _mesh_25_15_io_out_control_0_dataflow;
	wire _mesh_25_15_io_out_control_0_propagate;
	wire [4:0] _mesh_25_15_io_out_control_0_shift;
	wire [2:0] _mesh_25_15_io_out_id_0;
	wire _mesh_25_15_io_out_last_0;
	wire _mesh_25_15_io_out_valid_0;
	wire [31:0] _mesh_25_14_io_out_a_0;
	wire [31:0] _mesh_25_14_io_out_c_0;
	wire [31:0] _mesh_25_14_io_out_b_0;
	wire _mesh_25_14_io_out_control_0_dataflow;
	wire _mesh_25_14_io_out_control_0_propagate;
	wire [4:0] _mesh_25_14_io_out_control_0_shift;
	wire [2:0] _mesh_25_14_io_out_id_0;
	wire _mesh_25_14_io_out_last_0;
	wire _mesh_25_14_io_out_valid_0;
	wire [31:0] _mesh_25_13_io_out_a_0;
	wire [31:0] _mesh_25_13_io_out_c_0;
	wire [31:0] _mesh_25_13_io_out_b_0;
	wire _mesh_25_13_io_out_control_0_dataflow;
	wire _mesh_25_13_io_out_control_0_propagate;
	wire [4:0] _mesh_25_13_io_out_control_0_shift;
	wire [2:0] _mesh_25_13_io_out_id_0;
	wire _mesh_25_13_io_out_last_0;
	wire _mesh_25_13_io_out_valid_0;
	wire [31:0] _mesh_25_12_io_out_a_0;
	wire [31:0] _mesh_25_12_io_out_c_0;
	wire [31:0] _mesh_25_12_io_out_b_0;
	wire _mesh_25_12_io_out_control_0_dataflow;
	wire _mesh_25_12_io_out_control_0_propagate;
	wire [4:0] _mesh_25_12_io_out_control_0_shift;
	wire [2:0] _mesh_25_12_io_out_id_0;
	wire _mesh_25_12_io_out_last_0;
	wire _mesh_25_12_io_out_valid_0;
	wire [31:0] _mesh_25_11_io_out_a_0;
	wire [31:0] _mesh_25_11_io_out_c_0;
	wire [31:0] _mesh_25_11_io_out_b_0;
	wire _mesh_25_11_io_out_control_0_dataflow;
	wire _mesh_25_11_io_out_control_0_propagate;
	wire [4:0] _mesh_25_11_io_out_control_0_shift;
	wire [2:0] _mesh_25_11_io_out_id_0;
	wire _mesh_25_11_io_out_last_0;
	wire _mesh_25_11_io_out_valid_0;
	wire [31:0] _mesh_25_10_io_out_a_0;
	wire [31:0] _mesh_25_10_io_out_c_0;
	wire [31:0] _mesh_25_10_io_out_b_0;
	wire _mesh_25_10_io_out_control_0_dataflow;
	wire _mesh_25_10_io_out_control_0_propagate;
	wire [4:0] _mesh_25_10_io_out_control_0_shift;
	wire [2:0] _mesh_25_10_io_out_id_0;
	wire _mesh_25_10_io_out_last_0;
	wire _mesh_25_10_io_out_valid_0;
	wire [31:0] _mesh_25_9_io_out_a_0;
	wire [31:0] _mesh_25_9_io_out_c_0;
	wire [31:0] _mesh_25_9_io_out_b_0;
	wire _mesh_25_9_io_out_control_0_dataflow;
	wire _mesh_25_9_io_out_control_0_propagate;
	wire [4:0] _mesh_25_9_io_out_control_0_shift;
	wire [2:0] _mesh_25_9_io_out_id_0;
	wire _mesh_25_9_io_out_last_0;
	wire _mesh_25_9_io_out_valid_0;
	wire [31:0] _mesh_25_8_io_out_a_0;
	wire [31:0] _mesh_25_8_io_out_c_0;
	wire [31:0] _mesh_25_8_io_out_b_0;
	wire _mesh_25_8_io_out_control_0_dataflow;
	wire _mesh_25_8_io_out_control_0_propagate;
	wire [4:0] _mesh_25_8_io_out_control_0_shift;
	wire [2:0] _mesh_25_8_io_out_id_0;
	wire _mesh_25_8_io_out_last_0;
	wire _mesh_25_8_io_out_valid_0;
	wire [31:0] _mesh_25_7_io_out_a_0;
	wire [31:0] _mesh_25_7_io_out_c_0;
	wire [31:0] _mesh_25_7_io_out_b_0;
	wire _mesh_25_7_io_out_control_0_dataflow;
	wire _mesh_25_7_io_out_control_0_propagate;
	wire [4:0] _mesh_25_7_io_out_control_0_shift;
	wire [2:0] _mesh_25_7_io_out_id_0;
	wire _mesh_25_7_io_out_last_0;
	wire _mesh_25_7_io_out_valid_0;
	wire [31:0] _mesh_25_6_io_out_a_0;
	wire [31:0] _mesh_25_6_io_out_c_0;
	wire [31:0] _mesh_25_6_io_out_b_0;
	wire _mesh_25_6_io_out_control_0_dataflow;
	wire _mesh_25_6_io_out_control_0_propagate;
	wire [4:0] _mesh_25_6_io_out_control_0_shift;
	wire [2:0] _mesh_25_6_io_out_id_0;
	wire _mesh_25_6_io_out_last_0;
	wire _mesh_25_6_io_out_valid_0;
	wire [31:0] _mesh_25_5_io_out_a_0;
	wire [31:0] _mesh_25_5_io_out_c_0;
	wire [31:0] _mesh_25_5_io_out_b_0;
	wire _mesh_25_5_io_out_control_0_dataflow;
	wire _mesh_25_5_io_out_control_0_propagate;
	wire [4:0] _mesh_25_5_io_out_control_0_shift;
	wire [2:0] _mesh_25_5_io_out_id_0;
	wire _mesh_25_5_io_out_last_0;
	wire _mesh_25_5_io_out_valid_0;
	wire [31:0] _mesh_25_4_io_out_a_0;
	wire [31:0] _mesh_25_4_io_out_c_0;
	wire [31:0] _mesh_25_4_io_out_b_0;
	wire _mesh_25_4_io_out_control_0_dataflow;
	wire _mesh_25_4_io_out_control_0_propagate;
	wire [4:0] _mesh_25_4_io_out_control_0_shift;
	wire [2:0] _mesh_25_4_io_out_id_0;
	wire _mesh_25_4_io_out_last_0;
	wire _mesh_25_4_io_out_valid_0;
	wire [31:0] _mesh_25_3_io_out_a_0;
	wire [31:0] _mesh_25_3_io_out_c_0;
	wire [31:0] _mesh_25_3_io_out_b_0;
	wire _mesh_25_3_io_out_control_0_dataflow;
	wire _mesh_25_3_io_out_control_0_propagate;
	wire [4:0] _mesh_25_3_io_out_control_0_shift;
	wire [2:0] _mesh_25_3_io_out_id_0;
	wire _mesh_25_3_io_out_last_0;
	wire _mesh_25_3_io_out_valid_0;
	wire [31:0] _mesh_25_2_io_out_a_0;
	wire [31:0] _mesh_25_2_io_out_c_0;
	wire [31:0] _mesh_25_2_io_out_b_0;
	wire _mesh_25_2_io_out_control_0_dataflow;
	wire _mesh_25_2_io_out_control_0_propagate;
	wire [4:0] _mesh_25_2_io_out_control_0_shift;
	wire [2:0] _mesh_25_2_io_out_id_0;
	wire _mesh_25_2_io_out_last_0;
	wire _mesh_25_2_io_out_valid_0;
	wire [31:0] _mesh_25_1_io_out_a_0;
	wire [31:0] _mesh_25_1_io_out_c_0;
	wire [31:0] _mesh_25_1_io_out_b_0;
	wire _mesh_25_1_io_out_control_0_dataflow;
	wire _mesh_25_1_io_out_control_0_propagate;
	wire [4:0] _mesh_25_1_io_out_control_0_shift;
	wire [2:0] _mesh_25_1_io_out_id_0;
	wire _mesh_25_1_io_out_last_0;
	wire _mesh_25_1_io_out_valid_0;
	wire [31:0] _mesh_25_0_io_out_a_0;
	wire [31:0] _mesh_25_0_io_out_c_0;
	wire [31:0] _mesh_25_0_io_out_b_0;
	wire _mesh_25_0_io_out_control_0_dataflow;
	wire _mesh_25_0_io_out_control_0_propagate;
	wire [4:0] _mesh_25_0_io_out_control_0_shift;
	wire [2:0] _mesh_25_0_io_out_id_0;
	wire _mesh_25_0_io_out_last_0;
	wire _mesh_25_0_io_out_valid_0;
	wire [31:0] _mesh_24_31_io_out_a_0;
	wire [31:0] _mesh_24_31_io_out_c_0;
	wire [31:0] _mesh_24_31_io_out_b_0;
	wire _mesh_24_31_io_out_control_0_dataflow;
	wire _mesh_24_31_io_out_control_0_propagate;
	wire [4:0] _mesh_24_31_io_out_control_0_shift;
	wire [2:0] _mesh_24_31_io_out_id_0;
	wire _mesh_24_31_io_out_last_0;
	wire _mesh_24_31_io_out_valid_0;
	wire [31:0] _mesh_24_30_io_out_a_0;
	wire [31:0] _mesh_24_30_io_out_c_0;
	wire [31:0] _mesh_24_30_io_out_b_0;
	wire _mesh_24_30_io_out_control_0_dataflow;
	wire _mesh_24_30_io_out_control_0_propagate;
	wire [4:0] _mesh_24_30_io_out_control_0_shift;
	wire [2:0] _mesh_24_30_io_out_id_0;
	wire _mesh_24_30_io_out_last_0;
	wire _mesh_24_30_io_out_valid_0;
	wire [31:0] _mesh_24_29_io_out_a_0;
	wire [31:0] _mesh_24_29_io_out_c_0;
	wire [31:0] _mesh_24_29_io_out_b_0;
	wire _mesh_24_29_io_out_control_0_dataflow;
	wire _mesh_24_29_io_out_control_0_propagate;
	wire [4:0] _mesh_24_29_io_out_control_0_shift;
	wire [2:0] _mesh_24_29_io_out_id_0;
	wire _mesh_24_29_io_out_last_0;
	wire _mesh_24_29_io_out_valid_0;
	wire [31:0] _mesh_24_28_io_out_a_0;
	wire [31:0] _mesh_24_28_io_out_c_0;
	wire [31:0] _mesh_24_28_io_out_b_0;
	wire _mesh_24_28_io_out_control_0_dataflow;
	wire _mesh_24_28_io_out_control_0_propagate;
	wire [4:0] _mesh_24_28_io_out_control_0_shift;
	wire [2:0] _mesh_24_28_io_out_id_0;
	wire _mesh_24_28_io_out_last_0;
	wire _mesh_24_28_io_out_valid_0;
	wire [31:0] _mesh_24_27_io_out_a_0;
	wire [31:0] _mesh_24_27_io_out_c_0;
	wire [31:0] _mesh_24_27_io_out_b_0;
	wire _mesh_24_27_io_out_control_0_dataflow;
	wire _mesh_24_27_io_out_control_0_propagate;
	wire [4:0] _mesh_24_27_io_out_control_0_shift;
	wire [2:0] _mesh_24_27_io_out_id_0;
	wire _mesh_24_27_io_out_last_0;
	wire _mesh_24_27_io_out_valid_0;
	wire [31:0] _mesh_24_26_io_out_a_0;
	wire [31:0] _mesh_24_26_io_out_c_0;
	wire [31:0] _mesh_24_26_io_out_b_0;
	wire _mesh_24_26_io_out_control_0_dataflow;
	wire _mesh_24_26_io_out_control_0_propagate;
	wire [4:0] _mesh_24_26_io_out_control_0_shift;
	wire [2:0] _mesh_24_26_io_out_id_0;
	wire _mesh_24_26_io_out_last_0;
	wire _mesh_24_26_io_out_valid_0;
	wire [31:0] _mesh_24_25_io_out_a_0;
	wire [31:0] _mesh_24_25_io_out_c_0;
	wire [31:0] _mesh_24_25_io_out_b_0;
	wire _mesh_24_25_io_out_control_0_dataflow;
	wire _mesh_24_25_io_out_control_0_propagate;
	wire [4:0] _mesh_24_25_io_out_control_0_shift;
	wire [2:0] _mesh_24_25_io_out_id_0;
	wire _mesh_24_25_io_out_last_0;
	wire _mesh_24_25_io_out_valid_0;
	wire [31:0] _mesh_24_24_io_out_a_0;
	wire [31:0] _mesh_24_24_io_out_c_0;
	wire [31:0] _mesh_24_24_io_out_b_0;
	wire _mesh_24_24_io_out_control_0_dataflow;
	wire _mesh_24_24_io_out_control_0_propagate;
	wire [4:0] _mesh_24_24_io_out_control_0_shift;
	wire [2:0] _mesh_24_24_io_out_id_0;
	wire _mesh_24_24_io_out_last_0;
	wire _mesh_24_24_io_out_valid_0;
	wire [31:0] _mesh_24_23_io_out_a_0;
	wire [31:0] _mesh_24_23_io_out_c_0;
	wire [31:0] _mesh_24_23_io_out_b_0;
	wire _mesh_24_23_io_out_control_0_dataflow;
	wire _mesh_24_23_io_out_control_0_propagate;
	wire [4:0] _mesh_24_23_io_out_control_0_shift;
	wire [2:0] _mesh_24_23_io_out_id_0;
	wire _mesh_24_23_io_out_last_0;
	wire _mesh_24_23_io_out_valid_0;
	wire [31:0] _mesh_24_22_io_out_a_0;
	wire [31:0] _mesh_24_22_io_out_c_0;
	wire [31:0] _mesh_24_22_io_out_b_0;
	wire _mesh_24_22_io_out_control_0_dataflow;
	wire _mesh_24_22_io_out_control_0_propagate;
	wire [4:0] _mesh_24_22_io_out_control_0_shift;
	wire [2:0] _mesh_24_22_io_out_id_0;
	wire _mesh_24_22_io_out_last_0;
	wire _mesh_24_22_io_out_valid_0;
	wire [31:0] _mesh_24_21_io_out_a_0;
	wire [31:0] _mesh_24_21_io_out_c_0;
	wire [31:0] _mesh_24_21_io_out_b_0;
	wire _mesh_24_21_io_out_control_0_dataflow;
	wire _mesh_24_21_io_out_control_0_propagate;
	wire [4:0] _mesh_24_21_io_out_control_0_shift;
	wire [2:0] _mesh_24_21_io_out_id_0;
	wire _mesh_24_21_io_out_last_0;
	wire _mesh_24_21_io_out_valid_0;
	wire [31:0] _mesh_24_20_io_out_a_0;
	wire [31:0] _mesh_24_20_io_out_c_0;
	wire [31:0] _mesh_24_20_io_out_b_0;
	wire _mesh_24_20_io_out_control_0_dataflow;
	wire _mesh_24_20_io_out_control_0_propagate;
	wire [4:0] _mesh_24_20_io_out_control_0_shift;
	wire [2:0] _mesh_24_20_io_out_id_0;
	wire _mesh_24_20_io_out_last_0;
	wire _mesh_24_20_io_out_valid_0;
	wire [31:0] _mesh_24_19_io_out_a_0;
	wire [31:0] _mesh_24_19_io_out_c_0;
	wire [31:0] _mesh_24_19_io_out_b_0;
	wire _mesh_24_19_io_out_control_0_dataflow;
	wire _mesh_24_19_io_out_control_0_propagate;
	wire [4:0] _mesh_24_19_io_out_control_0_shift;
	wire [2:0] _mesh_24_19_io_out_id_0;
	wire _mesh_24_19_io_out_last_0;
	wire _mesh_24_19_io_out_valid_0;
	wire [31:0] _mesh_24_18_io_out_a_0;
	wire [31:0] _mesh_24_18_io_out_c_0;
	wire [31:0] _mesh_24_18_io_out_b_0;
	wire _mesh_24_18_io_out_control_0_dataflow;
	wire _mesh_24_18_io_out_control_0_propagate;
	wire [4:0] _mesh_24_18_io_out_control_0_shift;
	wire [2:0] _mesh_24_18_io_out_id_0;
	wire _mesh_24_18_io_out_last_0;
	wire _mesh_24_18_io_out_valid_0;
	wire [31:0] _mesh_24_17_io_out_a_0;
	wire [31:0] _mesh_24_17_io_out_c_0;
	wire [31:0] _mesh_24_17_io_out_b_0;
	wire _mesh_24_17_io_out_control_0_dataflow;
	wire _mesh_24_17_io_out_control_0_propagate;
	wire [4:0] _mesh_24_17_io_out_control_0_shift;
	wire [2:0] _mesh_24_17_io_out_id_0;
	wire _mesh_24_17_io_out_last_0;
	wire _mesh_24_17_io_out_valid_0;
	wire [31:0] _mesh_24_16_io_out_a_0;
	wire [31:0] _mesh_24_16_io_out_c_0;
	wire [31:0] _mesh_24_16_io_out_b_0;
	wire _mesh_24_16_io_out_control_0_dataflow;
	wire _mesh_24_16_io_out_control_0_propagate;
	wire [4:0] _mesh_24_16_io_out_control_0_shift;
	wire [2:0] _mesh_24_16_io_out_id_0;
	wire _mesh_24_16_io_out_last_0;
	wire _mesh_24_16_io_out_valid_0;
	wire [31:0] _mesh_24_15_io_out_a_0;
	wire [31:0] _mesh_24_15_io_out_c_0;
	wire [31:0] _mesh_24_15_io_out_b_0;
	wire _mesh_24_15_io_out_control_0_dataflow;
	wire _mesh_24_15_io_out_control_0_propagate;
	wire [4:0] _mesh_24_15_io_out_control_0_shift;
	wire [2:0] _mesh_24_15_io_out_id_0;
	wire _mesh_24_15_io_out_last_0;
	wire _mesh_24_15_io_out_valid_0;
	wire [31:0] _mesh_24_14_io_out_a_0;
	wire [31:0] _mesh_24_14_io_out_c_0;
	wire [31:0] _mesh_24_14_io_out_b_0;
	wire _mesh_24_14_io_out_control_0_dataflow;
	wire _mesh_24_14_io_out_control_0_propagate;
	wire [4:0] _mesh_24_14_io_out_control_0_shift;
	wire [2:0] _mesh_24_14_io_out_id_0;
	wire _mesh_24_14_io_out_last_0;
	wire _mesh_24_14_io_out_valid_0;
	wire [31:0] _mesh_24_13_io_out_a_0;
	wire [31:0] _mesh_24_13_io_out_c_0;
	wire [31:0] _mesh_24_13_io_out_b_0;
	wire _mesh_24_13_io_out_control_0_dataflow;
	wire _mesh_24_13_io_out_control_0_propagate;
	wire [4:0] _mesh_24_13_io_out_control_0_shift;
	wire [2:0] _mesh_24_13_io_out_id_0;
	wire _mesh_24_13_io_out_last_0;
	wire _mesh_24_13_io_out_valid_0;
	wire [31:0] _mesh_24_12_io_out_a_0;
	wire [31:0] _mesh_24_12_io_out_c_0;
	wire [31:0] _mesh_24_12_io_out_b_0;
	wire _mesh_24_12_io_out_control_0_dataflow;
	wire _mesh_24_12_io_out_control_0_propagate;
	wire [4:0] _mesh_24_12_io_out_control_0_shift;
	wire [2:0] _mesh_24_12_io_out_id_0;
	wire _mesh_24_12_io_out_last_0;
	wire _mesh_24_12_io_out_valid_0;
	wire [31:0] _mesh_24_11_io_out_a_0;
	wire [31:0] _mesh_24_11_io_out_c_0;
	wire [31:0] _mesh_24_11_io_out_b_0;
	wire _mesh_24_11_io_out_control_0_dataflow;
	wire _mesh_24_11_io_out_control_0_propagate;
	wire [4:0] _mesh_24_11_io_out_control_0_shift;
	wire [2:0] _mesh_24_11_io_out_id_0;
	wire _mesh_24_11_io_out_last_0;
	wire _mesh_24_11_io_out_valid_0;
	wire [31:0] _mesh_24_10_io_out_a_0;
	wire [31:0] _mesh_24_10_io_out_c_0;
	wire [31:0] _mesh_24_10_io_out_b_0;
	wire _mesh_24_10_io_out_control_0_dataflow;
	wire _mesh_24_10_io_out_control_0_propagate;
	wire [4:0] _mesh_24_10_io_out_control_0_shift;
	wire [2:0] _mesh_24_10_io_out_id_0;
	wire _mesh_24_10_io_out_last_0;
	wire _mesh_24_10_io_out_valid_0;
	wire [31:0] _mesh_24_9_io_out_a_0;
	wire [31:0] _mesh_24_9_io_out_c_0;
	wire [31:0] _mesh_24_9_io_out_b_0;
	wire _mesh_24_9_io_out_control_0_dataflow;
	wire _mesh_24_9_io_out_control_0_propagate;
	wire [4:0] _mesh_24_9_io_out_control_0_shift;
	wire [2:0] _mesh_24_9_io_out_id_0;
	wire _mesh_24_9_io_out_last_0;
	wire _mesh_24_9_io_out_valid_0;
	wire [31:0] _mesh_24_8_io_out_a_0;
	wire [31:0] _mesh_24_8_io_out_c_0;
	wire [31:0] _mesh_24_8_io_out_b_0;
	wire _mesh_24_8_io_out_control_0_dataflow;
	wire _mesh_24_8_io_out_control_0_propagate;
	wire [4:0] _mesh_24_8_io_out_control_0_shift;
	wire [2:0] _mesh_24_8_io_out_id_0;
	wire _mesh_24_8_io_out_last_0;
	wire _mesh_24_8_io_out_valid_0;
	wire [31:0] _mesh_24_7_io_out_a_0;
	wire [31:0] _mesh_24_7_io_out_c_0;
	wire [31:0] _mesh_24_7_io_out_b_0;
	wire _mesh_24_7_io_out_control_0_dataflow;
	wire _mesh_24_7_io_out_control_0_propagate;
	wire [4:0] _mesh_24_7_io_out_control_0_shift;
	wire [2:0] _mesh_24_7_io_out_id_0;
	wire _mesh_24_7_io_out_last_0;
	wire _mesh_24_7_io_out_valid_0;
	wire [31:0] _mesh_24_6_io_out_a_0;
	wire [31:0] _mesh_24_6_io_out_c_0;
	wire [31:0] _mesh_24_6_io_out_b_0;
	wire _mesh_24_6_io_out_control_0_dataflow;
	wire _mesh_24_6_io_out_control_0_propagate;
	wire [4:0] _mesh_24_6_io_out_control_0_shift;
	wire [2:0] _mesh_24_6_io_out_id_0;
	wire _mesh_24_6_io_out_last_0;
	wire _mesh_24_6_io_out_valid_0;
	wire [31:0] _mesh_24_5_io_out_a_0;
	wire [31:0] _mesh_24_5_io_out_c_0;
	wire [31:0] _mesh_24_5_io_out_b_0;
	wire _mesh_24_5_io_out_control_0_dataflow;
	wire _mesh_24_5_io_out_control_0_propagate;
	wire [4:0] _mesh_24_5_io_out_control_0_shift;
	wire [2:0] _mesh_24_5_io_out_id_0;
	wire _mesh_24_5_io_out_last_0;
	wire _mesh_24_5_io_out_valid_0;
	wire [31:0] _mesh_24_4_io_out_a_0;
	wire [31:0] _mesh_24_4_io_out_c_0;
	wire [31:0] _mesh_24_4_io_out_b_0;
	wire _mesh_24_4_io_out_control_0_dataflow;
	wire _mesh_24_4_io_out_control_0_propagate;
	wire [4:0] _mesh_24_4_io_out_control_0_shift;
	wire [2:0] _mesh_24_4_io_out_id_0;
	wire _mesh_24_4_io_out_last_0;
	wire _mesh_24_4_io_out_valid_0;
	wire [31:0] _mesh_24_3_io_out_a_0;
	wire [31:0] _mesh_24_3_io_out_c_0;
	wire [31:0] _mesh_24_3_io_out_b_0;
	wire _mesh_24_3_io_out_control_0_dataflow;
	wire _mesh_24_3_io_out_control_0_propagate;
	wire [4:0] _mesh_24_3_io_out_control_0_shift;
	wire [2:0] _mesh_24_3_io_out_id_0;
	wire _mesh_24_3_io_out_last_0;
	wire _mesh_24_3_io_out_valid_0;
	wire [31:0] _mesh_24_2_io_out_a_0;
	wire [31:0] _mesh_24_2_io_out_c_0;
	wire [31:0] _mesh_24_2_io_out_b_0;
	wire _mesh_24_2_io_out_control_0_dataflow;
	wire _mesh_24_2_io_out_control_0_propagate;
	wire [4:0] _mesh_24_2_io_out_control_0_shift;
	wire [2:0] _mesh_24_2_io_out_id_0;
	wire _mesh_24_2_io_out_last_0;
	wire _mesh_24_2_io_out_valid_0;
	wire [31:0] _mesh_24_1_io_out_a_0;
	wire [31:0] _mesh_24_1_io_out_c_0;
	wire [31:0] _mesh_24_1_io_out_b_0;
	wire _mesh_24_1_io_out_control_0_dataflow;
	wire _mesh_24_1_io_out_control_0_propagate;
	wire [4:0] _mesh_24_1_io_out_control_0_shift;
	wire [2:0] _mesh_24_1_io_out_id_0;
	wire _mesh_24_1_io_out_last_0;
	wire _mesh_24_1_io_out_valid_0;
	wire [31:0] _mesh_24_0_io_out_a_0;
	wire [31:0] _mesh_24_0_io_out_c_0;
	wire [31:0] _mesh_24_0_io_out_b_0;
	wire _mesh_24_0_io_out_control_0_dataflow;
	wire _mesh_24_0_io_out_control_0_propagate;
	wire [4:0] _mesh_24_0_io_out_control_0_shift;
	wire [2:0] _mesh_24_0_io_out_id_0;
	wire _mesh_24_0_io_out_last_0;
	wire _mesh_24_0_io_out_valid_0;
	wire [31:0] _mesh_23_31_io_out_a_0;
	wire [31:0] _mesh_23_31_io_out_c_0;
	wire [31:0] _mesh_23_31_io_out_b_0;
	wire _mesh_23_31_io_out_control_0_dataflow;
	wire _mesh_23_31_io_out_control_0_propagate;
	wire [4:0] _mesh_23_31_io_out_control_0_shift;
	wire [2:0] _mesh_23_31_io_out_id_0;
	wire _mesh_23_31_io_out_last_0;
	wire _mesh_23_31_io_out_valid_0;
	wire [31:0] _mesh_23_30_io_out_a_0;
	wire [31:0] _mesh_23_30_io_out_c_0;
	wire [31:0] _mesh_23_30_io_out_b_0;
	wire _mesh_23_30_io_out_control_0_dataflow;
	wire _mesh_23_30_io_out_control_0_propagate;
	wire [4:0] _mesh_23_30_io_out_control_0_shift;
	wire [2:0] _mesh_23_30_io_out_id_0;
	wire _mesh_23_30_io_out_last_0;
	wire _mesh_23_30_io_out_valid_0;
	wire [31:0] _mesh_23_29_io_out_a_0;
	wire [31:0] _mesh_23_29_io_out_c_0;
	wire [31:0] _mesh_23_29_io_out_b_0;
	wire _mesh_23_29_io_out_control_0_dataflow;
	wire _mesh_23_29_io_out_control_0_propagate;
	wire [4:0] _mesh_23_29_io_out_control_0_shift;
	wire [2:0] _mesh_23_29_io_out_id_0;
	wire _mesh_23_29_io_out_last_0;
	wire _mesh_23_29_io_out_valid_0;
	wire [31:0] _mesh_23_28_io_out_a_0;
	wire [31:0] _mesh_23_28_io_out_c_0;
	wire [31:0] _mesh_23_28_io_out_b_0;
	wire _mesh_23_28_io_out_control_0_dataflow;
	wire _mesh_23_28_io_out_control_0_propagate;
	wire [4:0] _mesh_23_28_io_out_control_0_shift;
	wire [2:0] _mesh_23_28_io_out_id_0;
	wire _mesh_23_28_io_out_last_0;
	wire _mesh_23_28_io_out_valid_0;
	wire [31:0] _mesh_23_27_io_out_a_0;
	wire [31:0] _mesh_23_27_io_out_c_0;
	wire [31:0] _mesh_23_27_io_out_b_0;
	wire _mesh_23_27_io_out_control_0_dataflow;
	wire _mesh_23_27_io_out_control_0_propagate;
	wire [4:0] _mesh_23_27_io_out_control_0_shift;
	wire [2:0] _mesh_23_27_io_out_id_0;
	wire _mesh_23_27_io_out_last_0;
	wire _mesh_23_27_io_out_valid_0;
	wire [31:0] _mesh_23_26_io_out_a_0;
	wire [31:0] _mesh_23_26_io_out_c_0;
	wire [31:0] _mesh_23_26_io_out_b_0;
	wire _mesh_23_26_io_out_control_0_dataflow;
	wire _mesh_23_26_io_out_control_0_propagate;
	wire [4:0] _mesh_23_26_io_out_control_0_shift;
	wire [2:0] _mesh_23_26_io_out_id_0;
	wire _mesh_23_26_io_out_last_0;
	wire _mesh_23_26_io_out_valid_0;
	wire [31:0] _mesh_23_25_io_out_a_0;
	wire [31:0] _mesh_23_25_io_out_c_0;
	wire [31:0] _mesh_23_25_io_out_b_0;
	wire _mesh_23_25_io_out_control_0_dataflow;
	wire _mesh_23_25_io_out_control_0_propagate;
	wire [4:0] _mesh_23_25_io_out_control_0_shift;
	wire [2:0] _mesh_23_25_io_out_id_0;
	wire _mesh_23_25_io_out_last_0;
	wire _mesh_23_25_io_out_valid_0;
	wire [31:0] _mesh_23_24_io_out_a_0;
	wire [31:0] _mesh_23_24_io_out_c_0;
	wire [31:0] _mesh_23_24_io_out_b_0;
	wire _mesh_23_24_io_out_control_0_dataflow;
	wire _mesh_23_24_io_out_control_0_propagate;
	wire [4:0] _mesh_23_24_io_out_control_0_shift;
	wire [2:0] _mesh_23_24_io_out_id_0;
	wire _mesh_23_24_io_out_last_0;
	wire _mesh_23_24_io_out_valid_0;
	wire [31:0] _mesh_23_23_io_out_a_0;
	wire [31:0] _mesh_23_23_io_out_c_0;
	wire [31:0] _mesh_23_23_io_out_b_0;
	wire _mesh_23_23_io_out_control_0_dataflow;
	wire _mesh_23_23_io_out_control_0_propagate;
	wire [4:0] _mesh_23_23_io_out_control_0_shift;
	wire [2:0] _mesh_23_23_io_out_id_0;
	wire _mesh_23_23_io_out_last_0;
	wire _mesh_23_23_io_out_valid_0;
	wire [31:0] _mesh_23_22_io_out_a_0;
	wire [31:0] _mesh_23_22_io_out_c_0;
	wire [31:0] _mesh_23_22_io_out_b_0;
	wire _mesh_23_22_io_out_control_0_dataflow;
	wire _mesh_23_22_io_out_control_0_propagate;
	wire [4:0] _mesh_23_22_io_out_control_0_shift;
	wire [2:0] _mesh_23_22_io_out_id_0;
	wire _mesh_23_22_io_out_last_0;
	wire _mesh_23_22_io_out_valid_0;
	wire [31:0] _mesh_23_21_io_out_a_0;
	wire [31:0] _mesh_23_21_io_out_c_0;
	wire [31:0] _mesh_23_21_io_out_b_0;
	wire _mesh_23_21_io_out_control_0_dataflow;
	wire _mesh_23_21_io_out_control_0_propagate;
	wire [4:0] _mesh_23_21_io_out_control_0_shift;
	wire [2:0] _mesh_23_21_io_out_id_0;
	wire _mesh_23_21_io_out_last_0;
	wire _mesh_23_21_io_out_valid_0;
	wire [31:0] _mesh_23_20_io_out_a_0;
	wire [31:0] _mesh_23_20_io_out_c_0;
	wire [31:0] _mesh_23_20_io_out_b_0;
	wire _mesh_23_20_io_out_control_0_dataflow;
	wire _mesh_23_20_io_out_control_0_propagate;
	wire [4:0] _mesh_23_20_io_out_control_0_shift;
	wire [2:0] _mesh_23_20_io_out_id_0;
	wire _mesh_23_20_io_out_last_0;
	wire _mesh_23_20_io_out_valid_0;
	wire [31:0] _mesh_23_19_io_out_a_0;
	wire [31:0] _mesh_23_19_io_out_c_0;
	wire [31:0] _mesh_23_19_io_out_b_0;
	wire _mesh_23_19_io_out_control_0_dataflow;
	wire _mesh_23_19_io_out_control_0_propagate;
	wire [4:0] _mesh_23_19_io_out_control_0_shift;
	wire [2:0] _mesh_23_19_io_out_id_0;
	wire _mesh_23_19_io_out_last_0;
	wire _mesh_23_19_io_out_valid_0;
	wire [31:0] _mesh_23_18_io_out_a_0;
	wire [31:0] _mesh_23_18_io_out_c_0;
	wire [31:0] _mesh_23_18_io_out_b_0;
	wire _mesh_23_18_io_out_control_0_dataflow;
	wire _mesh_23_18_io_out_control_0_propagate;
	wire [4:0] _mesh_23_18_io_out_control_0_shift;
	wire [2:0] _mesh_23_18_io_out_id_0;
	wire _mesh_23_18_io_out_last_0;
	wire _mesh_23_18_io_out_valid_0;
	wire [31:0] _mesh_23_17_io_out_a_0;
	wire [31:0] _mesh_23_17_io_out_c_0;
	wire [31:0] _mesh_23_17_io_out_b_0;
	wire _mesh_23_17_io_out_control_0_dataflow;
	wire _mesh_23_17_io_out_control_0_propagate;
	wire [4:0] _mesh_23_17_io_out_control_0_shift;
	wire [2:0] _mesh_23_17_io_out_id_0;
	wire _mesh_23_17_io_out_last_0;
	wire _mesh_23_17_io_out_valid_0;
	wire [31:0] _mesh_23_16_io_out_a_0;
	wire [31:0] _mesh_23_16_io_out_c_0;
	wire [31:0] _mesh_23_16_io_out_b_0;
	wire _mesh_23_16_io_out_control_0_dataflow;
	wire _mesh_23_16_io_out_control_0_propagate;
	wire [4:0] _mesh_23_16_io_out_control_0_shift;
	wire [2:0] _mesh_23_16_io_out_id_0;
	wire _mesh_23_16_io_out_last_0;
	wire _mesh_23_16_io_out_valid_0;
	wire [31:0] _mesh_23_15_io_out_a_0;
	wire [31:0] _mesh_23_15_io_out_c_0;
	wire [31:0] _mesh_23_15_io_out_b_0;
	wire _mesh_23_15_io_out_control_0_dataflow;
	wire _mesh_23_15_io_out_control_0_propagate;
	wire [4:0] _mesh_23_15_io_out_control_0_shift;
	wire [2:0] _mesh_23_15_io_out_id_0;
	wire _mesh_23_15_io_out_last_0;
	wire _mesh_23_15_io_out_valid_0;
	wire [31:0] _mesh_23_14_io_out_a_0;
	wire [31:0] _mesh_23_14_io_out_c_0;
	wire [31:0] _mesh_23_14_io_out_b_0;
	wire _mesh_23_14_io_out_control_0_dataflow;
	wire _mesh_23_14_io_out_control_0_propagate;
	wire [4:0] _mesh_23_14_io_out_control_0_shift;
	wire [2:0] _mesh_23_14_io_out_id_0;
	wire _mesh_23_14_io_out_last_0;
	wire _mesh_23_14_io_out_valid_0;
	wire [31:0] _mesh_23_13_io_out_a_0;
	wire [31:0] _mesh_23_13_io_out_c_0;
	wire [31:0] _mesh_23_13_io_out_b_0;
	wire _mesh_23_13_io_out_control_0_dataflow;
	wire _mesh_23_13_io_out_control_0_propagate;
	wire [4:0] _mesh_23_13_io_out_control_0_shift;
	wire [2:0] _mesh_23_13_io_out_id_0;
	wire _mesh_23_13_io_out_last_0;
	wire _mesh_23_13_io_out_valid_0;
	wire [31:0] _mesh_23_12_io_out_a_0;
	wire [31:0] _mesh_23_12_io_out_c_0;
	wire [31:0] _mesh_23_12_io_out_b_0;
	wire _mesh_23_12_io_out_control_0_dataflow;
	wire _mesh_23_12_io_out_control_0_propagate;
	wire [4:0] _mesh_23_12_io_out_control_0_shift;
	wire [2:0] _mesh_23_12_io_out_id_0;
	wire _mesh_23_12_io_out_last_0;
	wire _mesh_23_12_io_out_valid_0;
	wire [31:0] _mesh_23_11_io_out_a_0;
	wire [31:0] _mesh_23_11_io_out_c_0;
	wire [31:0] _mesh_23_11_io_out_b_0;
	wire _mesh_23_11_io_out_control_0_dataflow;
	wire _mesh_23_11_io_out_control_0_propagate;
	wire [4:0] _mesh_23_11_io_out_control_0_shift;
	wire [2:0] _mesh_23_11_io_out_id_0;
	wire _mesh_23_11_io_out_last_0;
	wire _mesh_23_11_io_out_valid_0;
	wire [31:0] _mesh_23_10_io_out_a_0;
	wire [31:0] _mesh_23_10_io_out_c_0;
	wire [31:0] _mesh_23_10_io_out_b_0;
	wire _mesh_23_10_io_out_control_0_dataflow;
	wire _mesh_23_10_io_out_control_0_propagate;
	wire [4:0] _mesh_23_10_io_out_control_0_shift;
	wire [2:0] _mesh_23_10_io_out_id_0;
	wire _mesh_23_10_io_out_last_0;
	wire _mesh_23_10_io_out_valid_0;
	wire [31:0] _mesh_23_9_io_out_a_0;
	wire [31:0] _mesh_23_9_io_out_c_0;
	wire [31:0] _mesh_23_9_io_out_b_0;
	wire _mesh_23_9_io_out_control_0_dataflow;
	wire _mesh_23_9_io_out_control_0_propagate;
	wire [4:0] _mesh_23_9_io_out_control_0_shift;
	wire [2:0] _mesh_23_9_io_out_id_0;
	wire _mesh_23_9_io_out_last_0;
	wire _mesh_23_9_io_out_valid_0;
	wire [31:0] _mesh_23_8_io_out_a_0;
	wire [31:0] _mesh_23_8_io_out_c_0;
	wire [31:0] _mesh_23_8_io_out_b_0;
	wire _mesh_23_8_io_out_control_0_dataflow;
	wire _mesh_23_8_io_out_control_0_propagate;
	wire [4:0] _mesh_23_8_io_out_control_0_shift;
	wire [2:0] _mesh_23_8_io_out_id_0;
	wire _mesh_23_8_io_out_last_0;
	wire _mesh_23_8_io_out_valid_0;
	wire [31:0] _mesh_23_7_io_out_a_0;
	wire [31:0] _mesh_23_7_io_out_c_0;
	wire [31:0] _mesh_23_7_io_out_b_0;
	wire _mesh_23_7_io_out_control_0_dataflow;
	wire _mesh_23_7_io_out_control_0_propagate;
	wire [4:0] _mesh_23_7_io_out_control_0_shift;
	wire [2:0] _mesh_23_7_io_out_id_0;
	wire _mesh_23_7_io_out_last_0;
	wire _mesh_23_7_io_out_valid_0;
	wire [31:0] _mesh_23_6_io_out_a_0;
	wire [31:0] _mesh_23_6_io_out_c_0;
	wire [31:0] _mesh_23_6_io_out_b_0;
	wire _mesh_23_6_io_out_control_0_dataflow;
	wire _mesh_23_6_io_out_control_0_propagate;
	wire [4:0] _mesh_23_6_io_out_control_0_shift;
	wire [2:0] _mesh_23_6_io_out_id_0;
	wire _mesh_23_6_io_out_last_0;
	wire _mesh_23_6_io_out_valid_0;
	wire [31:0] _mesh_23_5_io_out_a_0;
	wire [31:0] _mesh_23_5_io_out_c_0;
	wire [31:0] _mesh_23_5_io_out_b_0;
	wire _mesh_23_5_io_out_control_0_dataflow;
	wire _mesh_23_5_io_out_control_0_propagate;
	wire [4:0] _mesh_23_5_io_out_control_0_shift;
	wire [2:0] _mesh_23_5_io_out_id_0;
	wire _mesh_23_5_io_out_last_0;
	wire _mesh_23_5_io_out_valid_0;
	wire [31:0] _mesh_23_4_io_out_a_0;
	wire [31:0] _mesh_23_4_io_out_c_0;
	wire [31:0] _mesh_23_4_io_out_b_0;
	wire _mesh_23_4_io_out_control_0_dataflow;
	wire _mesh_23_4_io_out_control_0_propagate;
	wire [4:0] _mesh_23_4_io_out_control_0_shift;
	wire [2:0] _mesh_23_4_io_out_id_0;
	wire _mesh_23_4_io_out_last_0;
	wire _mesh_23_4_io_out_valid_0;
	wire [31:0] _mesh_23_3_io_out_a_0;
	wire [31:0] _mesh_23_3_io_out_c_0;
	wire [31:0] _mesh_23_3_io_out_b_0;
	wire _mesh_23_3_io_out_control_0_dataflow;
	wire _mesh_23_3_io_out_control_0_propagate;
	wire [4:0] _mesh_23_3_io_out_control_0_shift;
	wire [2:0] _mesh_23_3_io_out_id_0;
	wire _mesh_23_3_io_out_last_0;
	wire _mesh_23_3_io_out_valid_0;
	wire [31:0] _mesh_23_2_io_out_a_0;
	wire [31:0] _mesh_23_2_io_out_c_0;
	wire [31:0] _mesh_23_2_io_out_b_0;
	wire _mesh_23_2_io_out_control_0_dataflow;
	wire _mesh_23_2_io_out_control_0_propagate;
	wire [4:0] _mesh_23_2_io_out_control_0_shift;
	wire [2:0] _mesh_23_2_io_out_id_0;
	wire _mesh_23_2_io_out_last_0;
	wire _mesh_23_2_io_out_valid_0;
	wire [31:0] _mesh_23_1_io_out_a_0;
	wire [31:0] _mesh_23_1_io_out_c_0;
	wire [31:0] _mesh_23_1_io_out_b_0;
	wire _mesh_23_1_io_out_control_0_dataflow;
	wire _mesh_23_1_io_out_control_0_propagate;
	wire [4:0] _mesh_23_1_io_out_control_0_shift;
	wire [2:0] _mesh_23_1_io_out_id_0;
	wire _mesh_23_1_io_out_last_0;
	wire _mesh_23_1_io_out_valid_0;
	wire [31:0] _mesh_23_0_io_out_a_0;
	wire [31:0] _mesh_23_0_io_out_c_0;
	wire [31:0] _mesh_23_0_io_out_b_0;
	wire _mesh_23_0_io_out_control_0_dataflow;
	wire _mesh_23_0_io_out_control_0_propagate;
	wire [4:0] _mesh_23_0_io_out_control_0_shift;
	wire [2:0] _mesh_23_0_io_out_id_0;
	wire _mesh_23_0_io_out_last_0;
	wire _mesh_23_0_io_out_valid_0;
	wire [31:0] _mesh_22_31_io_out_a_0;
	wire [31:0] _mesh_22_31_io_out_c_0;
	wire [31:0] _mesh_22_31_io_out_b_0;
	wire _mesh_22_31_io_out_control_0_dataflow;
	wire _mesh_22_31_io_out_control_0_propagate;
	wire [4:0] _mesh_22_31_io_out_control_0_shift;
	wire [2:0] _mesh_22_31_io_out_id_0;
	wire _mesh_22_31_io_out_last_0;
	wire _mesh_22_31_io_out_valid_0;
	wire [31:0] _mesh_22_30_io_out_a_0;
	wire [31:0] _mesh_22_30_io_out_c_0;
	wire [31:0] _mesh_22_30_io_out_b_0;
	wire _mesh_22_30_io_out_control_0_dataflow;
	wire _mesh_22_30_io_out_control_0_propagate;
	wire [4:0] _mesh_22_30_io_out_control_0_shift;
	wire [2:0] _mesh_22_30_io_out_id_0;
	wire _mesh_22_30_io_out_last_0;
	wire _mesh_22_30_io_out_valid_0;
	wire [31:0] _mesh_22_29_io_out_a_0;
	wire [31:0] _mesh_22_29_io_out_c_0;
	wire [31:0] _mesh_22_29_io_out_b_0;
	wire _mesh_22_29_io_out_control_0_dataflow;
	wire _mesh_22_29_io_out_control_0_propagate;
	wire [4:0] _mesh_22_29_io_out_control_0_shift;
	wire [2:0] _mesh_22_29_io_out_id_0;
	wire _mesh_22_29_io_out_last_0;
	wire _mesh_22_29_io_out_valid_0;
	wire [31:0] _mesh_22_28_io_out_a_0;
	wire [31:0] _mesh_22_28_io_out_c_0;
	wire [31:0] _mesh_22_28_io_out_b_0;
	wire _mesh_22_28_io_out_control_0_dataflow;
	wire _mesh_22_28_io_out_control_0_propagate;
	wire [4:0] _mesh_22_28_io_out_control_0_shift;
	wire [2:0] _mesh_22_28_io_out_id_0;
	wire _mesh_22_28_io_out_last_0;
	wire _mesh_22_28_io_out_valid_0;
	wire [31:0] _mesh_22_27_io_out_a_0;
	wire [31:0] _mesh_22_27_io_out_c_0;
	wire [31:0] _mesh_22_27_io_out_b_0;
	wire _mesh_22_27_io_out_control_0_dataflow;
	wire _mesh_22_27_io_out_control_0_propagate;
	wire [4:0] _mesh_22_27_io_out_control_0_shift;
	wire [2:0] _mesh_22_27_io_out_id_0;
	wire _mesh_22_27_io_out_last_0;
	wire _mesh_22_27_io_out_valid_0;
	wire [31:0] _mesh_22_26_io_out_a_0;
	wire [31:0] _mesh_22_26_io_out_c_0;
	wire [31:0] _mesh_22_26_io_out_b_0;
	wire _mesh_22_26_io_out_control_0_dataflow;
	wire _mesh_22_26_io_out_control_0_propagate;
	wire [4:0] _mesh_22_26_io_out_control_0_shift;
	wire [2:0] _mesh_22_26_io_out_id_0;
	wire _mesh_22_26_io_out_last_0;
	wire _mesh_22_26_io_out_valid_0;
	wire [31:0] _mesh_22_25_io_out_a_0;
	wire [31:0] _mesh_22_25_io_out_c_0;
	wire [31:0] _mesh_22_25_io_out_b_0;
	wire _mesh_22_25_io_out_control_0_dataflow;
	wire _mesh_22_25_io_out_control_0_propagate;
	wire [4:0] _mesh_22_25_io_out_control_0_shift;
	wire [2:0] _mesh_22_25_io_out_id_0;
	wire _mesh_22_25_io_out_last_0;
	wire _mesh_22_25_io_out_valid_0;
	wire [31:0] _mesh_22_24_io_out_a_0;
	wire [31:0] _mesh_22_24_io_out_c_0;
	wire [31:0] _mesh_22_24_io_out_b_0;
	wire _mesh_22_24_io_out_control_0_dataflow;
	wire _mesh_22_24_io_out_control_0_propagate;
	wire [4:0] _mesh_22_24_io_out_control_0_shift;
	wire [2:0] _mesh_22_24_io_out_id_0;
	wire _mesh_22_24_io_out_last_0;
	wire _mesh_22_24_io_out_valid_0;
	wire [31:0] _mesh_22_23_io_out_a_0;
	wire [31:0] _mesh_22_23_io_out_c_0;
	wire [31:0] _mesh_22_23_io_out_b_0;
	wire _mesh_22_23_io_out_control_0_dataflow;
	wire _mesh_22_23_io_out_control_0_propagate;
	wire [4:0] _mesh_22_23_io_out_control_0_shift;
	wire [2:0] _mesh_22_23_io_out_id_0;
	wire _mesh_22_23_io_out_last_0;
	wire _mesh_22_23_io_out_valid_0;
	wire [31:0] _mesh_22_22_io_out_a_0;
	wire [31:0] _mesh_22_22_io_out_c_0;
	wire [31:0] _mesh_22_22_io_out_b_0;
	wire _mesh_22_22_io_out_control_0_dataflow;
	wire _mesh_22_22_io_out_control_0_propagate;
	wire [4:0] _mesh_22_22_io_out_control_0_shift;
	wire [2:0] _mesh_22_22_io_out_id_0;
	wire _mesh_22_22_io_out_last_0;
	wire _mesh_22_22_io_out_valid_0;
	wire [31:0] _mesh_22_21_io_out_a_0;
	wire [31:0] _mesh_22_21_io_out_c_0;
	wire [31:0] _mesh_22_21_io_out_b_0;
	wire _mesh_22_21_io_out_control_0_dataflow;
	wire _mesh_22_21_io_out_control_0_propagate;
	wire [4:0] _mesh_22_21_io_out_control_0_shift;
	wire [2:0] _mesh_22_21_io_out_id_0;
	wire _mesh_22_21_io_out_last_0;
	wire _mesh_22_21_io_out_valid_0;
	wire [31:0] _mesh_22_20_io_out_a_0;
	wire [31:0] _mesh_22_20_io_out_c_0;
	wire [31:0] _mesh_22_20_io_out_b_0;
	wire _mesh_22_20_io_out_control_0_dataflow;
	wire _mesh_22_20_io_out_control_0_propagate;
	wire [4:0] _mesh_22_20_io_out_control_0_shift;
	wire [2:0] _mesh_22_20_io_out_id_0;
	wire _mesh_22_20_io_out_last_0;
	wire _mesh_22_20_io_out_valid_0;
	wire [31:0] _mesh_22_19_io_out_a_0;
	wire [31:0] _mesh_22_19_io_out_c_0;
	wire [31:0] _mesh_22_19_io_out_b_0;
	wire _mesh_22_19_io_out_control_0_dataflow;
	wire _mesh_22_19_io_out_control_0_propagate;
	wire [4:0] _mesh_22_19_io_out_control_0_shift;
	wire [2:0] _mesh_22_19_io_out_id_0;
	wire _mesh_22_19_io_out_last_0;
	wire _mesh_22_19_io_out_valid_0;
	wire [31:0] _mesh_22_18_io_out_a_0;
	wire [31:0] _mesh_22_18_io_out_c_0;
	wire [31:0] _mesh_22_18_io_out_b_0;
	wire _mesh_22_18_io_out_control_0_dataflow;
	wire _mesh_22_18_io_out_control_0_propagate;
	wire [4:0] _mesh_22_18_io_out_control_0_shift;
	wire [2:0] _mesh_22_18_io_out_id_0;
	wire _mesh_22_18_io_out_last_0;
	wire _mesh_22_18_io_out_valid_0;
	wire [31:0] _mesh_22_17_io_out_a_0;
	wire [31:0] _mesh_22_17_io_out_c_0;
	wire [31:0] _mesh_22_17_io_out_b_0;
	wire _mesh_22_17_io_out_control_0_dataflow;
	wire _mesh_22_17_io_out_control_0_propagate;
	wire [4:0] _mesh_22_17_io_out_control_0_shift;
	wire [2:0] _mesh_22_17_io_out_id_0;
	wire _mesh_22_17_io_out_last_0;
	wire _mesh_22_17_io_out_valid_0;
	wire [31:0] _mesh_22_16_io_out_a_0;
	wire [31:0] _mesh_22_16_io_out_c_0;
	wire [31:0] _mesh_22_16_io_out_b_0;
	wire _mesh_22_16_io_out_control_0_dataflow;
	wire _mesh_22_16_io_out_control_0_propagate;
	wire [4:0] _mesh_22_16_io_out_control_0_shift;
	wire [2:0] _mesh_22_16_io_out_id_0;
	wire _mesh_22_16_io_out_last_0;
	wire _mesh_22_16_io_out_valid_0;
	wire [31:0] _mesh_22_15_io_out_a_0;
	wire [31:0] _mesh_22_15_io_out_c_0;
	wire [31:0] _mesh_22_15_io_out_b_0;
	wire _mesh_22_15_io_out_control_0_dataflow;
	wire _mesh_22_15_io_out_control_0_propagate;
	wire [4:0] _mesh_22_15_io_out_control_0_shift;
	wire [2:0] _mesh_22_15_io_out_id_0;
	wire _mesh_22_15_io_out_last_0;
	wire _mesh_22_15_io_out_valid_0;
	wire [31:0] _mesh_22_14_io_out_a_0;
	wire [31:0] _mesh_22_14_io_out_c_0;
	wire [31:0] _mesh_22_14_io_out_b_0;
	wire _mesh_22_14_io_out_control_0_dataflow;
	wire _mesh_22_14_io_out_control_0_propagate;
	wire [4:0] _mesh_22_14_io_out_control_0_shift;
	wire [2:0] _mesh_22_14_io_out_id_0;
	wire _mesh_22_14_io_out_last_0;
	wire _mesh_22_14_io_out_valid_0;
	wire [31:0] _mesh_22_13_io_out_a_0;
	wire [31:0] _mesh_22_13_io_out_c_0;
	wire [31:0] _mesh_22_13_io_out_b_0;
	wire _mesh_22_13_io_out_control_0_dataflow;
	wire _mesh_22_13_io_out_control_0_propagate;
	wire [4:0] _mesh_22_13_io_out_control_0_shift;
	wire [2:0] _mesh_22_13_io_out_id_0;
	wire _mesh_22_13_io_out_last_0;
	wire _mesh_22_13_io_out_valid_0;
	wire [31:0] _mesh_22_12_io_out_a_0;
	wire [31:0] _mesh_22_12_io_out_c_0;
	wire [31:0] _mesh_22_12_io_out_b_0;
	wire _mesh_22_12_io_out_control_0_dataflow;
	wire _mesh_22_12_io_out_control_0_propagate;
	wire [4:0] _mesh_22_12_io_out_control_0_shift;
	wire [2:0] _mesh_22_12_io_out_id_0;
	wire _mesh_22_12_io_out_last_0;
	wire _mesh_22_12_io_out_valid_0;
	wire [31:0] _mesh_22_11_io_out_a_0;
	wire [31:0] _mesh_22_11_io_out_c_0;
	wire [31:0] _mesh_22_11_io_out_b_0;
	wire _mesh_22_11_io_out_control_0_dataflow;
	wire _mesh_22_11_io_out_control_0_propagate;
	wire [4:0] _mesh_22_11_io_out_control_0_shift;
	wire [2:0] _mesh_22_11_io_out_id_0;
	wire _mesh_22_11_io_out_last_0;
	wire _mesh_22_11_io_out_valid_0;
	wire [31:0] _mesh_22_10_io_out_a_0;
	wire [31:0] _mesh_22_10_io_out_c_0;
	wire [31:0] _mesh_22_10_io_out_b_0;
	wire _mesh_22_10_io_out_control_0_dataflow;
	wire _mesh_22_10_io_out_control_0_propagate;
	wire [4:0] _mesh_22_10_io_out_control_0_shift;
	wire [2:0] _mesh_22_10_io_out_id_0;
	wire _mesh_22_10_io_out_last_0;
	wire _mesh_22_10_io_out_valid_0;
	wire [31:0] _mesh_22_9_io_out_a_0;
	wire [31:0] _mesh_22_9_io_out_c_0;
	wire [31:0] _mesh_22_9_io_out_b_0;
	wire _mesh_22_9_io_out_control_0_dataflow;
	wire _mesh_22_9_io_out_control_0_propagate;
	wire [4:0] _mesh_22_9_io_out_control_0_shift;
	wire [2:0] _mesh_22_9_io_out_id_0;
	wire _mesh_22_9_io_out_last_0;
	wire _mesh_22_9_io_out_valid_0;
	wire [31:0] _mesh_22_8_io_out_a_0;
	wire [31:0] _mesh_22_8_io_out_c_0;
	wire [31:0] _mesh_22_8_io_out_b_0;
	wire _mesh_22_8_io_out_control_0_dataflow;
	wire _mesh_22_8_io_out_control_0_propagate;
	wire [4:0] _mesh_22_8_io_out_control_0_shift;
	wire [2:0] _mesh_22_8_io_out_id_0;
	wire _mesh_22_8_io_out_last_0;
	wire _mesh_22_8_io_out_valid_0;
	wire [31:0] _mesh_22_7_io_out_a_0;
	wire [31:0] _mesh_22_7_io_out_c_0;
	wire [31:0] _mesh_22_7_io_out_b_0;
	wire _mesh_22_7_io_out_control_0_dataflow;
	wire _mesh_22_7_io_out_control_0_propagate;
	wire [4:0] _mesh_22_7_io_out_control_0_shift;
	wire [2:0] _mesh_22_7_io_out_id_0;
	wire _mesh_22_7_io_out_last_0;
	wire _mesh_22_7_io_out_valid_0;
	wire [31:0] _mesh_22_6_io_out_a_0;
	wire [31:0] _mesh_22_6_io_out_c_0;
	wire [31:0] _mesh_22_6_io_out_b_0;
	wire _mesh_22_6_io_out_control_0_dataflow;
	wire _mesh_22_6_io_out_control_0_propagate;
	wire [4:0] _mesh_22_6_io_out_control_0_shift;
	wire [2:0] _mesh_22_6_io_out_id_0;
	wire _mesh_22_6_io_out_last_0;
	wire _mesh_22_6_io_out_valid_0;
	wire [31:0] _mesh_22_5_io_out_a_0;
	wire [31:0] _mesh_22_5_io_out_c_0;
	wire [31:0] _mesh_22_5_io_out_b_0;
	wire _mesh_22_5_io_out_control_0_dataflow;
	wire _mesh_22_5_io_out_control_0_propagate;
	wire [4:0] _mesh_22_5_io_out_control_0_shift;
	wire [2:0] _mesh_22_5_io_out_id_0;
	wire _mesh_22_5_io_out_last_0;
	wire _mesh_22_5_io_out_valid_0;
	wire [31:0] _mesh_22_4_io_out_a_0;
	wire [31:0] _mesh_22_4_io_out_c_0;
	wire [31:0] _mesh_22_4_io_out_b_0;
	wire _mesh_22_4_io_out_control_0_dataflow;
	wire _mesh_22_4_io_out_control_0_propagate;
	wire [4:0] _mesh_22_4_io_out_control_0_shift;
	wire [2:0] _mesh_22_4_io_out_id_0;
	wire _mesh_22_4_io_out_last_0;
	wire _mesh_22_4_io_out_valid_0;
	wire [31:0] _mesh_22_3_io_out_a_0;
	wire [31:0] _mesh_22_3_io_out_c_0;
	wire [31:0] _mesh_22_3_io_out_b_0;
	wire _mesh_22_3_io_out_control_0_dataflow;
	wire _mesh_22_3_io_out_control_0_propagate;
	wire [4:0] _mesh_22_3_io_out_control_0_shift;
	wire [2:0] _mesh_22_3_io_out_id_0;
	wire _mesh_22_3_io_out_last_0;
	wire _mesh_22_3_io_out_valid_0;
	wire [31:0] _mesh_22_2_io_out_a_0;
	wire [31:0] _mesh_22_2_io_out_c_0;
	wire [31:0] _mesh_22_2_io_out_b_0;
	wire _mesh_22_2_io_out_control_0_dataflow;
	wire _mesh_22_2_io_out_control_0_propagate;
	wire [4:0] _mesh_22_2_io_out_control_0_shift;
	wire [2:0] _mesh_22_2_io_out_id_0;
	wire _mesh_22_2_io_out_last_0;
	wire _mesh_22_2_io_out_valid_0;
	wire [31:0] _mesh_22_1_io_out_a_0;
	wire [31:0] _mesh_22_1_io_out_c_0;
	wire [31:0] _mesh_22_1_io_out_b_0;
	wire _mesh_22_1_io_out_control_0_dataflow;
	wire _mesh_22_1_io_out_control_0_propagate;
	wire [4:0] _mesh_22_1_io_out_control_0_shift;
	wire [2:0] _mesh_22_1_io_out_id_0;
	wire _mesh_22_1_io_out_last_0;
	wire _mesh_22_1_io_out_valid_0;
	wire [31:0] _mesh_22_0_io_out_a_0;
	wire [31:0] _mesh_22_0_io_out_c_0;
	wire [31:0] _mesh_22_0_io_out_b_0;
	wire _mesh_22_0_io_out_control_0_dataflow;
	wire _mesh_22_0_io_out_control_0_propagate;
	wire [4:0] _mesh_22_0_io_out_control_0_shift;
	wire [2:0] _mesh_22_0_io_out_id_0;
	wire _mesh_22_0_io_out_last_0;
	wire _mesh_22_0_io_out_valid_0;
	wire [31:0] _mesh_21_31_io_out_a_0;
	wire [31:0] _mesh_21_31_io_out_c_0;
	wire [31:0] _mesh_21_31_io_out_b_0;
	wire _mesh_21_31_io_out_control_0_dataflow;
	wire _mesh_21_31_io_out_control_0_propagate;
	wire [4:0] _mesh_21_31_io_out_control_0_shift;
	wire [2:0] _mesh_21_31_io_out_id_0;
	wire _mesh_21_31_io_out_last_0;
	wire _mesh_21_31_io_out_valid_0;
	wire [31:0] _mesh_21_30_io_out_a_0;
	wire [31:0] _mesh_21_30_io_out_c_0;
	wire [31:0] _mesh_21_30_io_out_b_0;
	wire _mesh_21_30_io_out_control_0_dataflow;
	wire _mesh_21_30_io_out_control_0_propagate;
	wire [4:0] _mesh_21_30_io_out_control_0_shift;
	wire [2:0] _mesh_21_30_io_out_id_0;
	wire _mesh_21_30_io_out_last_0;
	wire _mesh_21_30_io_out_valid_0;
	wire [31:0] _mesh_21_29_io_out_a_0;
	wire [31:0] _mesh_21_29_io_out_c_0;
	wire [31:0] _mesh_21_29_io_out_b_0;
	wire _mesh_21_29_io_out_control_0_dataflow;
	wire _mesh_21_29_io_out_control_0_propagate;
	wire [4:0] _mesh_21_29_io_out_control_0_shift;
	wire [2:0] _mesh_21_29_io_out_id_0;
	wire _mesh_21_29_io_out_last_0;
	wire _mesh_21_29_io_out_valid_0;
	wire [31:0] _mesh_21_28_io_out_a_0;
	wire [31:0] _mesh_21_28_io_out_c_0;
	wire [31:0] _mesh_21_28_io_out_b_0;
	wire _mesh_21_28_io_out_control_0_dataflow;
	wire _mesh_21_28_io_out_control_0_propagate;
	wire [4:0] _mesh_21_28_io_out_control_0_shift;
	wire [2:0] _mesh_21_28_io_out_id_0;
	wire _mesh_21_28_io_out_last_0;
	wire _mesh_21_28_io_out_valid_0;
	wire [31:0] _mesh_21_27_io_out_a_0;
	wire [31:0] _mesh_21_27_io_out_c_0;
	wire [31:0] _mesh_21_27_io_out_b_0;
	wire _mesh_21_27_io_out_control_0_dataflow;
	wire _mesh_21_27_io_out_control_0_propagate;
	wire [4:0] _mesh_21_27_io_out_control_0_shift;
	wire [2:0] _mesh_21_27_io_out_id_0;
	wire _mesh_21_27_io_out_last_0;
	wire _mesh_21_27_io_out_valid_0;
	wire [31:0] _mesh_21_26_io_out_a_0;
	wire [31:0] _mesh_21_26_io_out_c_0;
	wire [31:0] _mesh_21_26_io_out_b_0;
	wire _mesh_21_26_io_out_control_0_dataflow;
	wire _mesh_21_26_io_out_control_0_propagate;
	wire [4:0] _mesh_21_26_io_out_control_0_shift;
	wire [2:0] _mesh_21_26_io_out_id_0;
	wire _mesh_21_26_io_out_last_0;
	wire _mesh_21_26_io_out_valid_0;
	wire [31:0] _mesh_21_25_io_out_a_0;
	wire [31:0] _mesh_21_25_io_out_c_0;
	wire [31:0] _mesh_21_25_io_out_b_0;
	wire _mesh_21_25_io_out_control_0_dataflow;
	wire _mesh_21_25_io_out_control_0_propagate;
	wire [4:0] _mesh_21_25_io_out_control_0_shift;
	wire [2:0] _mesh_21_25_io_out_id_0;
	wire _mesh_21_25_io_out_last_0;
	wire _mesh_21_25_io_out_valid_0;
	wire [31:0] _mesh_21_24_io_out_a_0;
	wire [31:0] _mesh_21_24_io_out_c_0;
	wire [31:0] _mesh_21_24_io_out_b_0;
	wire _mesh_21_24_io_out_control_0_dataflow;
	wire _mesh_21_24_io_out_control_0_propagate;
	wire [4:0] _mesh_21_24_io_out_control_0_shift;
	wire [2:0] _mesh_21_24_io_out_id_0;
	wire _mesh_21_24_io_out_last_0;
	wire _mesh_21_24_io_out_valid_0;
	wire [31:0] _mesh_21_23_io_out_a_0;
	wire [31:0] _mesh_21_23_io_out_c_0;
	wire [31:0] _mesh_21_23_io_out_b_0;
	wire _mesh_21_23_io_out_control_0_dataflow;
	wire _mesh_21_23_io_out_control_0_propagate;
	wire [4:0] _mesh_21_23_io_out_control_0_shift;
	wire [2:0] _mesh_21_23_io_out_id_0;
	wire _mesh_21_23_io_out_last_0;
	wire _mesh_21_23_io_out_valid_0;
	wire [31:0] _mesh_21_22_io_out_a_0;
	wire [31:0] _mesh_21_22_io_out_c_0;
	wire [31:0] _mesh_21_22_io_out_b_0;
	wire _mesh_21_22_io_out_control_0_dataflow;
	wire _mesh_21_22_io_out_control_0_propagate;
	wire [4:0] _mesh_21_22_io_out_control_0_shift;
	wire [2:0] _mesh_21_22_io_out_id_0;
	wire _mesh_21_22_io_out_last_0;
	wire _mesh_21_22_io_out_valid_0;
	wire [31:0] _mesh_21_21_io_out_a_0;
	wire [31:0] _mesh_21_21_io_out_c_0;
	wire [31:0] _mesh_21_21_io_out_b_0;
	wire _mesh_21_21_io_out_control_0_dataflow;
	wire _mesh_21_21_io_out_control_0_propagate;
	wire [4:0] _mesh_21_21_io_out_control_0_shift;
	wire [2:0] _mesh_21_21_io_out_id_0;
	wire _mesh_21_21_io_out_last_0;
	wire _mesh_21_21_io_out_valid_0;
	wire [31:0] _mesh_21_20_io_out_a_0;
	wire [31:0] _mesh_21_20_io_out_c_0;
	wire [31:0] _mesh_21_20_io_out_b_0;
	wire _mesh_21_20_io_out_control_0_dataflow;
	wire _mesh_21_20_io_out_control_0_propagate;
	wire [4:0] _mesh_21_20_io_out_control_0_shift;
	wire [2:0] _mesh_21_20_io_out_id_0;
	wire _mesh_21_20_io_out_last_0;
	wire _mesh_21_20_io_out_valid_0;
	wire [31:0] _mesh_21_19_io_out_a_0;
	wire [31:0] _mesh_21_19_io_out_c_0;
	wire [31:0] _mesh_21_19_io_out_b_0;
	wire _mesh_21_19_io_out_control_0_dataflow;
	wire _mesh_21_19_io_out_control_0_propagate;
	wire [4:0] _mesh_21_19_io_out_control_0_shift;
	wire [2:0] _mesh_21_19_io_out_id_0;
	wire _mesh_21_19_io_out_last_0;
	wire _mesh_21_19_io_out_valid_0;
	wire [31:0] _mesh_21_18_io_out_a_0;
	wire [31:0] _mesh_21_18_io_out_c_0;
	wire [31:0] _mesh_21_18_io_out_b_0;
	wire _mesh_21_18_io_out_control_0_dataflow;
	wire _mesh_21_18_io_out_control_0_propagate;
	wire [4:0] _mesh_21_18_io_out_control_0_shift;
	wire [2:0] _mesh_21_18_io_out_id_0;
	wire _mesh_21_18_io_out_last_0;
	wire _mesh_21_18_io_out_valid_0;
	wire [31:0] _mesh_21_17_io_out_a_0;
	wire [31:0] _mesh_21_17_io_out_c_0;
	wire [31:0] _mesh_21_17_io_out_b_0;
	wire _mesh_21_17_io_out_control_0_dataflow;
	wire _mesh_21_17_io_out_control_0_propagate;
	wire [4:0] _mesh_21_17_io_out_control_0_shift;
	wire [2:0] _mesh_21_17_io_out_id_0;
	wire _mesh_21_17_io_out_last_0;
	wire _mesh_21_17_io_out_valid_0;
	wire [31:0] _mesh_21_16_io_out_a_0;
	wire [31:0] _mesh_21_16_io_out_c_0;
	wire [31:0] _mesh_21_16_io_out_b_0;
	wire _mesh_21_16_io_out_control_0_dataflow;
	wire _mesh_21_16_io_out_control_0_propagate;
	wire [4:0] _mesh_21_16_io_out_control_0_shift;
	wire [2:0] _mesh_21_16_io_out_id_0;
	wire _mesh_21_16_io_out_last_0;
	wire _mesh_21_16_io_out_valid_0;
	wire [31:0] _mesh_21_15_io_out_a_0;
	wire [31:0] _mesh_21_15_io_out_c_0;
	wire [31:0] _mesh_21_15_io_out_b_0;
	wire _mesh_21_15_io_out_control_0_dataflow;
	wire _mesh_21_15_io_out_control_0_propagate;
	wire [4:0] _mesh_21_15_io_out_control_0_shift;
	wire [2:0] _mesh_21_15_io_out_id_0;
	wire _mesh_21_15_io_out_last_0;
	wire _mesh_21_15_io_out_valid_0;
	wire [31:0] _mesh_21_14_io_out_a_0;
	wire [31:0] _mesh_21_14_io_out_c_0;
	wire [31:0] _mesh_21_14_io_out_b_0;
	wire _mesh_21_14_io_out_control_0_dataflow;
	wire _mesh_21_14_io_out_control_0_propagate;
	wire [4:0] _mesh_21_14_io_out_control_0_shift;
	wire [2:0] _mesh_21_14_io_out_id_0;
	wire _mesh_21_14_io_out_last_0;
	wire _mesh_21_14_io_out_valid_0;
	wire [31:0] _mesh_21_13_io_out_a_0;
	wire [31:0] _mesh_21_13_io_out_c_0;
	wire [31:0] _mesh_21_13_io_out_b_0;
	wire _mesh_21_13_io_out_control_0_dataflow;
	wire _mesh_21_13_io_out_control_0_propagate;
	wire [4:0] _mesh_21_13_io_out_control_0_shift;
	wire [2:0] _mesh_21_13_io_out_id_0;
	wire _mesh_21_13_io_out_last_0;
	wire _mesh_21_13_io_out_valid_0;
	wire [31:0] _mesh_21_12_io_out_a_0;
	wire [31:0] _mesh_21_12_io_out_c_0;
	wire [31:0] _mesh_21_12_io_out_b_0;
	wire _mesh_21_12_io_out_control_0_dataflow;
	wire _mesh_21_12_io_out_control_0_propagate;
	wire [4:0] _mesh_21_12_io_out_control_0_shift;
	wire [2:0] _mesh_21_12_io_out_id_0;
	wire _mesh_21_12_io_out_last_0;
	wire _mesh_21_12_io_out_valid_0;
	wire [31:0] _mesh_21_11_io_out_a_0;
	wire [31:0] _mesh_21_11_io_out_c_0;
	wire [31:0] _mesh_21_11_io_out_b_0;
	wire _mesh_21_11_io_out_control_0_dataflow;
	wire _mesh_21_11_io_out_control_0_propagate;
	wire [4:0] _mesh_21_11_io_out_control_0_shift;
	wire [2:0] _mesh_21_11_io_out_id_0;
	wire _mesh_21_11_io_out_last_0;
	wire _mesh_21_11_io_out_valid_0;
	wire [31:0] _mesh_21_10_io_out_a_0;
	wire [31:0] _mesh_21_10_io_out_c_0;
	wire [31:0] _mesh_21_10_io_out_b_0;
	wire _mesh_21_10_io_out_control_0_dataflow;
	wire _mesh_21_10_io_out_control_0_propagate;
	wire [4:0] _mesh_21_10_io_out_control_0_shift;
	wire [2:0] _mesh_21_10_io_out_id_0;
	wire _mesh_21_10_io_out_last_0;
	wire _mesh_21_10_io_out_valid_0;
	wire [31:0] _mesh_21_9_io_out_a_0;
	wire [31:0] _mesh_21_9_io_out_c_0;
	wire [31:0] _mesh_21_9_io_out_b_0;
	wire _mesh_21_9_io_out_control_0_dataflow;
	wire _mesh_21_9_io_out_control_0_propagate;
	wire [4:0] _mesh_21_9_io_out_control_0_shift;
	wire [2:0] _mesh_21_9_io_out_id_0;
	wire _mesh_21_9_io_out_last_0;
	wire _mesh_21_9_io_out_valid_0;
	wire [31:0] _mesh_21_8_io_out_a_0;
	wire [31:0] _mesh_21_8_io_out_c_0;
	wire [31:0] _mesh_21_8_io_out_b_0;
	wire _mesh_21_8_io_out_control_0_dataflow;
	wire _mesh_21_8_io_out_control_0_propagate;
	wire [4:0] _mesh_21_8_io_out_control_0_shift;
	wire [2:0] _mesh_21_8_io_out_id_0;
	wire _mesh_21_8_io_out_last_0;
	wire _mesh_21_8_io_out_valid_0;
	wire [31:0] _mesh_21_7_io_out_a_0;
	wire [31:0] _mesh_21_7_io_out_c_0;
	wire [31:0] _mesh_21_7_io_out_b_0;
	wire _mesh_21_7_io_out_control_0_dataflow;
	wire _mesh_21_7_io_out_control_0_propagate;
	wire [4:0] _mesh_21_7_io_out_control_0_shift;
	wire [2:0] _mesh_21_7_io_out_id_0;
	wire _mesh_21_7_io_out_last_0;
	wire _mesh_21_7_io_out_valid_0;
	wire [31:0] _mesh_21_6_io_out_a_0;
	wire [31:0] _mesh_21_6_io_out_c_0;
	wire [31:0] _mesh_21_6_io_out_b_0;
	wire _mesh_21_6_io_out_control_0_dataflow;
	wire _mesh_21_6_io_out_control_0_propagate;
	wire [4:0] _mesh_21_6_io_out_control_0_shift;
	wire [2:0] _mesh_21_6_io_out_id_0;
	wire _mesh_21_6_io_out_last_0;
	wire _mesh_21_6_io_out_valid_0;
	wire [31:0] _mesh_21_5_io_out_a_0;
	wire [31:0] _mesh_21_5_io_out_c_0;
	wire [31:0] _mesh_21_5_io_out_b_0;
	wire _mesh_21_5_io_out_control_0_dataflow;
	wire _mesh_21_5_io_out_control_0_propagate;
	wire [4:0] _mesh_21_5_io_out_control_0_shift;
	wire [2:0] _mesh_21_5_io_out_id_0;
	wire _mesh_21_5_io_out_last_0;
	wire _mesh_21_5_io_out_valid_0;
	wire [31:0] _mesh_21_4_io_out_a_0;
	wire [31:0] _mesh_21_4_io_out_c_0;
	wire [31:0] _mesh_21_4_io_out_b_0;
	wire _mesh_21_4_io_out_control_0_dataflow;
	wire _mesh_21_4_io_out_control_0_propagate;
	wire [4:0] _mesh_21_4_io_out_control_0_shift;
	wire [2:0] _mesh_21_4_io_out_id_0;
	wire _mesh_21_4_io_out_last_0;
	wire _mesh_21_4_io_out_valid_0;
	wire [31:0] _mesh_21_3_io_out_a_0;
	wire [31:0] _mesh_21_3_io_out_c_0;
	wire [31:0] _mesh_21_3_io_out_b_0;
	wire _mesh_21_3_io_out_control_0_dataflow;
	wire _mesh_21_3_io_out_control_0_propagate;
	wire [4:0] _mesh_21_3_io_out_control_0_shift;
	wire [2:0] _mesh_21_3_io_out_id_0;
	wire _mesh_21_3_io_out_last_0;
	wire _mesh_21_3_io_out_valid_0;
	wire [31:0] _mesh_21_2_io_out_a_0;
	wire [31:0] _mesh_21_2_io_out_c_0;
	wire [31:0] _mesh_21_2_io_out_b_0;
	wire _mesh_21_2_io_out_control_0_dataflow;
	wire _mesh_21_2_io_out_control_0_propagate;
	wire [4:0] _mesh_21_2_io_out_control_0_shift;
	wire [2:0] _mesh_21_2_io_out_id_0;
	wire _mesh_21_2_io_out_last_0;
	wire _mesh_21_2_io_out_valid_0;
	wire [31:0] _mesh_21_1_io_out_a_0;
	wire [31:0] _mesh_21_1_io_out_c_0;
	wire [31:0] _mesh_21_1_io_out_b_0;
	wire _mesh_21_1_io_out_control_0_dataflow;
	wire _mesh_21_1_io_out_control_0_propagate;
	wire [4:0] _mesh_21_1_io_out_control_0_shift;
	wire [2:0] _mesh_21_1_io_out_id_0;
	wire _mesh_21_1_io_out_last_0;
	wire _mesh_21_1_io_out_valid_0;
	wire [31:0] _mesh_21_0_io_out_a_0;
	wire [31:0] _mesh_21_0_io_out_c_0;
	wire [31:0] _mesh_21_0_io_out_b_0;
	wire _mesh_21_0_io_out_control_0_dataflow;
	wire _mesh_21_0_io_out_control_0_propagate;
	wire [4:0] _mesh_21_0_io_out_control_0_shift;
	wire [2:0] _mesh_21_0_io_out_id_0;
	wire _mesh_21_0_io_out_last_0;
	wire _mesh_21_0_io_out_valid_0;
	wire [31:0] _mesh_20_31_io_out_a_0;
	wire [31:0] _mesh_20_31_io_out_c_0;
	wire [31:0] _mesh_20_31_io_out_b_0;
	wire _mesh_20_31_io_out_control_0_dataflow;
	wire _mesh_20_31_io_out_control_0_propagate;
	wire [4:0] _mesh_20_31_io_out_control_0_shift;
	wire [2:0] _mesh_20_31_io_out_id_0;
	wire _mesh_20_31_io_out_last_0;
	wire _mesh_20_31_io_out_valid_0;
	wire [31:0] _mesh_20_30_io_out_a_0;
	wire [31:0] _mesh_20_30_io_out_c_0;
	wire [31:0] _mesh_20_30_io_out_b_0;
	wire _mesh_20_30_io_out_control_0_dataflow;
	wire _mesh_20_30_io_out_control_0_propagate;
	wire [4:0] _mesh_20_30_io_out_control_0_shift;
	wire [2:0] _mesh_20_30_io_out_id_0;
	wire _mesh_20_30_io_out_last_0;
	wire _mesh_20_30_io_out_valid_0;
	wire [31:0] _mesh_20_29_io_out_a_0;
	wire [31:0] _mesh_20_29_io_out_c_0;
	wire [31:0] _mesh_20_29_io_out_b_0;
	wire _mesh_20_29_io_out_control_0_dataflow;
	wire _mesh_20_29_io_out_control_0_propagate;
	wire [4:0] _mesh_20_29_io_out_control_0_shift;
	wire [2:0] _mesh_20_29_io_out_id_0;
	wire _mesh_20_29_io_out_last_0;
	wire _mesh_20_29_io_out_valid_0;
	wire [31:0] _mesh_20_28_io_out_a_0;
	wire [31:0] _mesh_20_28_io_out_c_0;
	wire [31:0] _mesh_20_28_io_out_b_0;
	wire _mesh_20_28_io_out_control_0_dataflow;
	wire _mesh_20_28_io_out_control_0_propagate;
	wire [4:0] _mesh_20_28_io_out_control_0_shift;
	wire [2:0] _mesh_20_28_io_out_id_0;
	wire _mesh_20_28_io_out_last_0;
	wire _mesh_20_28_io_out_valid_0;
	wire [31:0] _mesh_20_27_io_out_a_0;
	wire [31:0] _mesh_20_27_io_out_c_0;
	wire [31:0] _mesh_20_27_io_out_b_0;
	wire _mesh_20_27_io_out_control_0_dataflow;
	wire _mesh_20_27_io_out_control_0_propagate;
	wire [4:0] _mesh_20_27_io_out_control_0_shift;
	wire [2:0] _mesh_20_27_io_out_id_0;
	wire _mesh_20_27_io_out_last_0;
	wire _mesh_20_27_io_out_valid_0;
	wire [31:0] _mesh_20_26_io_out_a_0;
	wire [31:0] _mesh_20_26_io_out_c_0;
	wire [31:0] _mesh_20_26_io_out_b_0;
	wire _mesh_20_26_io_out_control_0_dataflow;
	wire _mesh_20_26_io_out_control_0_propagate;
	wire [4:0] _mesh_20_26_io_out_control_0_shift;
	wire [2:0] _mesh_20_26_io_out_id_0;
	wire _mesh_20_26_io_out_last_0;
	wire _mesh_20_26_io_out_valid_0;
	wire [31:0] _mesh_20_25_io_out_a_0;
	wire [31:0] _mesh_20_25_io_out_c_0;
	wire [31:0] _mesh_20_25_io_out_b_0;
	wire _mesh_20_25_io_out_control_0_dataflow;
	wire _mesh_20_25_io_out_control_0_propagate;
	wire [4:0] _mesh_20_25_io_out_control_0_shift;
	wire [2:0] _mesh_20_25_io_out_id_0;
	wire _mesh_20_25_io_out_last_0;
	wire _mesh_20_25_io_out_valid_0;
	wire [31:0] _mesh_20_24_io_out_a_0;
	wire [31:0] _mesh_20_24_io_out_c_0;
	wire [31:0] _mesh_20_24_io_out_b_0;
	wire _mesh_20_24_io_out_control_0_dataflow;
	wire _mesh_20_24_io_out_control_0_propagate;
	wire [4:0] _mesh_20_24_io_out_control_0_shift;
	wire [2:0] _mesh_20_24_io_out_id_0;
	wire _mesh_20_24_io_out_last_0;
	wire _mesh_20_24_io_out_valid_0;
	wire [31:0] _mesh_20_23_io_out_a_0;
	wire [31:0] _mesh_20_23_io_out_c_0;
	wire [31:0] _mesh_20_23_io_out_b_0;
	wire _mesh_20_23_io_out_control_0_dataflow;
	wire _mesh_20_23_io_out_control_0_propagate;
	wire [4:0] _mesh_20_23_io_out_control_0_shift;
	wire [2:0] _mesh_20_23_io_out_id_0;
	wire _mesh_20_23_io_out_last_0;
	wire _mesh_20_23_io_out_valid_0;
	wire [31:0] _mesh_20_22_io_out_a_0;
	wire [31:0] _mesh_20_22_io_out_c_0;
	wire [31:0] _mesh_20_22_io_out_b_0;
	wire _mesh_20_22_io_out_control_0_dataflow;
	wire _mesh_20_22_io_out_control_0_propagate;
	wire [4:0] _mesh_20_22_io_out_control_0_shift;
	wire [2:0] _mesh_20_22_io_out_id_0;
	wire _mesh_20_22_io_out_last_0;
	wire _mesh_20_22_io_out_valid_0;
	wire [31:0] _mesh_20_21_io_out_a_0;
	wire [31:0] _mesh_20_21_io_out_c_0;
	wire [31:0] _mesh_20_21_io_out_b_0;
	wire _mesh_20_21_io_out_control_0_dataflow;
	wire _mesh_20_21_io_out_control_0_propagate;
	wire [4:0] _mesh_20_21_io_out_control_0_shift;
	wire [2:0] _mesh_20_21_io_out_id_0;
	wire _mesh_20_21_io_out_last_0;
	wire _mesh_20_21_io_out_valid_0;
	wire [31:0] _mesh_20_20_io_out_a_0;
	wire [31:0] _mesh_20_20_io_out_c_0;
	wire [31:0] _mesh_20_20_io_out_b_0;
	wire _mesh_20_20_io_out_control_0_dataflow;
	wire _mesh_20_20_io_out_control_0_propagate;
	wire [4:0] _mesh_20_20_io_out_control_0_shift;
	wire [2:0] _mesh_20_20_io_out_id_0;
	wire _mesh_20_20_io_out_last_0;
	wire _mesh_20_20_io_out_valid_0;
	wire [31:0] _mesh_20_19_io_out_a_0;
	wire [31:0] _mesh_20_19_io_out_c_0;
	wire [31:0] _mesh_20_19_io_out_b_0;
	wire _mesh_20_19_io_out_control_0_dataflow;
	wire _mesh_20_19_io_out_control_0_propagate;
	wire [4:0] _mesh_20_19_io_out_control_0_shift;
	wire [2:0] _mesh_20_19_io_out_id_0;
	wire _mesh_20_19_io_out_last_0;
	wire _mesh_20_19_io_out_valid_0;
	wire [31:0] _mesh_20_18_io_out_a_0;
	wire [31:0] _mesh_20_18_io_out_c_0;
	wire [31:0] _mesh_20_18_io_out_b_0;
	wire _mesh_20_18_io_out_control_0_dataflow;
	wire _mesh_20_18_io_out_control_0_propagate;
	wire [4:0] _mesh_20_18_io_out_control_0_shift;
	wire [2:0] _mesh_20_18_io_out_id_0;
	wire _mesh_20_18_io_out_last_0;
	wire _mesh_20_18_io_out_valid_0;
	wire [31:0] _mesh_20_17_io_out_a_0;
	wire [31:0] _mesh_20_17_io_out_c_0;
	wire [31:0] _mesh_20_17_io_out_b_0;
	wire _mesh_20_17_io_out_control_0_dataflow;
	wire _mesh_20_17_io_out_control_0_propagate;
	wire [4:0] _mesh_20_17_io_out_control_0_shift;
	wire [2:0] _mesh_20_17_io_out_id_0;
	wire _mesh_20_17_io_out_last_0;
	wire _mesh_20_17_io_out_valid_0;
	wire [31:0] _mesh_20_16_io_out_a_0;
	wire [31:0] _mesh_20_16_io_out_c_0;
	wire [31:0] _mesh_20_16_io_out_b_0;
	wire _mesh_20_16_io_out_control_0_dataflow;
	wire _mesh_20_16_io_out_control_0_propagate;
	wire [4:0] _mesh_20_16_io_out_control_0_shift;
	wire [2:0] _mesh_20_16_io_out_id_0;
	wire _mesh_20_16_io_out_last_0;
	wire _mesh_20_16_io_out_valid_0;
	wire [31:0] _mesh_20_15_io_out_a_0;
	wire [31:0] _mesh_20_15_io_out_c_0;
	wire [31:0] _mesh_20_15_io_out_b_0;
	wire _mesh_20_15_io_out_control_0_dataflow;
	wire _mesh_20_15_io_out_control_0_propagate;
	wire [4:0] _mesh_20_15_io_out_control_0_shift;
	wire [2:0] _mesh_20_15_io_out_id_0;
	wire _mesh_20_15_io_out_last_0;
	wire _mesh_20_15_io_out_valid_0;
	wire [31:0] _mesh_20_14_io_out_a_0;
	wire [31:0] _mesh_20_14_io_out_c_0;
	wire [31:0] _mesh_20_14_io_out_b_0;
	wire _mesh_20_14_io_out_control_0_dataflow;
	wire _mesh_20_14_io_out_control_0_propagate;
	wire [4:0] _mesh_20_14_io_out_control_0_shift;
	wire [2:0] _mesh_20_14_io_out_id_0;
	wire _mesh_20_14_io_out_last_0;
	wire _mesh_20_14_io_out_valid_0;
	wire [31:0] _mesh_20_13_io_out_a_0;
	wire [31:0] _mesh_20_13_io_out_c_0;
	wire [31:0] _mesh_20_13_io_out_b_0;
	wire _mesh_20_13_io_out_control_0_dataflow;
	wire _mesh_20_13_io_out_control_0_propagate;
	wire [4:0] _mesh_20_13_io_out_control_0_shift;
	wire [2:0] _mesh_20_13_io_out_id_0;
	wire _mesh_20_13_io_out_last_0;
	wire _mesh_20_13_io_out_valid_0;
	wire [31:0] _mesh_20_12_io_out_a_0;
	wire [31:0] _mesh_20_12_io_out_c_0;
	wire [31:0] _mesh_20_12_io_out_b_0;
	wire _mesh_20_12_io_out_control_0_dataflow;
	wire _mesh_20_12_io_out_control_0_propagate;
	wire [4:0] _mesh_20_12_io_out_control_0_shift;
	wire [2:0] _mesh_20_12_io_out_id_0;
	wire _mesh_20_12_io_out_last_0;
	wire _mesh_20_12_io_out_valid_0;
	wire [31:0] _mesh_20_11_io_out_a_0;
	wire [31:0] _mesh_20_11_io_out_c_0;
	wire [31:0] _mesh_20_11_io_out_b_0;
	wire _mesh_20_11_io_out_control_0_dataflow;
	wire _mesh_20_11_io_out_control_0_propagate;
	wire [4:0] _mesh_20_11_io_out_control_0_shift;
	wire [2:0] _mesh_20_11_io_out_id_0;
	wire _mesh_20_11_io_out_last_0;
	wire _mesh_20_11_io_out_valid_0;
	wire [31:0] _mesh_20_10_io_out_a_0;
	wire [31:0] _mesh_20_10_io_out_c_0;
	wire [31:0] _mesh_20_10_io_out_b_0;
	wire _mesh_20_10_io_out_control_0_dataflow;
	wire _mesh_20_10_io_out_control_0_propagate;
	wire [4:0] _mesh_20_10_io_out_control_0_shift;
	wire [2:0] _mesh_20_10_io_out_id_0;
	wire _mesh_20_10_io_out_last_0;
	wire _mesh_20_10_io_out_valid_0;
	wire [31:0] _mesh_20_9_io_out_a_0;
	wire [31:0] _mesh_20_9_io_out_c_0;
	wire [31:0] _mesh_20_9_io_out_b_0;
	wire _mesh_20_9_io_out_control_0_dataflow;
	wire _mesh_20_9_io_out_control_0_propagate;
	wire [4:0] _mesh_20_9_io_out_control_0_shift;
	wire [2:0] _mesh_20_9_io_out_id_0;
	wire _mesh_20_9_io_out_last_0;
	wire _mesh_20_9_io_out_valid_0;
	wire [31:0] _mesh_20_8_io_out_a_0;
	wire [31:0] _mesh_20_8_io_out_c_0;
	wire [31:0] _mesh_20_8_io_out_b_0;
	wire _mesh_20_8_io_out_control_0_dataflow;
	wire _mesh_20_8_io_out_control_0_propagate;
	wire [4:0] _mesh_20_8_io_out_control_0_shift;
	wire [2:0] _mesh_20_8_io_out_id_0;
	wire _mesh_20_8_io_out_last_0;
	wire _mesh_20_8_io_out_valid_0;
	wire [31:0] _mesh_20_7_io_out_a_0;
	wire [31:0] _mesh_20_7_io_out_c_0;
	wire [31:0] _mesh_20_7_io_out_b_0;
	wire _mesh_20_7_io_out_control_0_dataflow;
	wire _mesh_20_7_io_out_control_0_propagate;
	wire [4:0] _mesh_20_7_io_out_control_0_shift;
	wire [2:0] _mesh_20_7_io_out_id_0;
	wire _mesh_20_7_io_out_last_0;
	wire _mesh_20_7_io_out_valid_0;
	wire [31:0] _mesh_20_6_io_out_a_0;
	wire [31:0] _mesh_20_6_io_out_c_0;
	wire [31:0] _mesh_20_6_io_out_b_0;
	wire _mesh_20_6_io_out_control_0_dataflow;
	wire _mesh_20_6_io_out_control_0_propagate;
	wire [4:0] _mesh_20_6_io_out_control_0_shift;
	wire [2:0] _mesh_20_6_io_out_id_0;
	wire _mesh_20_6_io_out_last_0;
	wire _mesh_20_6_io_out_valid_0;
	wire [31:0] _mesh_20_5_io_out_a_0;
	wire [31:0] _mesh_20_5_io_out_c_0;
	wire [31:0] _mesh_20_5_io_out_b_0;
	wire _mesh_20_5_io_out_control_0_dataflow;
	wire _mesh_20_5_io_out_control_0_propagate;
	wire [4:0] _mesh_20_5_io_out_control_0_shift;
	wire [2:0] _mesh_20_5_io_out_id_0;
	wire _mesh_20_5_io_out_last_0;
	wire _mesh_20_5_io_out_valid_0;
	wire [31:0] _mesh_20_4_io_out_a_0;
	wire [31:0] _mesh_20_4_io_out_c_0;
	wire [31:0] _mesh_20_4_io_out_b_0;
	wire _mesh_20_4_io_out_control_0_dataflow;
	wire _mesh_20_4_io_out_control_0_propagate;
	wire [4:0] _mesh_20_4_io_out_control_0_shift;
	wire [2:0] _mesh_20_4_io_out_id_0;
	wire _mesh_20_4_io_out_last_0;
	wire _mesh_20_4_io_out_valid_0;
	wire [31:0] _mesh_20_3_io_out_a_0;
	wire [31:0] _mesh_20_3_io_out_c_0;
	wire [31:0] _mesh_20_3_io_out_b_0;
	wire _mesh_20_3_io_out_control_0_dataflow;
	wire _mesh_20_3_io_out_control_0_propagate;
	wire [4:0] _mesh_20_3_io_out_control_0_shift;
	wire [2:0] _mesh_20_3_io_out_id_0;
	wire _mesh_20_3_io_out_last_0;
	wire _mesh_20_3_io_out_valid_0;
	wire [31:0] _mesh_20_2_io_out_a_0;
	wire [31:0] _mesh_20_2_io_out_c_0;
	wire [31:0] _mesh_20_2_io_out_b_0;
	wire _mesh_20_2_io_out_control_0_dataflow;
	wire _mesh_20_2_io_out_control_0_propagate;
	wire [4:0] _mesh_20_2_io_out_control_0_shift;
	wire [2:0] _mesh_20_2_io_out_id_0;
	wire _mesh_20_2_io_out_last_0;
	wire _mesh_20_2_io_out_valid_0;
	wire [31:0] _mesh_20_1_io_out_a_0;
	wire [31:0] _mesh_20_1_io_out_c_0;
	wire [31:0] _mesh_20_1_io_out_b_0;
	wire _mesh_20_1_io_out_control_0_dataflow;
	wire _mesh_20_1_io_out_control_0_propagate;
	wire [4:0] _mesh_20_1_io_out_control_0_shift;
	wire [2:0] _mesh_20_1_io_out_id_0;
	wire _mesh_20_1_io_out_last_0;
	wire _mesh_20_1_io_out_valid_0;
	wire [31:0] _mesh_20_0_io_out_a_0;
	wire [31:0] _mesh_20_0_io_out_c_0;
	wire [31:0] _mesh_20_0_io_out_b_0;
	wire _mesh_20_0_io_out_control_0_dataflow;
	wire _mesh_20_0_io_out_control_0_propagate;
	wire [4:0] _mesh_20_0_io_out_control_0_shift;
	wire [2:0] _mesh_20_0_io_out_id_0;
	wire _mesh_20_0_io_out_last_0;
	wire _mesh_20_0_io_out_valid_0;
	wire [31:0] _mesh_19_31_io_out_a_0;
	wire [31:0] _mesh_19_31_io_out_c_0;
	wire [31:0] _mesh_19_31_io_out_b_0;
	wire _mesh_19_31_io_out_control_0_dataflow;
	wire _mesh_19_31_io_out_control_0_propagate;
	wire [4:0] _mesh_19_31_io_out_control_0_shift;
	wire [2:0] _mesh_19_31_io_out_id_0;
	wire _mesh_19_31_io_out_last_0;
	wire _mesh_19_31_io_out_valid_0;
	wire [31:0] _mesh_19_30_io_out_a_0;
	wire [31:0] _mesh_19_30_io_out_c_0;
	wire [31:0] _mesh_19_30_io_out_b_0;
	wire _mesh_19_30_io_out_control_0_dataflow;
	wire _mesh_19_30_io_out_control_0_propagate;
	wire [4:0] _mesh_19_30_io_out_control_0_shift;
	wire [2:0] _mesh_19_30_io_out_id_0;
	wire _mesh_19_30_io_out_last_0;
	wire _mesh_19_30_io_out_valid_0;
	wire [31:0] _mesh_19_29_io_out_a_0;
	wire [31:0] _mesh_19_29_io_out_c_0;
	wire [31:0] _mesh_19_29_io_out_b_0;
	wire _mesh_19_29_io_out_control_0_dataflow;
	wire _mesh_19_29_io_out_control_0_propagate;
	wire [4:0] _mesh_19_29_io_out_control_0_shift;
	wire [2:0] _mesh_19_29_io_out_id_0;
	wire _mesh_19_29_io_out_last_0;
	wire _mesh_19_29_io_out_valid_0;
	wire [31:0] _mesh_19_28_io_out_a_0;
	wire [31:0] _mesh_19_28_io_out_c_0;
	wire [31:0] _mesh_19_28_io_out_b_0;
	wire _mesh_19_28_io_out_control_0_dataflow;
	wire _mesh_19_28_io_out_control_0_propagate;
	wire [4:0] _mesh_19_28_io_out_control_0_shift;
	wire [2:0] _mesh_19_28_io_out_id_0;
	wire _mesh_19_28_io_out_last_0;
	wire _mesh_19_28_io_out_valid_0;
	wire [31:0] _mesh_19_27_io_out_a_0;
	wire [31:0] _mesh_19_27_io_out_c_0;
	wire [31:0] _mesh_19_27_io_out_b_0;
	wire _mesh_19_27_io_out_control_0_dataflow;
	wire _mesh_19_27_io_out_control_0_propagate;
	wire [4:0] _mesh_19_27_io_out_control_0_shift;
	wire [2:0] _mesh_19_27_io_out_id_0;
	wire _mesh_19_27_io_out_last_0;
	wire _mesh_19_27_io_out_valid_0;
	wire [31:0] _mesh_19_26_io_out_a_0;
	wire [31:0] _mesh_19_26_io_out_c_0;
	wire [31:0] _mesh_19_26_io_out_b_0;
	wire _mesh_19_26_io_out_control_0_dataflow;
	wire _mesh_19_26_io_out_control_0_propagate;
	wire [4:0] _mesh_19_26_io_out_control_0_shift;
	wire [2:0] _mesh_19_26_io_out_id_0;
	wire _mesh_19_26_io_out_last_0;
	wire _mesh_19_26_io_out_valid_0;
	wire [31:0] _mesh_19_25_io_out_a_0;
	wire [31:0] _mesh_19_25_io_out_c_0;
	wire [31:0] _mesh_19_25_io_out_b_0;
	wire _mesh_19_25_io_out_control_0_dataflow;
	wire _mesh_19_25_io_out_control_0_propagate;
	wire [4:0] _mesh_19_25_io_out_control_0_shift;
	wire [2:0] _mesh_19_25_io_out_id_0;
	wire _mesh_19_25_io_out_last_0;
	wire _mesh_19_25_io_out_valid_0;
	wire [31:0] _mesh_19_24_io_out_a_0;
	wire [31:0] _mesh_19_24_io_out_c_0;
	wire [31:0] _mesh_19_24_io_out_b_0;
	wire _mesh_19_24_io_out_control_0_dataflow;
	wire _mesh_19_24_io_out_control_0_propagate;
	wire [4:0] _mesh_19_24_io_out_control_0_shift;
	wire [2:0] _mesh_19_24_io_out_id_0;
	wire _mesh_19_24_io_out_last_0;
	wire _mesh_19_24_io_out_valid_0;
	wire [31:0] _mesh_19_23_io_out_a_0;
	wire [31:0] _mesh_19_23_io_out_c_0;
	wire [31:0] _mesh_19_23_io_out_b_0;
	wire _mesh_19_23_io_out_control_0_dataflow;
	wire _mesh_19_23_io_out_control_0_propagate;
	wire [4:0] _mesh_19_23_io_out_control_0_shift;
	wire [2:0] _mesh_19_23_io_out_id_0;
	wire _mesh_19_23_io_out_last_0;
	wire _mesh_19_23_io_out_valid_0;
	wire [31:0] _mesh_19_22_io_out_a_0;
	wire [31:0] _mesh_19_22_io_out_c_0;
	wire [31:0] _mesh_19_22_io_out_b_0;
	wire _mesh_19_22_io_out_control_0_dataflow;
	wire _mesh_19_22_io_out_control_0_propagate;
	wire [4:0] _mesh_19_22_io_out_control_0_shift;
	wire [2:0] _mesh_19_22_io_out_id_0;
	wire _mesh_19_22_io_out_last_0;
	wire _mesh_19_22_io_out_valid_0;
	wire [31:0] _mesh_19_21_io_out_a_0;
	wire [31:0] _mesh_19_21_io_out_c_0;
	wire [31:0] _mesh_19_21_io_out_b_0;
	wire _mesh_19_21_io_out_control_0_dataflow;
	wire _mesh_19_21_io_out_control_0_propagate;
	wire [4:0] _mesh_19_21_io_out_control_0_shift;
	wire [2:0] _mesh_19_21_io_out_id_0;
	wire _mesh_19_21_io_out_last_0;
	wire _mesh_19_21_io_out_valid_0;
	wire [31:0] _mesh_19_20_io_out_a_0;
	wire [31:0] _mesh_19_20_io_out_c_0;
	wire [31:0] _mesh_19_20_io_out_b_0;
	wire _mesh_19_20_io_out_control_0_dataflow;
	wire _mesh_19_20_io_out_control_0_propagate;
	wire [4:0] _mesh_19_20_io_out_control_0_shift;
	wire [2:0] _mesh_19_20_io_out_id_0;
	wire _mesh_19_20_io_out_last_0;
	wire _mesh_19_20_io_out_valid_0;
	wire [31:0] _mesh_19_19_io_out_a_0;
	wire [31:0] _mesh_19_19_io_out_c_0;
	wire [31:0] _mesh_19_19_io_out_b_0;
	wire _mesh_19_19_io_out_control_0_dataflow;
	wire _mesh_19_19_io_out_control_0_propagate;
	wire [4:0] _mesh_19_19_io_out_control_0_shift;
	wire [2:0] _mesh_19_19_io_out_id_0;
	wire _mesh_19_19_io_out_last_0;
	wire _mesh_19_19_io_out_valid_0;
	wire [31:0] _mesh_19_18_io_out_a_0;
	wire [31:0] _mesh_19_18_io_out_c_0;
	wire [31:0] _mesh_19_18_io_out_b_0;
	wire _mesh_19_18_io_out_control_0_dataflow;
	wire _mesh_19_18_io_out_control_0_propagate;
	wire [4:0] _mesh_19_18_io_out_control_0_shift;
	wire [2:0] _mesh_19_18_io_out_id_0;
	wire _mesh_19_18_io_out_last_0;
	wire _mesh_19_18_io_out_valid_0;
	wire [31:0] _mesh_19_17_io_out_a_0;
	wire [31:0] _mesh_19_17_io_out_c_0;
	wire [31:0] _mesh_19_17_io_out_b_0;
	wire _mesh_19_17_io_out_control_0_dataflow;
	wire _mesh_19_17_io_out_control_0_propagate;
	wire [4:0] _mesh_19_17_io_out_control_0_shift;
	wire [2:0] _mesh_19_17_io_out_id_0;
	wire _mesh_19_17_io_out_last_0;
	wire _mesh_19_17_io_out_valid_0;
	wire [31:0] _mesh_19_16_io_out_a_0;
	wire [31:0] _mesh_19_16_io_out_c_0;
	wire [31:0] _mesh_19_16_io_out_b_0;
	wire _mesh_19_16_io_out_control_0_dataflow;
	wire _mesh_19_16_io_out_control_0_propagate;
	wire [4:0] _mesh_19_16_io_out_control_0_shift;
	wire [2:0] _mesh_19_16_io_out_id_0;
	wire _mesh_19_16_io_out_last_0;
	wire _mesh_19_16_io_out_valid_0;
	wire [31:0] _mesh_19_15_io_out_a_0;
	wire [31:0] _mesh_19_15_io_out_c_0;
	wire [31:0] _mesh_19_15_io_out_b_0;
	wire _mesh_19_15_io_out_control_0_dataflow;
	wire _mesh_19_15_io_out_control_0_propagate;
	wire [4:0] _mesh_19_15_io_out_control_0_shift;
	wire [2:0] _mesh_19_15_io_out_id_0;
	wire _mesh_19_15_io_out_last_0;
	wire _mesh_19_15_io_out_valid_0;
	wire [31:0] _mesh_19_14_io_out_a_0;
	wire [31:0] _mesh_19_14_io_out_c_0;
	wire [31:0] _mesh_19_14_io_out_b_0;
	wire _mesh_19_14_io_out_control_0_dataflow;
	wire _mesh_19_14_io_out_control_0_propagate;
	wire [4:0] _mesh_19_14_io_out_control_0_shift;
	wire [2:0] _mesh_19_14_io_out_id_0;
	wire _mesh_19_14_io_out_last_0;
	wire _mesh_19_14_io_out_valid_0;
	wire [31:0] _mesh_19_13_io_out_a_0;
	wire [31:0] _mesh_19_13_io_out_c_0;
	wire [31:0] _mesh_19_13_io_out_b_0;
	wire _mesh_19_13_io_out_control_0_dataflow;
	wire _mesh_19_13_io_out_control_0_propagate;
	wire [4:0] _mesh_19_13_io_out_control_0_shift;
	wire [2:0] _mesh_19_13_io_out_id_0;
	wire _mesh_19_13_io_out_last_0;
	wire _mesh_19_13_io_out_valid_0;
	wire [31:0] _mesh_19_12_io_out_a_0;
	wire [31:0] _mesh_19_12_io_out_c_0;
	wire [31:0] _mesh_19_12_io_out_b_0;
	wire _mesh_19_12_io_out_control_0_dataflow;
	wire _mesh_19_12_io_out_control_0_propagate;
	wire [4:0] _mesh_19_12_io_out_control_0_shift;
	wire [2:0] _mesh_19_12_io_out_id_0;
	wire _mesh_19_12_io_out_last_0;
	wire _mesh_19_12_io_out_valid_0;
	wire [31:0] _mesh_19_11_io_out_a_0;
	wire [31:0] _mesh_19_11_io_out_c_0;
	wire [31:0] _mesh_19_11_io_out_b_0;
	wire _mesh_19_11_io_out_control_0_dataflow;
	wire _mesh_19_11_io_out_control_0_propagate;
	wire [4:0] _mesh_19_11_io_out_control_0_shift;
	wire [2:0] _mesh_19_11_io_out_id_0;
	wire _mesh_19_11_io_out_last_0;
	wire _mesh_19_11_io_out_valid_0;
	wire [31:0] _mesh_19_10_io_out_a_0;
	wire [31:0] _mesh_19_10_io_out_c_0;
	wire [31:0] _mesh_19_10_io_out_b_0;
	wire _mesh_19_10_io_out_control_0_dataflow;
	wire _mesh_19_10_io_out_control_0_propagate;
	wire [4:0] _mesh_19_10_io_out_control_0_shift;
	wire [2:0] _mesh_19_10_io_out_id_0;
	wire _mesh_19_10_io_out_last_0;
	wire _mesh_19_10_io_out_valid_0;
	wire [31:0] _mesh_19_9_io_out_a_0;
	wire [31:0] _mesh_19_9_io_out_c_0;
	wire [31:0] _mesh_19_9_io_out_b_0;
	wire _mesh_19_9_io_out_control_0_dataflow;
	wire _mesh_19_9_io_out_control_0_propagate;
	wire [4:0] _mesh_19_9_io_out_control_0_shift;
	wire [2:0] _mesh_19_9_io_out_id_0;
	wire _mesh_19_9_io_out_last_0;
	wire _mesh_19_9_io_out_valid_0;
	wire [31:0] _mesh_19_8_io_out_a_0;
	wire [31:0] _mesh_19_8_io_out_c_0;
	wire [31:0] _mesh_19_8_io_out_b_0;
	wire _mesh_19_8_io_out_control_0_dataflow;
	wire _mesh_19_8_io_out_control_0_propagate;
	wire [4:0] _mesh_19_8_io_out_control_0_shift;
	wire [2:0] _mesh_19_8_io_out_id_0;
	wire _mesh_19_8_io_out_last_0;
	wire _mesh_19_8_io_out_valid_0;
	wire [31:0] _mesh_19_7_io_out_a_0;
	wire [31:0] _mesh_19_7_io_out_c_0;
	wire [31:0] _mesh_19_7_io_out_b_0;
	wire _mesh_19_7_io_out_control_0_dataflow;
	wire _mesh_19_7_io_out_control_0_propagate;
	wire [4:0] _mesh_19_7_io_out_control_0_shift;
	wire [2:0] _mesh_19_7_io_out_id_0;
	wire _mesh_19_7_io_out_last_0;
	wire _mesh_19_7_io_out_valid_0;
	wire [31:0] _mesh_19_6_io_out_a_0;
	wire [31:0] _mesh_19_6_io_out_c_0;
	wire [31:0] _mesh_19_6_io_out_b_0;
	wire _mesh_19_6_io_out_control_0_dataflow;
	wire _mesh_19_6_io_out_control_0_propagate;
	wire [4:0] _mesh_19_6_io_out_control_0_shift;
	wire [2:0] _mesh_19_6_io_out_id_0;
	wire _mesh_19_6_io_out_last_0;
	wire _mesh_19_6_io_out_valid_0;
	wire [31:0] _mesh_19_5_io_out_a_0;
	wire [31:0] _mesh_19_5_io_out_c_0;
	wire [31:0] _mesh_19_5_io_out_b_0;
	wire _mesh_19_5_io_out_control_0_dataflow;
	wire _mesh_19_5_io_out_control_0_propagate;
	wire [4:0] _mesh_19_5_io_out_control_0_shift;
	wire [2:0] _mesh_19_5_io_out_id_0;
	wire _mesh_19_5_io_out_last_0;
	wire _mesh_19_5_io_out_valid_0;
	wire [31:0] _mesh_19_4_io_out_a_0;
	wire [31:0] _mesh_19_4_io_out_c_0;
	wire [31:0] _mesh_19_4_io_out_b_0;
	wire _mesh_19_4_io_out_control_0_dataflow;
	wire _mesh_19_4_io_out_control_0_propagate;
	wire [4:0] _mesh_19_4_io_out_control_0_shift;
	wire [2:0] _mesh_19_4_io_out_id_0;
	wire _mesh_19_4_io_out_last_0;
	wire _mesh_19_4_io_out_valid_0;
	wire [31:0] _mesh_19_3_io_out_a_0;
	wire [31:0] _mesh_19_3_io_out_c_0;
	wire [31:0] _mesh_19_3_io_out_b_0;
	wire _mesh_19_3_io_out_control_0_dataflow;
	wire _mesh_19_3_io_out_control_0_propagate;
	wire [4:0] _mesh_19_3_io_out_control_0_shift;
	wire [2:0] _mesh_19_3_io_out_id_0;
	wire _mesh_19_3_io_out_last_0;
	wire _mesh_19_3_io_out_valid_0;
	wire [31:0] _mesh_19_2_io_out_a_0;
	wire [31:0] _mesh_19_2_io_out_c_0;
	wire [31:0] _mesh_19_2_io_out_b_0;
	wire _mesh_19_2_io_out_control_0_dataflow;
	wire _mesh_19_2_io_out_control_0_propagate;
	wire [4:0] _mesh_19_2_io_out_control_0_shift;
	wire [2:0] _mesh_19_2_io_out_id_0;
	wire _mesh_19_2_io_out_last_0;
	wire _mesh_19_2_io_out_valid_0;
	wire [31:0] _mesh_19_1_io_out_a_0;
	wire [31:0] _mesh_19_1_io_out_c_0;
	wire [31:0] _mesh_19_1_io_out_b_0;
	wire _mesh_19_1_io_out_control_0_dataflow;
	wire _mesh_19_1_io_out_control_0_propagate;
	wire [4:0] _mesh_19_1_io_out_control_0_shift;
	wire [2:0] _mesh_19_1_io_out_id_0;
	wire _mesh_19_1_io_out_last_0;
	wire _mesh_19_1_io_out_valid_0;
	wire [31:0] _mesh_19_0_io_out_a_0;
	wire [31:0] _mesh_19_0_io_out_c_0;
	wire [31:0] _mesh_19_0_io_out_b_0;
	wire _mesh_19_0_io_out_control_0_dataflow;
	wire _mesh_19_0_io_out_control_0_propagate;
	wire [4:0] _mesh_19_0_io_out_control_0_shift;
	wire [2:0] _mesh_19_0_io_out_id_0;
	wire _mesh_19_0_io_out_last_0;
	wire _mesh_19_0_io_out_valid_0;
	wire [31:0] _mesh_18_31_io_out_a_0;
	wire [31:0] _mesh_18_31_io_out_c_0;
	wire [31:0] _mesh_18_31_io_out_b_0;
	wire _mesh_18_31_io_out_control_0_dataflow;
	wire _mesh_18_31_io_out_control_0_propagate;
	wire [4:0] _mesh_18_31_io_out_control_0_shift;
	wire [2:0] _mesh_18_31_io_out_id_0;
	wire _mesh_18_31_io_out_last_0;
	wire _mesh_18_31_io_out_valid_0;
	wire [31:0] _mesh_18_30_io_out_a_0;
	wire [31:0] _mesh_18_30_io_out_c_0;
	wire [31:0] _mesh_18_30_io_out_b_0;
	wire _mesh_18_30_io_out_control_0_dataflow;
	wire _mesh_18_30_io_out_control_0_propagate;
	wire [4:0] _mesh_18_30_io_out_control_0_shift;
	wire [2:0] _mesh_18_30_io_out_id_0;
	wire _mesh_18_30_io_out_last_0;
	wire _mesh_18_30_io_out_valid_0;
	wire [31:0] _mesh_18_29_io_out_a_0;
	wire [31:0] _mesh_18_29_io_out_c_0;
	wire [31:0] _mesh_18_29_io_out_b_0;
	wire _mesh_18_29_io_out_control_0_dataflow;
	wire _mesh_18_29_io_out_control_0_propagate;
	wire [4:0] _mesh_18_29_io_out_control_0_shift;
	wire [2:0] _mesh_18_29_io_out_id_0;
	wire _mesh_18_29_io_out_last_0;
	wire _mesh_18_29_io_out_valid_0;
	wire [31:0] _mesh_18_28_io_out_a_0;
	wire [31:0] _mesh_18_28_io_out_c_0;
	wire [31:0] _mesh_18_28_io_out_b_0;
	wire _mesh_18_28_io_out_control_0_dataflow;
	wire _mesh_18_28_io_out_control_0_propagate;
	wire [4:0] _mesh_18_28_io_out_control_0_shift;
	wire [2:0] _mesh_18_28_io_out_id_0;
	wire _mesh_18_28_io_out_last_0;
	wire _mesh_18_28_io_out_valid_0;
	wire [31:0] _mesh_18_27_io_out_a_0;
	wire [31:0] _mesh_18_27_io_out_c_0;
	wire [31:0] _mesh_18_27_io_out_b_0;
	wire _mesh_18_27_io_out_control_0_dataflow;
	wire _mesh_18_27_io_out_control_0_propagate;
	wire [4:0] _mesh_18_27_io_out_control_0_shift;
	wire [2:0] _mesh_18_27_io_out_id_0;
	wire _mesh_18_27_io_out_last_0;
	wire _mesh_18_27_io_out_valid_0;
	wire [31:0] _mesh_18_26_io_out_a_0;
	wire [31:0] _mesh_18_26_io_out_c_0;
	wire [31:0] _mesh_18_26_io_out_b_0;
	wire _mesh_18_26_io_out_control_0_dataflow;
	wire _mesh_18_26_io_out_control_0_propagate;
	wire [4:0] _mesh_18_26_io_out_control_0_shift;
	wire [2:0] _mesh_18_26_io_out_id_0;
	wire _mesh_18_26_io_out_last_0;
	wire _mesh_18_26_io_out_valid_0;
	wire [31:0] _mesh_18_25_io_out_a_0;
	wire [31:0] _mesh_18_25_io_out_c_0;
	wire [31:0] _mesh_18_25_io_out_b_0;
	wire _mesh_18_25_io_out_control_0_dataflow;
	wire _mesh_18_25_io_out_control_0_propagate;
	wire [4:0] _mesh_18_25_io_out_control_0_shift;
	wire [2:0] _mesh_18_25_io_out_id_0;
	wire _mesh_18_25_io_out_last_0;
	wire _mesh_18_25_io_out_valid_0;
	wire [31:0] _mesh_18_24_io_out_a_0;
	wire [31:0] _mesh_18_24_io_out_c_0;
	wire [31:0] _mesh_18_24_io_out_b_0;
	wire _mesh_18_24_io_out_control_0_dataflow;
	wire _mesh_18_24_io_out_control_0_propagate;
	wire [4:0] _mesh_18_24_io_out_control_0_shift;
	wire [2:0] _mesh_18_24_io_out_id_0;
	wire _mesh_18_24_io_out_last_0;
	wire _mesh_18_24_io_out_valid_0;
	wire [31:0] _mesh_18_23_io_out_a_0;
	wire [31:0] _mesh_18_23_io_out_c_0;
	wire [31:0] _mesh_18_23_io_out_b_0;
	wire _mesh_18_23_io_out_control_0_dataflow;
	wire _mesh_18_23_io_out_control_0_propagate;
	wire [4:0] _mesh_18_23_io_out_control_0_shift;
	wire [2:0] _mesh_18_23_io_out_id_0;
	wire _mesh_18_23_io_out_last_0;
	wire _mesh_18_23_io_out_valid_0;
	wire [31:0] _mesh_18_22_io_out_a_0;
	wire [31:0] _mesh_18_22_io_out_c_0;
	wire [31:0] _mesh_18_22_io_out_b_0;
	wire _mesh_18_22_io_out_control_0_dataflow;
	wire _mesh_18_22_io_out_control_0_propagate;
	wire [4:0] _mesh_18_22_io_out_control_0_shift;
	wire [2:0] _mesh_18_22_io_out_id_0;
	wire _mesh_18_22_io_out_last_0;
	wire _mesh_18_22_io_out_valid_0;
	wire [31:0] _mesh_18_21_io_out_a_0;
	wire [31:0] _mesh_18_21_io_out_c_0;
	wire [31:0] _mesh_18_21_io_out_b_0;
	wire _mesh_18_21_io_out_control_0_dataflow;
	wire _mesh_18_21_io_out_control_0_propagate;
	wire [4:0] _mesh_18_21_io_out_control_0_shift;
	wire [2:0] _mesh_18_21_io_out_id_0;
	wire _mesh_18_21_io_out_last_0;
	wire _mesh_18_21_io_out_valid_0;
	wire [31:0] _mesh_18_20_io_out_a_0;
	wire [31:0] _mesh_18_20_io_out_c_0;
	wire [31:0] _mesh_18_20_io_out_b_0;
	wire _mesh_18_20_io_out_control_0_dataflow;
	wire _mesh_18_20_io_out_control_0_propagate;
	wire [4:0] _mesh_18_20_io_out_control_0_shift;
	wire [2:0] _mesh_18_20_io_out_id_0;
	wire _mesh_18_20_io_out_last_0;
	wire _mesh_18_20_io_out_valid_0;
	wire [31:0] _mesh_18_19_io_out_a_0;
	wire [31:0] _mesh_18_19_io_out_c_0;
	wire [31:0] _mesh_18_19_io_out_b_0;
	wire _mesh_18_19_io_out_control_0_dataflow;
	wire _mesh_18_19_io_out_control_0_propagate;
	wire [4:0] _mesh_18_19_io_out_control_0_shift;
	wire [2:0] _mesh_18_19_io_out_id_0;
	wire _mesh_18_19_io_out_last_0;
	wire _mesh_18_19_io_out_valid_0;
	wire [31:0] _mesh_18_18_io_out_a_0;
	wire [31:0] _mesh_18_18_io_out_c_0;
	wire [31:0] _mesh_18_18_io_out_b_0;
	wire _mesh_18_18_io_out_control_0_dataflow;
	wire _mesh_18_18_io_out_control_0_propagate;
	wire [4:0] _mesh_18_18_io_out_control_0_shift;
	wire [2:0] _mesh_18_18_io_out_id_0;
	wire _mesh_18_18_io_out_last_0;
	wire _mesh_18_18_io_out_valid_0;
	wire [31:0] _mesh_18_17_io_out_a_0;
	wire [31:0] _mesh_18_17_io_out_c_0;
	wire [31:0] _mesh_18_17_io_out_b_0;
	wire _mesh_18_17_io_out_control_0_dataflow;
	wire _mesh_18_17_io_out_control_0_propagate;
	wire [4:0] _mesh_18_17_io_out_control_0_shift;
	wire [2:0] _mesh_18_17_io_out_id_0;
	wire _mesh_18_17_io_out_last_0;
	wire _mesh_18_17_io_out_valid_0;
	wire [31:0] _mesh_18_16_io_out_a_0;
	wire [31:0] _mesh_18_16_io_out_c_0;
	wire [31:0] _mesh_18_16_io_out_b_0;
	wire _mesh_18_16_io_out_control_0_dataflow;
	wire _mesh_18_16_io_out_control_0_propagate;
	wire [4:0] _mesh_18_16_io_out_control_0_shift;
	wire [2:0] _mesh_18_16_io_out_id_0;
	wire _mesh_18_16_io_out_last_0;
	wire _mesh_18_16_io_out_valid_0;
	wire [31:0] _mesh_18_15_io_out_a_0;
	wire [31:0] _mesh_18_15_io_out_c_0;
	wire [31:0] _mesh_18_15_io_out_b_0;
	wire _mesh_18_15_io_out_control_0_dataflow;
	wire _mesh_18_15_io_out_control_0_propagate;
	wire [4:0] _mesh_18_15_io_out_control_0_shift;
	wire [2:0] _mesh_18_15_io_out_id_0;
	wire _mesh_18_15_io_out_last_0;
	wire _mesh_18_15_io_out_valid_0;
	wire [31:0] _mesh_18_14_io_out_a_0;
	wire [31:0] _mesh_18_14_io_out_c_0;
	wire [31:0] _mesh_18_14_io_out_b_0;
	wire _mesh_18_14_io_out_control_0_dataflow;
	wire _mesh_18_14_io_out_control_0_propagate;
	wire [4:0] _mesh_18_14_io_out_control_0_shift;
	wire [2:0] _mesh_18_14_io_out_id_0;
	wire _mesh_18_14_io_out_last_0;
	wire _mesh_18_14_io_out_valid_0;
	wire [31:0] _mesh_18_13_io_out_a_0;
	wire [31:0] _mesh_18_13_io_out_c_0;
	wire [31:0] _mesh_18_13_io_out_b_0;
	wire _mesh_18_13_io_out_control_0_dataflow;
	wire _mesh_18_13_io_out_control_0_propagate;
	wire [4:0] _mesh_18_13_io_out_control_0_shift;
	wire [2:0] _mesh_18_13_io_out_id_0;
	wire _mesh_18_13_io_out_last_0;
	wire _mesh_18_13_io_out_valid_0;
	wire [31:0] _mesh_18_12_io_out_a_0;
	wire [31:0] _mesh_18_12_io_out_c_0;
	wire [31:0] _mesh_18_12_io_out_b_0;
	wire _mesh_18_12_io_out_control_0_dataflow;
	wire _mesh_18_12_io_out_control_0_propagate;
	wire [4:0] _mesh_18_12_io_out_control_0_shift;
	wire [2:0] _mesh_18_12_io_out_id_0;
	wire _mesh_18_12_io_out_last_0;
	wire _mesh_18_12_io_out_valid_0;
	wire [31:0] _mesh_18_11_io_out_a_0;
	wire [31:0] _mesh_18_11_io_out_c_0;
	wire [31:0] _mesh_18_11_io_out_b_0;
	wire _mesh_18_11_io_out_control_0_dataflow;
	wire _mesh_18_11_io_out_control_0_propagate;
	wire [4:0] _mesh_18_11_io_out_control_0_shift;
	wire [2:0] _mesh_18_11_io_out_id_0;
	wire _mesh_18_11_io_out_last_0;
	wire _mesh_18_11_io_out_valid_0;
	wire [31:0] _mesh_18_10_io_out_a_0;
	wire [31:0] _mesh_18_10_io_out_c_0;
	wire [31:0] _mesh_18_10_io_out_b_0;
	wire _mesh_18_10_io_out_control_0_dataflow;
	wire _mesh_18_10_io_out_control_0_propagate;
	wire [4:0] _mesh_18_10_io_out_control_0_shift;
	wire [2:0] _mesh_18_10_io_out_id_0;
	wire _mesh_18_10_io_out_last_0;
	wire _mesh_18_10_io_out_valid_0;
	wire [31:0] _mesh_18_9_io_out_a_0;
	wire [31:0] _mesh_18_9_io_out_c_0;
	wire [31:0] _mesh_18_9_io_out_b_0;
	wire _mesh_18_9_io_out_control_0_dataflow;
	wire _mesh_18_9_io_out_control_0_propagate;
	wire [4:0] _mesh_18_9_io_out_control_0_shift;
	wire [2:0] _mesh_18_9_io_out_id_0;
	wire _mesh_18_9_io_out_last_0;
	wire _mesh_18_9_io_out_valid_0;
	wire [31:0] _mesh_18_8_io_out_a_0;
	wire [31:0] _mesh_18_8_io_out_c_0;
	wire [31:0] _mesh_18_8_io_out_b_0;
	wire _mesh_18_8_io_out_control_0_dataflow;
	wire _mesh_18_8_io_out_control_0_propagate;
	wire [4:0] _mesh_18_8_io_out_control_0_shift;
	wire [2:0] _mesh_18_8_io_out_id_0;
	wire _mesh_18_8_io_out_last_0;
	wire _mesh_18_8_io_out_valid_0;
	wire [31:0] _mesh_18_7_io_out_a_0;
	wire [31:0] _mesh_18_7_io_out_c_0;
	wire [31:0] _mesh_18_7_io_out_b_0;
	wire _mesh_18_7_io_out_control_0_dataflow;
	wire _mesh_18_7_io_out_control_0_propagate;
	wire [4:0] _mesh_18_7_io_out_control_0_shift;
	wire [2:0] _mesh_18_7_io_out_id_0;
	wire _mesh_18_7_io_out_last_0;
	wire _mesh_18_7_io_out_valid_0;
	wire [31:0] _mesh_18_6_io_out_a_0;
	wire [31:0] _mesh_18_6_io_out_c_0;
	wire [31:0] _mesh_18_6_io_out_b_0;
	wire _mesh_18_6_io_out_control_0_dataflow;
	wire _mesh_18_6_io_out_control_0_propagate;
	wire [4:0] _mesh_18_6_io_out_control_0_shift;
	wire [2:0] _mesh_18_6_io_out_id_0;
	wire _mesh_18_6_io_out_last_0;
	wire _mesh_18_6_io_out_valid_0;
	wire [31:0] _mesh_18_5_io_out_a_0;
	wire [31:0] _mesh_18_5_io_out_c_0;
	wire [31:0] _mesh_18_5_io_out_b_0;
	wire _mesh_18_5_io_out_control_0_dataflow;
	wire _mesh_18_5_io_out_control_0_propagate;
	wire [4:0] _mesh_18_5_io_out_control_0_shift;
	wire [2:0] _mesh_18_5_io_out_id_0;
	wire _mesh_18_5_io_out_last_0;
	wire _mesh_18_5_io_out_valid_0;
	wire [31:0] _mesh_18_4_io_out_a_0;
	wire [31:0] _mesh_18_4_io_out_c_0;
	wire [31:0] _mesh_18_4_io_out_b_0;
	wire _mesh_18_4_io_out_control_0_dataflow;
	wire _mesh_18_4_io_out_control_0_propagate;
	wire [4:0] _mesh_18_4_io_out_control_0_shift;
	wire [2:0] _mesh_18_4_io_out_id_0;
	wire _mesh_18_4_io_out_last_0;
	wire _mesh_18_4_io_out_valid_0;
	wire [31:0] _mesh_18_3_io_out_a_0;
	wire [31:0] _mesh_18_3_io_out_c_0;
	wire [31:0] _mesh_18_3_io_out_b_0;
	wire _mesh_18_3_io_out_control_0_dataflow;
	wire _mesh_18_3_io_out_control_0_propagate;
	wire [4:0] _mesh_18_3_io_out_control_0_shift;
	wire [2:0] _mesh_18_3_io_out_id_0;
	wire _mesh_18_3_io_out_last_0;
	wire _mesh_18_3_io_out_valid_0;
	wire [31:0] _mesh_18_2_io_out_a_0;
	wire [31:0] _mesh_18_2_io_out_c_0;
	wire [31:0] _mesh_18_2_io_out_b_0;
	wire _mesh_18_2_io_out_control_0_dataflow;
	wire _mesh_18_2_io_out_control_0_propagate;
	wire [4:0] _mesh_18_2_io_out_control_0_shift;
	wire [2:0] _mesh_18_2_io_out_id_0;
	wire _mesh_18_2_io_out_last_0;
	wire _mesh_18_2_io_out_valid_0;
	wire [31:0] _mesh_18_1_io_out_a_0;
	wire [31:0] _mesh_18_1_io_out_c_0;
	wire [31:0] _mesh_18_1_io_out_b_0;
	wire _mesh_18_1_io_out_control_0_dataflow;
	wire _mesh_18_1_io_out_control_0_propagate;
	wire [4:0] _mesh_18_1_io_out_control_0_shift;
	wire [2:0] _mesh_18_1_io_out_id_0;
	wire _mesh_18_1_io_out_last_0;
	wire _mesh_18_1_io_out_valid_0;
	wire [31:0] _mesh_18_0_io_out_a_0;
	wire [31:0] _mesh_18_0_io_out_c_0;
	wire [31:0] _mesh_18_0_io_out_b_0;
	wire _mesh_18_0_io_out_control_0_dataflow;
	wire _mesh_18_0_io_out_control_0_propagate;
	wire [4:0] _mesh_18_0_io_out_control_0_shift;
	wire [2:0] _mesh_18_0_io_out_id_0;
	wire _mesh_18_0_io_out_last_0;
	wire _mesh_18_0_io_out_valid_0;
	wire [31:0] _mesh_17_31_io_out_a_0;
	wire [31:0] _mesh_17_31_io_out_c_0;
	wire [31:0] _mesh_17_31_io_out_b_0;
	wire _mesh_17_31_io_out_control_0_dataflow;
	wire _mesh_17_31_io_out_control_0_propagate;
	wire [4:0] _mesh_17_31_io_out_control_0_shift;
	wire [2:0] _mesh_17_31_io_out_id_0;
	wire _mesh_17_31_io_out_last_0;
	wire _mesh_17_31_io_out_valid_0;
	wire [31:0] _mesh_17_30_io_out_a_0;
	wire [31:0] _mesh_17_30_io_out_c_0;
	wire [31:0] _mesh_17_30_io_out_b_0;
	wire _mesh_17_30_io_out_control_0_dataflow;
	wire _mesh_17_30_io_out_control_0_propagate;
	wire [4:0] _mesh_17_30_io_out_control_0_shift;
	wire [2:0] _mesh_17_30_io_out_id_0;
	wire _mesh_17_30_io_out_last_0;
	wire _mesh_17_30_io_out_valid_0;
	wire [31:0] _mesh_17_29_io_out_a_0;
	wire [31:0] _mesh_17_29_io_out_c_0;
	wire [31:0] _mesh_17_29_io_out_b_0;
	wire _mesh_17_29_io_out_control_0_dataflow;
	wire _mesh_17_29_io_out_control_0_propagate;
	wire [4:0] _mesh_17_29_io_out_control_0_shift;
	wire [2:0] _mesh_17_29_io_out_id_0;
	wire _mesh_17_29_io_out_last_0;
	wire _mesh_17_29_io_out_valid_0;
	wire [31:0] _mesh_17_28_io_out_a_0;
	wire [31:0] _mesh_17_28_io_out_c_0;
	wire [31:0] _mesh_17_28_io_out_b_0;
	wire _mesh_17_28_io_out_control_0_dataflow;
	wire _mesh_17_28_io_out_control_0_propagate;
	wire [4:0] _mesh_17_28_io_out_control_0_shift;
	wire [2:0] _mesh_17_28_io_out_id_0;
	wire _mesh_17_28_io_out_last_0;
	wire _mesh_17_28_io_out_valid_0;
	wire [31:0] _mesh_17_27_io_out_a_0;
	wire [31:0] _mesh_17_27_io_out_c_0;
	wire [31:0] _mesh_17_27_io_out_b_0;
	wire _mesh_17_27_io_out_control_0_dataflow;
	wire _mesh_17_27_io_out_control_0_propagate;
	wire [4:0] _mesh_17_27_io_out_control_0_shift;
	wire [2:0] _mesh_17_27_io_out_id_0;
	wire _mesh_17_27_io_out_last_0;
	wire _mesh_17_27_io_out_valid_0;
	wire [31:0] _mesh_17_26_io_out_a_0;
	wire [31:0] _mesh_17_26_io_out_c_0;
	wire [31:0] _mesh_17_26_io_out_b_0;
	wire _mesh_17_26_io_out_control_0_dataflow;
	wire _mesh_17_26_io_out_control_0_propagate;
	wire [4:0] _mesh_17_26_io_out_control_0_shift;
	wire [2:0] _mesh_17_26_io_out_id_0;
	wire _mesh_17_26_io_out_last_0;
	wire _mesh_17_26_io_out_valid_0;
	wire [31:0] _mesh_17_25_io_out_a_0;
	wire [31:0] _mesh_17_25_io_out_c_0;
	wire [31:0] _mesh_17_25_io_out_b_0;
	wire _mesh_17_25_io_out_control_0_dataflow;
	wire _mesh_17_25_io_out_control_0_propagate;
	wire [4:0] _mesh_17_25_io_out_control_0_shift;
	wire [2:0] _mesh_17_25_io_out_id_0;
	wire _mesh_17_25_io_out_last_0;
	wire _mesh_17_25_io_out_valid_0;
	wire [31:0] _mesh_17_24_io_out_a_0;
	wire [31:0] _mesh_17_24_io_out_c_0;
	wire [31:0] _mesh_17_24_io_out_b_0;
	wire _mesh_17_24_io_out_control_0_dataflow;
	wire _mesh_17_24_io_out_control_0_propagate;
	wire [4:0] _mesh_17_24_io_out_control_0_shift;
	wire [2:0] _mesh_17_24_io_out_id_0;
	wire _mesh_17_24_io_out_last_0;
	wire _mesh_17_24_io_out_valid_0;
	wire [31:0] _mesh_17_23_io_out_a_0;
	wire [31:0] _mesh_17_23_io_out_c_0;
	wire [31:0] _mesh_17_23_io_out_b_0;
	wire _mesh_17_23_io_out_control_0_dataflow;
	wire _mesh_17_23_io_out_control_0_propagate;
	wire [4:0] _mesh_17_23_io_out_control_0_shift;
	wire [2:0] _mesh_17_23_io_out_id_0;
	wire _mesh_17_23_io_out_last_0;
	wire _mesh_17_23_io_out_valid_0;
	wire [31:0] _mesh_17_22_io_out_a_0;
	wire [31:0] _mesh_17_22_io_out_c_0;
	wire [31:0] _mesh_17_22_io_out_b_0;
	wire _mesh_17_22_io_out_control_0_dataflow;
	wire _mesh_17_22_io_out_control_0_propagate;
	wire [4:0] _mesh_17_22_io_out_control_0_shift;
	wire [2:0] _mesh_17_22_io_out_id_0;
	wire _mesh_17_22_io_out_last_0;
	wire _mesh_17_22_io_out_valid_0;
	wire [31:0] _mesh_17_21_io_out_a_0;
	wire [31:0] _mesh_17_21_io_out_c_0;
	wire [31:0] _mesh_17_21_io_out_b_0;
	wire _mesh_17_21_io_out_control_0_dataflow;
	wire _mesh_17_21_io_out_control_0_propagate;
	wire [4:0] _mesh_17_21_io_out_control_0_shift;
	wire [2:0] _mesh_17_21_io_out_id_0;
	wire _mesh_17_21_io_out_last_0;
	wire _mesh_17_21_io_out_valid_0;
	wire [31:0] _mesh_17_20_io_out_a_0;
	wire [31:0] _mesh_17_20_io_out_c_0;
	wire [31:0] _mesh_17_20_io_out_b_0;
	wire _mesh_17_20_io_out_control_0_dataflow;
	wire _mesh_17_20_io_out_control_0_propagate;
	wire [4:0] _mesh_17_20_io_out_control_0_shift;
	wire [2:0] _mesh_17_20_io_out_id_0;
	wire _mesh_17_20_io_out_last_0;
	wire _mesh_17_20_io_out_valid_0;
	wire [31:0] _mesh_17_19_io_out_a_0;
	wire [31:0] _mesh_17_19_io_out_c_0;
	wire [31:0] _mesh_17_19_io_out_b_0;
	wire _mesh_17_19_io_out_control_0_dataflow;
	wire _mesh_17_19_io_out_control_0_propagate;
	wire [4:0] _mesh_17_19_io_out_control_0_shift;
	wire [2:0] _mesh_17_19_io_out_id_0;
	wire _mesh_17_19_io_out_last_0;
	wire _mesh_17_19_io_out_valid_0;
	wire [31:0] _mesh_17_18_io_out_a_0;
	wire [31:0] _mesh_17_18_io_out_c_0;
	wire [31:0] _mesh_17_18_io_out_b_0;
	wire _mesh_17_18_io_out_control_0_dataflow;
	wire _mesh_17_18_io_out_control_0_propagate;
	wire [4:0] _mesh_17_18_io_out_control_0_shift;
	wire [2:0] _mesh_17_18_io_out_id_0;
	wire _mesh_17_18_io_out_last_0;
	wire _mesh_17_18_io_out_valid_0;
	wire [31:0] _mesh_17_17_io_out_a_0;
	wire [31:0] _mesh_17_17_io_out_c_0;
	wire [31:0] _mesh_17_17_io_out_b_0;
	wire _mesh_17_17_io_out_control_0_dataflow;
	wire _mesh_17_17_io_out_control_0_propagate;
	wire [4:0] _mesh_17_17_io_out_control_0_shift;
	wire [2:0] _mesh_17_17_io_out_id_0;
	wire _mesh_17_17_io_out_last_0;
	wire _mesh_17_17_io_out_valid_0;
	wire [31:0] _mesh_17_16_io_out_a_0;
	wire [31:0] _mesh_17_16_io_out_c_0;
	wire [31:0] _mesh_17_16_io_out_b_0;
	wire _mesh_17_16_io_out_control_0_dataflow;
	wire _mesh_17_16_io_out_control_0_propagate;
	wire [4:0] _mesh_17_16_io_out_control_0_shift;
	wire [2:0] _mesh_17_16_io_out_id_0;
	wire _mesh_17_16_io_out_last_0;
	wire _mesh_17_16_io_out_valid_0;
	wire [31:0] _mesh_17_15_io_out_a_0;
	wire [31:0] _mesh_17_15_io_out_c_0;
	wire [31:0] _mesh_17_15_io_out_b_0;
	wire _mesh_17_15_io_out_control_0_dataflow;
	wire _mesh_17_15_io_out_control_0_propagate;
	wire [4:0] _mesh_17_15_io_out_control_0_shift;
	wire [2:0] _mesh_17_15_io_out_id_0;
	wire _mesh_17_15_io_out_last_0;
	wire _mesh_17_15_io_out_valid_0;
	wire [31:0] _mesh_17_14_io_out_a_0;
	wire [31:0] _mesh_17_14_io_out_c_0;
	wire [31:0] _mesh_17_14_io_out_b_0;
	wire _mesh_17_14_io_out_control_0_dataflow;
	wire _mesh_17_14_io_out_control_0_propagate;
	wire [4:0] _mesh_17_14_io_out_control_0_shift;
	wire [2:0] _mesh_17_14_io_out_id_0;
	wire _mesh_17_14_io_out_last_0;
	wire _mesh_17_14_io_out_valid_0;
	wire [31:0] _mesh_17_13_io_out_a_0;
	wire [31:0] _mesh_17_13_io_out_c_0;
	wire [31:0] _mesh_17_13_io_out_b_0;
	wire _mesh_17_13_io_out_control_0_dataflow;
	wire _mesh_17_13_io_out_control_0_propagate;
	wire [4:0] _mesh_17_13_io_out_control_0_shift;
	wire [2:0] _mesh_17_13_io_out_id_0;
	wire _mesh_17_13_io_out_last_0;
	wire _mesh_17_13_io_out_valid_0;
	wire [31:0] _mesh_17_12_io_out_a_0;
	wire [31:0] _mesh_17_12_io_out_c_0;
	wire [31:0] _mesh_17_12_io_out_b_0;
	wire _mesh_17_12_io_out_control_0_dataflow;
	wire _mesh_17_12_io_out_control_0_propagate;
	wire [4:0] _mesh_17_12_io_out_control_0_shift;
	wire [2:0] _mesh_17_12_io_out_id_0;
	wire _mesh_17_12_io_out_last_0;
	wire _mesh_17_12_io_out_valid_0;
	wire [31:0] _mesh_17_11_io_out_a_0;
	wire [31:0] _mesh_17_11_io_out_c_0;
	wire [31:0] _mesh_17_11_io_out_b_0;
	wire _mesh_17_11_io_out_control_0_dataflow;
	wire _mesh_17_11_io_out_control_0_propagate;
	wire [4:0] _mesh_17_11_io_out_control_0_shift;
	wire [2:0] _mesh_17_11_io_out_id_0;
	wire _mesh_17_11_io_out_last_0;
	wire _mesh_17_11_io_out_valid_0;
	wire [31:0] _mesh_17_10_io_out_a_0;
	wire [31:0] _mesh_17_10_io_out_c_0;
	wire [31:0] _mesh_17_10_io_out_b_0;
	wire _mesh_17_10_io_out_control_0_dataflow;
	wire _mesh_17_10_io_out_control_0_propagate;
	wire [4:0] _mesh_17_10_io_out_control_0_shift;
	wire [2:0] _mesh_17_10_io_out_id_0;
	wire _mesh_17_10_io_out_last_0;
	wire _mesh_17_10_io_out_valid_0;
	wire [31:0] _mesh_17_9_io_out_a_0;
	wire [31:0] _mesh_17_9_io_out_c_0;
	wire [31:0] _mesh_17_9_io_out_b_0;
	wire _mesh_17_9_io_out_control_0_dataflow;
	wire _mesh_17_9_io_out_control_0_propagate;
	wire [4:0] _mesh_17_9_io_out_control_0_shift;
	wire [2:0] _mesh_17_9_io_out_id_0;
	wire _mesh_17_9_io_out_last_0;
	wire _mesh_17_9_io_out_valid_0;
	wire [31:0] _mesh_17_8_io_out_a_0;
	wire [31:0] _mesh_17_8_io_out_c_0;
	wire [31:0] _mesh_17_8_io_out_b_0;
	wire _mesh_17_8_io_out_control_0_dataflow;
	wire _mesh_17_8_io_out_control_0_propagate;
	wire [4:0] _mesh_17_8_io_out_control_0_shift;
	wire [2:0] _mesh_17_8_io_out_id_0;
	wire _mesh_17_8_io_out_last_0;
	wire _mesh_17_8_io_out_valid_0;
	wire [31:0] _mesh_17_7_io_out_a_0;
	wire [31:0] _mesh_17_7_io_out_c_0;
	wire [31:0] _mesh_17_7_io_out_b_0;
	wire _mesh_17_7_io_out_control_0_dataflow;
	wire _mesh_17_7_io_out_control_0_propagate;
	wire [4:0] _mesh_17_7_io_out_control_0_shift;
	wire [2:0] _mesh_17_7_io_out_id_0;
	wire _mesh_17_7_io_out_last_0;
	wire _mesh_17_7_io_out_valid_0;
	wire [31:0] _mesh_17_6_io_out_a_0;
	wire [31:0] _mesh_17_6_io_out_c_0;
	wire [31:0] _mesh_17_6_io_out_b_0;
	wire _mesh_17_6_io_out_control_0_dataflow;
	wire _mesh_17_6_io_out_control_0_propagate;
	wire [4:0] _mesh_17_6_io_out_control_0_shift;
	wire [2:0] _mesh_17_6_io_out_id_0;
	wire _mesh_17_6_io_out_last_0;
	wire _mesh_17_6_io_out_valid_0;
	wire [31:0] _mesh_17_5_io_out_a_0;
	wire [31:0] _mesh_17_5_io_out_c_0;
	wire [31:0] _mesh_17_5_io_out_b_0;
	wire _mesh_17_5_io_out_control_0_dataflow;
	wire _mesh_17_5_io_out_control_0_propagate;
	wire [4:0] _mesh_17_5_io_out_control_0_shift;
	wire [2:0] _mesh_17_5_io_out_id_0;
	wire _mesh_17_5_io_out_last_0;
	wire _mesh_17_5_io_out_valid_0;
	wire [31:0] _mesh_17_4_io_out_a_0;
	wire [31:0] _mesh_17_4_io_out_c_0;
	wire [31:0] _mesh_17_4_io_out_b_0;
	wire _mesh_17_4_io_out_control_0_dataflow;
	wire _mesh_17_4_io_out_control_0_propagate;
	wire [4:0] _mesh_17_4_io_out_control_0_shift;
	wire [2:0] _mesh_17_4_io_out_id_0;
	wire _mesh_17_4_io_out_last_0;
	wire _mesh_17_4_io_out_valid_0;
	wire [31:0] _mesh_17_3_io_out_a_0;
	wire [31:0] _mesh_17_3_io_out_c_0;
	wire [31:0] _mesh_17_3_io_out_b_0;
	wire _mesh_17_3_io_out_control_0_dataflow;
	wire _mesh_17_3_io_out_control_0_propagate;
	wire [4:0] _mesh_17_3_io_out_control_0_shift;
	wire [2:0] _mesh_17_3_io_out_id_0;
	wire _mesh_17_3_io_out_last_0;
	wire _mesh_17_3_io_out_valid_0;
	wire [31:0] _mesh_17_2_io_out_a_0;
	wire [31:0] _mesh_17_2_io_out_c_0;
	wire [31:0] _mesh_17_2_io_out_b_0;
	wire _mesh_17_2_io_out_control_0_dataflow;
	wire _mesh_17_2_io_out_control_0_propagate;
	wire [4:0] _mesh_17_2_io_out_control_0_shift;
	wire [2:0] _mesh_17_2_io_out_id_0;
	wire _mesh_17_2_io_out_last_0;
	wire _mesh_17_2_io_out_valid_0;
	wire [31:0] _mesh_17_1_io_out_a_0;
	wire [31:0] _mesh_17_1_io_out_c_0;
	wire [31:0] _mesh_17_1_io_out_b_0;
	wire _mesh_17_1_io_out_control_0_dataflow;
	wire _mesh_17_1_io_out_control_0_propagate;
	wire [4:0] _mesh_17_1_io_out_control_0_shift;
	wire [2:0] _mesh_17_1_io_out_id_0;
	wire _mesh_17_1_io_out_last_0;
	wire _mesh_17_1_io_out_valid_0;
	wire [31:0] _mesh_17_0_io_out_a_0;
	wire [31:0] _mesh_17_0_io_out_c_0;
	wire [31:0] _mesh_17_0_io_out_b_0;
	wire _mesh_17_0_io_out_control_0_dataflow;
	wire _mesh_17_0_io_out_control_0_propagate;
	wire [4:0] _mesh_17_0_io_out_control_0_shift;
	wire [2:0] _mesh_17_0_io_out_id_0;
	wire _mesh_17_0_io_out_last_0;
	wire _mesh_17_0_io_out_valid_0;
	wire [31:0] _mesh_16_31_io_out_a_0;
	wire [31:0] _mesh_16_31_io_out_c_0;
	wire [31:0] _mesh_16_31_io_out_b_0;
	wire _mesh_16_31_io_out_control_0_dataflow;
	wire _mesh_16_31_io_out_control_0_propagate;
	wire [4:0] _mesh_16_31_io_out_control_0_shift;
	wire [2:0] _mesh_16_31_io_out_id_0;
	wire _mesh_16_31_io_out_last_0;
	wire _mesh_16_31_io_out_valid_0;
	wire [31:0] _mesh_16_30_io_out_a_0;
	wire [31:0] _mesh_16_30_io_out_c_0;
	wire [31:0] _mesh_16_30_io_out_b_0;
	wire _mesh_16_30_io_out_control_0_dataflow;
	wire _mesh_16_30_io_out_control_0_propagate;
	wire [4:0] _mesh_16_30_io_out_control_0_shift;
	wire [2:0] _mesh_16_30_io_out_id_0;
	wire _mesh_16_30_io_out_last_0;
	wire _mesh_16_30_io_out_valid_0;
	wire [31:0] _mesh_16_29_io_out_a_0;
	wire [31:0] _mesh_16_29_io_out_c_0;
	wire [31:0] _mesh_16_29_io_out_b_0;
	wire _mesh_16_29_io_out_control_0_dataflow;
	wire _mesh_16_29_io_out_control_0_propagate;
	wire [4:0] _mesh_16_29_io_out_control_0_shift;
	wire [2:0] _mesh_16_29_io_out_id_0;
	wire _mesh_16_29_io_out_last_0;
	wire _mesh_16_29_io_out_valid_0;
	wire [31:0] _mesh_16_28_io_out_a_0;
	wire [31:0] _mesh_16_28_io_out_c_0;
	wire [31:0] _mesh_16_28_io_out_b_0;
	wire _mesh_16_28_io_out_control_0_dataflow;
	wire _mesh_16_28_io_out_control_0_propagate;
	wire [4:0] _mesh_16_28_io_out_control_0_shift;
	wire [2:0] _mesh_16_28_io_out_id_0;
	wire _mesh_16_28_io_out_last_0;
	wire _mesh_16_28_io_out_valid_0;
	wire [31:0] _mesh_16_27_io_out_a_0;
	wire [31:0] _mesh_16_27_io_out_c_0;
	wire [31:0] _mesh_16_27_io_out_b_0;
	wire _mesh_16_27_io_out_control_0_dataflow;
	wire _mesh_16_27_io_out_control_0_propagate;
	wire [4:0] _mesh_16_27_io_out_control_0_shift;
	wire [2:0] _mesh_16_27_io_out_id_0;
	wire _mesh_16_27_io_out_last_0;
	wire _mesh_16_27_io_out_valid_0;
	wire [31:0] _mesh_16_26_io_out_a_0;
	wire [31:0] _mesh_16_26_io_out_c_0;
	wire [31:0] _mesh_16_26_io_out_b_0;
	wire _mesh_16_26_io_out_control_0_dataflow;
	wire _mesh_16_26_io_out_control_0_propagate;
	wire [4:0] _mesh_16_26_io_out_control_0_shift;
	wire [2:0] _mesh_16_26_io_out_id_0;
	wire _mesh_16_26_io_out_last_0;
	wire _mesh_16_26_io_out_valid_0;
	wire [31:0] _mesh_16_25_io_out_a_0;
	wire [31:0] _mesh_16_25_io_out_c_0;
	wire [31:0] _mesh_16_25_io_out_b_0;
	wire _mesh_16_25_io_out_control_0_dataflow;
	wire _mesh_16_25_io_out_control_0_propagate;
	wire [4:0] _mesh_16_25_io_out_control_0_shift;
	wire [2:0] _mesh_16_25_io_out_id_0;
	wire _mesh_16_25_io_out_last_0;
	wire _mesh_16_25_io_out_valid_0;
	wire [31:0] _mesh_16_24_io_out_a_0;
	wire [31:0] _mesh_16_24_io_out_c_0;
	wire [31:0] _mesh_16_24_io_out_b_0;
	wire _mesh_16_24_io_out_control_0_dataflow;
	wire _mesh_16_24_io_out_control_0_propagate;
	wire [4:0] _mesh_16_24_io_out_control_0_shift;
	wire [2:0] _mesh_16_24_io_out_id_0;
	wire _mesh_16_24_io_out_last_0;
	wire _mesh_16_24_io_out_valid_0;
	wire [31:0] _mesh_16_23_io_out_a_0;
	wire [31:0] _mesh_16_23_io_out_c_0;
	wire [31:0] _mesh_16_23_io_out_b_0;
	wire _mesh_16_23_io_out_control_0_dataflow;
	wire _mesh_16_23_io_out_control_0_propagate;
	wire [4:0] _mesh_16_23_io_out_control_0_shift;
	wire [2:0] _mesh_16_23_io_out_id_0;
	wire _mesh_16_23_io_out_last_0;
	wire _mesh_16_23_io_out_valid_0;
	wire [31:0] _mesh_16_22_io_out_a_0;
	wire [31:0] _mesh_16_22_io_out_c_0;
	wire [31:0] _mesh_16_22_io_out_b_0;
	wire _mesh_16_22_io_out_control_0_dataflow;
	wire _mesh_16_22_io_out_control_0_propagate;
	wire [4:0] _mesh_16_22_io_out_control_0_shift;
	wire [2:0] _mesh_16_22_io_out_id_0;
	wire _mesh_16_22_io_out_last_0;
	wire _mesh_16_22_io_out_valid_0;
	wire [31:0] _mesh_16_21_io_out_a_0;
	wire [31:0] _mesh_16_21_io_out_c_0;
	wire [31:0] _mesh_16_21_io_out_b_0;
	wire _mesh_16_21_io_out_control_0_dataflow;
	wire _mesh_16_21_io_out_control_0_propagate;
	wire [4:0] _mesh_16_21_io_out_control_0_shift;
	wire [2:0] _mesh_16_21_io_out_id_0;
	wire _mesh_16_21_io_out_last_0;
	wire _mesh_16_21_io_out_valid_0;
	wire [31:0] _mesh_16_20_io_out_a_0;
	wire [31:0] _mesh_16_20_io_out_c_0;
	wire [31:0] _mesh_16_20_io_out_b_0;
	wire _mesh_16_20_io_out_control_0_dataflow;
	wire _mesh_16_20_io_out_control_0_propagate;
	wire [4:0] _mesh_16_20_io_out_control_0_shift;
	wire [2:0] _mesh_16_20_io_out_id_0;
	wire _mesh_16_20_io_out_last_0;
	wire _mesh_16_20_io_out_valid_0;
	wire [31:0] _mesh_16_19_io_out_a_0;
	wire [31:0] _mesh_16_19_io_out_c_0;
	wire [31:0] _mesh_16_19_io_out_b_0;
	wire _mesh_16_19_io_out_control_0_dataflow;
	wire _mesh_16_19_io_out_control_0_propagate;
	wire [4:0] _mesh_16_19_io_out_control_0_shift;
	wire [2:0] _mesh_16_19_io_out_id_0;
	wire _mesh_16_19_io_out_last_0;
	wire _mesh_16_19_io_out_valid_0;
	wire [31:0] _mesh_16_18_io_out_a_0;
	wire [31:0] _mesh_16_18_io_out_c_0;
	wire [31:0] _mesh_16_18_io_out_b_0;
	wire _mesh_16_18_io_out_control_0_dataflow;
	wire _mesh_16_18_io_out_control_0_propagate;
	wire [4:0] _mesh_16_18_io_out_control_0_shift;
	wire [2:0] _mesh_16_18_io_out_id_0;
	wire _mesh_16_18_io_out_last_0;
	wire _mesh_16_18_io_out_valid_0;
	wire [31:0] _mesh_16_17_io_out_a_0;
	wire [31:0] _mesh_16_17_io_out_c_0;
	wire [31:0] _mesh_16_17_io_out_b_0;
	wire _mesh_16_17_io_out_control_0_dataflow;
	wire _mesh_16_17_io_out_control_0_propagate;
	wire [4:0] _mesh_16_17_io_out_control_0_shift;
	wire [2:0] _mesh_16_17_io_out_id_0;
	wire _mesh_16_17_io_out_last_0;
	wire _mesh_16_17_io_out_valid_0;
	wire [31:0] _mesh_16_16_io_out_a_0;
	wire [31:0] _mesh_16_16_io_out_c_0;
	wire [31:0] _mesh_16_16_io_out_b_0;
	wire _mesh_16_16_io_out_control_0_dataflow;
	wire _mesh_16_16_io_out_control_0_propagate;
	wire [4:0] _mesh_16_16_io_out_control_0_shift;
	wire [2:0] _mesh_16_16_io_out_id_0;
	wire _mesh_16_16_io_out_last_0;
	wire _mesh_16_16_io_out_valid_0;
	wire [31:0] _mesh_16_15_io_out_a_0;
	wire [31:0] _mesh_16_15_io_out_c_0;
	wire [31:0] _mesh_16_15_io_out_b_0;
	wire _mesh_16_15_io_out_control_0_dataflow;
	wire _mesh_16_15_io_out_control_0_propagate;
	wire [4:0] _mesh_16_15_io_out_control_0_shift;
	wire [2:0] _mesh_16_15_io_out_id_0;
	wire _mesh_16_15_io_out_last_0;
	wire _mesh_16_15_io_out_valid_0;
	wire [31:0] _mesh_16_14_io_out_a_0;
	wire [31:0] _mesh_16_14_io_out_c_0;
	wire [31:0] _mesh_16_14_io_out_b_0;
	wire _mesh_16_14_io_out_control_0_dataflow;
	wire _mesh_16_14_io_out_control_0_propagate;
	wire [4:0] _mesh_16_14_io_out_control_0_shift;
	wire [2:0] _mesh_16_14_io_out_id_0;
	wire _mesh_16_14_io_out_last_0;
	wire _mesh_16_14_io_out_valid_0;
	wire [31:0] _mesh_16_13_io_out_a_0;
	wire [31:0] _mesh_16_13_io_out_c_0;
	wire [31:0] _mesh_16_13_io_out_b_0;
	wire _mesh_16_13_io_out_control_0_dataflow;
	wire _mesh_16_13_io_out_control_0_propagate;
	wire [4:0] _mesh_16_13_io_out_control_0_shift;
	wire [2:0] _mesh_16_13_io_out_id_0;
	wire _mesh_16_13_io_out_last_0;
	wire _mesh_16_13_io_out_valid_0;
	wire [31:0] _mesh_16_12_io_out_a_0;
	wire [31:0] _mesh_16_12_io_out_c_0;
	wire [31:0] _mesh_16_12_io_out_b_0;
	wire _mesh_16_12_io_out_control_0_dataflow;
	wire _mesh_16_12_io_out_control_0_propagate;
	wire [4:0] _mesh_16_12_io_out_control_0_shift;
	wire [2:0] _mesh_16_12_io_out_id_0;
	wire _mesh_16_12_io_out_last_0;
	wire _mesh_16_12_io_out_valid_0;
	wire [31:0] _mesh_16_11_io_out_a_0;
	wire [31:0] _mesh_16_11_io_out_c_0;
	wire [31:0] _mesh_16_11_io_out_b_0;
	wire _mesh_16_11_io_out_control_0_dataflow;
	wire _mesh_16_11_io_out_control_0_propagate;
	wire [4:0] _mesh_16_11_io_out_control_0_shift;
	wire [2:0] _mesh_16_11_io_out_id_0;
	wire _mesh_16_11_io_out_last_0;
	wire _mesh_16_11_io_out_valid_0;
	wire [31:0] _mesh_16_10_io_out_a_0;
	wire [31:0] _mesh_16_10_io_out_c_0;
	wire [31:0] _mesh_16_10_io_out_b_0;
	wire _mesh_16_10_io_out_control_0_dataflow;
	wire _mesh_16_10_io_out_control_0_propagate;
	wire [4:0] _mesh_16_10_io_out_control_0_shift;
	wire [2:0] _mesh_16_10_io_out_id_0;
	wire _mesh_16_10_io_out_last_0;
	wire _mesh_16_10_io_out_valid_0;
	wire [31:0] _mesh_16_9_io_out_a_0;
	wire [31:0] _mesh_16_9_io_out_c_0;
	wire [31:0] _mesh_16_9_io_out_b_0;
	wire _mesh_16_9_io_out_control_0_dataflow;
	wire _mesh_16_9_io_out_control_0_propagate;
	wire [4:0] _mesh_16_9_io_out_control_0_shift;
	wire [2:0] _mesh_16_9_io_out_id_0;
	wire _mesh_16_9_io_out_last_0;
	wire _mesh_16_9_io_out_valid_0;
	wire [31:0] _mesh_16_8_io_out_a_0;
	wire [31:0] _mesh_16_8_io_out_c_0;
	wire [31:0] _mesh_16_8_io_out_b_0;
	wire _mesh_16_8_io_out_control_0_dataflow;
	wire _mesh_16_8_io_out_control_0_propagate;
	wire [4:0] _mesh_16_8_io_out_control_0_shift;
	wire [2:0] _mesh_16_8_io_out_id_0;
	wire _mesh_16_8_io_out_last_0;
	wire _mesh_16_8_io_out_valid_0;
	wire [31:0] _mesh_16_7_io_out_a_0;
	wire [31:0] _mesh_16_7_io_out_c_0;
	wire [31:0] _mesh_16_7_io_out_b_0;
	wire _mesh_16_7_io_out_control_0_dataflow;
	wire _mesh_16_7_io_out_control_0_propagate;
	wire [4:0] _mesh_16_7_io_out_control_0_shift;
	wire [2:0] _mesh_16_7_io_out_id_0;
	wire _mesh_16_7_io_out_last_0;
	wire _mesh_16_7_io_out_valid_0;
	wire [31:0] _mesh_16_6_io_out_a_0;
	wire [31:0] _mesh_16_6_io_out_c_0;
	wire [31:0] _mesh_16_6_io_out_b_0;
	wire _mesh_16_6_io_out_control_0_dataflow;
	wire _mesh_16_6_io_out_control_0_propagate;
	wire [4:0] _mesh_16_6_io_out_control_0_shift;
	wire [2:0] _mesh_16_6_io_out_id_0;
	wire _mesh_16_6_io_out_last_0;
	wire _mesh_16_6_io_out_valid_0;
	wire [31:0] _mesh_16_5_io_out_a_0;
	wire [31:0] _mesh_16_5_io_out_c_0;
	wire [31:0] _mesh_16_5_io_out_b_0;
	wire _mesh_16_5_io_out_control_0_dataflow;
	wire _mesh_16_5_io_out_control_0_propagate;
	wire [4:0] _mesh_16_5_io_out_control_0_shift;
	wire [2:0] _mesh_16_5_io_out_id_0;
	wire _mesh_16_5_io_out_last_0;
	wire _mesh_16_5_io_out_valid_0;
	wire [31:0] _mesh_16_4_io_out_a_0;
	wire [31:0] _mesh_16_4_io_out_c_0;
	wire [31:0] _mesh_16_4_io_out_b_0;
	wire _mesh_16_4_io_out_control_0_dataflow;
	wire _mesh_16_4_io_out_control_0_propagate;
	wire [4:0] _mesh_16_4_io_out_control_0_shift;
	wire [2:0] _mesh_16_4_io_out_id_0;
	wire _mesh_16_4_io_out_last_0;
	wire _mesh_16_4_io_out_valid_0;
	wire [31:0] _mesh_16_3_io_out_a_0;
	wire [31:0] _mesh_16_3_io_out_c_0;
	wire [31:0] _mesh_16_3_io_out_b_0;
	wire _mesh_16_3_io_out_control_0_dataflow;
	wire _mesh_16_3_io_out_control_0_propagate;
	wire [4:0] _mesh_16_3_io_out_control_0_shift;
	wire [2:0] _mesh_16_3_io_out_id_0;
	wire _mesh_16_3_io_out_last_0;
	wire _mesh_16_3_io_out_valid_0;
	wire [31:0] _mesh_16_2_io_out_a_0;
	wire [31:0] _mesh_16_2_io_out_c_0;
	wire [31:0] _mesh_16_2_io_out_b_0;
	wire _mesh_16_2_io_out_control_0_dataflow;
	wire _mesh_16_2_io_out_control_0_propagate;
	wire [4:0] _mesh_16_2_io_out_control_0_shift;
	wire [2:0] _mesh_16_2_io_out_id_0;
	wire _mesh_16_2_io_out_last_0;
	wire _mesh_16_2_io_out_valid_0;
	wire [31:0] _mesh_16_1_io_out_a_0;
	wire [31:0] _mesh_16_1_io_out_c_0;
	wire [31:0] _mesh_16_1_io_out_b_0;
	wire _mesh_16_1_io_out_control_0_dataflow;
	wire _mesh_16_1_io_out_control_0_propagate;
	wire [4:0] _mesh_16_1_io_out_control_0_shift;
	wire [2:0] _mesh_16_1_io_out_id_0;
	wire _mesh_16_1_io_out_last_0;
	wire _mesh_16_1_io_out_valid_0;
	wire [31:0] _mesh_16_0_io_out_a_0;
	wire [31:0] _mesh_16_0_io_out_c_0;
	wire [31:0] _mesh_16_0_io_out_b_0;
	wire _mesh_16_0_io_out_control_0_dataflow;
	wire _mesh_16_0_io_out_control_0_propagate;
	wire [4:0] _mesh_16_0_io_out_control_0_shift;
	wire [2:0] _mesh_16_0_io_out_id_0;
	wire _mesh_16_0_io_out_last_0;
	wire _mesh_16_0_io_out_valid_0;
	wire [31:0] _mesh_15_31_io_out_a_0;
	wire [31:0] _mesh_15_31_io_out_c_0;
	wire [31:0] _mesh_15_31_io_out_b_0;
	wire _mesh_15_31_io_out_control_0_dataflow;
	wire _mesh_15_31_io_out_control_0_propagate;
	wire [4:0] _mesh_15_31_io_out_control_0_shift;
	wire [2:0] _mesh_15_31_io_out_id_0;
	wire _mesh_15_31_io_out_last_0;
	wire _mesh_15_31_io_out_valid_0;
	wire [31:0] _mesh_15_30_io_out_a_0;
	wire [31:0] _mesh_15_30_io_out_c_0;
	wire [31:0] _mesh_15_30_io_out_b_0;
	wire _mesh_15_30_io_out_control_0_dataflow;
	wire _mesh_15_30_io_out_control_0_propagate;
	wire [4:0] _mesh_15_30_io_out_control_0_shift;
	wire [2:0] _mesh_15_30_io_out_id_0;
	wire _mesh_15_30_io_out_last_0;
	wire _mesh_15_30_io_out_valid_0;
	wire [31:0] _mesh_15_29_io_out_a_0;
	wire [31:0] _mesh_15_29_io_out_c_0;
	wire [31:0] _mesh_15_29_io_out_b_0;
	wire _mesh_15_29_io_out_control_0_dataflow;
	wire _mesh_15_29_io_out_control_0_propagate;
	wire [4:0] _mesh_15_29_io_out_control_0_shift;
	wire [2:0] _mesh_15_29_io_out_id_0;
	wire _mesh_15_29_io_out_last_0;
	wire _mesh_15_29_io_out_valid_0;
	wire [31:0] _mesh_15_28_io_out_a_0;
	wire [31:0] _mesh_15_28_io_out_c_0;
	wire [31:0] _mesh_15_28_io_out_b_0;
	wire _mesh_15_28_io_out_control_0_dataflow;
	wire _mesh_15_28_io_out_control_0_propagate;
	wire [4:0] _mesh_15_28_io_out_control_0_shift;
	wire [2:0] _mesh_15_28_io_out_id_0;
	wire _mesh_15_28_io_out_last_0;
	wire _mesh_15_28_io_out_valid_0;
	wire [31:0] _mesh_15_27_io_out_a_0;
	wire [31:0] _mesh_15_27_io_out_c_0;
	wire [31:0] _mesh_15_27_io_out_b_0;
	wire _mesh_15_27_io_out_control_0_dataflow;
	wire _mesh_15_27_io_out_control_0_propagate;
	wire [4:0] _mesh_15_27_io_out_control_0_shift;
	wire [2:0] _mesh_15_27_io_out_id_0;
	wire _mesh_15_27_io_out_last_0;
	wire _mesh_15_27_io_out_valid_0;
	wire [31:0] _mesh_15_26_io_out_a_0;
	wire [31:0] _mesh_15_26_io_out_c_0;
	wire [31:0] _mesh_15_26_io_out_b_0;
	wire _mesh_15_26_io_out_control_0_dataflow;
	wire _mesh_15_26_io_out_control_0_propagate;
	wire [4:0] _mesh_15_26_io_out_control_0_shift;
	wire [2:0] _mesh_15_26_io_out_id_0;
	wire _mesh_15_26_io_out_last_0;
	wire _mesh_15_26_io_out_valid_0;
	wire [31:0] _mesh_15_25_io_out_a_0;
	wire [31:0] _mesh_15_25_io_out_c_0;
	wire [31:0] _mesh_15_25_io_out_b_0;
	wire _mesh_15_25_io_out_control_0_dataflow;
	wire _mesh_15_25_io_out_control_0_propagate;
	wire [4:0] _mesh_15_25_io_out_control_0_shift;
	wire [2:0] _mesh_15_25_io_out_id_0;
	wire _mesh_15_25_io_out_last_0;
	wire _mesh_15_25_io_out_valid_0;
	wire [31:0] _mesh_15_24_io_out_a_0;
	wire [31:0] _mesh_15_24_io_out_c_0;
	wire [31:0] _mesh_15_24_io_out_b_0;
	wire _mesh_15_24_io_out_control_0_dataflow;
	wire _mesh_15_24_io_out_control_0_propagate;
	wire [4:0] _mesh_15_24_io_out_control_0_shift;
	wire [2:0] _mesh_15_24_io_out_id_0;
	wire _mesh_15_24_io_out_last_0;
	wire _mesh_15_24_io_out_valid_0;
	wire [31:0] _mesh_15_23_io_out_a_0;
	wire [31:0] _mesh_15_23_io_out_c_0;
	wire [31:0] _mesh_15_23_io_out_b_0;
	wire _mesh_15_23_io_out_control_0_dataflow;
	wire _mesh_15_23_io_out_control_0_propagate;
	wire [4:0] _mesh_15_23_io_out_control_0_shift;
	wire [2:0] _mesh_15_23_io_out_id_0;
	wire _mesh_15_23_io_out_last_0;
	wire _mesh_15_23_io_out_valid_0;
	wire [31:0] _mesh_15_22_io_out_a_0;
	wire [31:0] _mesh_15_22_io_out_c_0;
	wire [31:0] _mesh_15_22_io_out_b_0;
	wire _mesh_15_22_io_out_control_0_dataflow;
	wire _mesh_15_22_io_out_control_0_propagate;
	wire [4:0] _mesh_15_22_io_out_control_0_shift;
	wire [2:0] _mesh_15_22_io_out_id_0;
	wire _mesh_15_22_io_out_last_0;
	wire _mesh_15_22_io_out_valid_0;
	wire [31:0] _mesh_15_21_io_out_a_0;
	wire [31:0] _mesh_15_21_io_out_c_0;
	wire [31:0] _mesh_15_21_io_out_b_0;
	wire _mesh_15_21_io_out_control_0_dataflow;
	wire _mesh_15_21_io_out_control_0_propagate;
	wire [4:0] _mesh_15_21_io_out_control_0_shift;
	wire [2:0] _mesh_15_21_io_out_id_0;
	wire _mesh_15_21_io_out_last_0;
	wire _mesh_15_21_io_out_valid_0;
	wire [31:0] _mesh_15_20_io_out_a_0;
	wire [31:0] _mesh_15_20_io_out_c_0;
	wire [31:0] _mesh_15_20_io_out_b_0;
	wire _mesh_15_20_io_out_control_0_dataflow;
	wire _mesh_15_20_io_out_control_0_propagate;
	wire [4:0] _mesh_15_20_io_out_control_0_shift;
	wire [2:0] _mesh_15_20_io_out_id_0;
	wire _mesh_15_20_io_out_last_0;
	wire _mesh_15_20_io_out_valid_0;
	wire [31:0] _mesh_15_19_io_out_a_0;
	wire [31:0] _mesh_15_19_io_out_c_0;
	wire [31:0] _mesh_15_19_io_out_b_0;
	wire _mesh_15_19_io_out_control_0_dataflow;
	wire _mesh_15_19_io_out_control_0_propagate;
	wire [4:0] _mesh_15_19_io_out_control_0_shift;
	wire [2:0] _mesh_15_19_io_out_id_0;
	wire _mesh_15_19_io_out_last_0;
	wire _mesh_15_19_io_out_valid_0;
	wire [31:0] _mesh_15_18_io_out_a_0;
	wire [31:0] _mesh_15_18_io_out_c_0;
	wire [31:0] _mesh_15_18_io_out_b_0;
	wire _mesh_15_18_io_out_control_0_dataflow;
	wire _mesh_15_18_io_out_control_0_propagate;
	wire [4:0] _mesh_15_18_io_out_control_0_shift;
	wire [2:0] _mesh_15_18_io_out_id_0;
	wire _mesh_15_18_io_out_last_0;
	wire _mesh_15_18_io_out_valid_0;
	wire [31:0] _mesh_15_17_io_out_a_0;
	wire [31:0] _mesh_15_17_io_out_c_0;
	wire [31:0] _mesh_15_17_io_out_b_0;
	wire _mesh_15_17_io_out_control_0_dataflow;
	wire _mesh_15_17_io_out_control_0_propagate;
	wire [4:0] _mesh_15_17_io_out_control_0_shift;
	wire [2:0] _mesh_15_17_io_out_id_0;
	wire _mesh_15_17_io_out_last_0;
	wire _mesh_15_17_io_out_valid_0;
	wire [31:0] _mesh_15_16_io_out_a_0;
	wire [31:0] _mesh_15_16_io_out_c_0;
	wire [31:0] _mesh_15_16_io_out_b_0;
	wire _mesh_15_16_io_out_control_0_dataflow;
	wire _mesh_15_16_io_out_control_0_propagate;
	wire [4:0] _mesh_15_16_io_out_control_0_shift;
	wire [2:0] _mesh_15_16_io_out_id_0;
	wire _mesh_15_16_io_out_last_0;
	wire _mesh_15_16_io_out_valid_0;
	wire [31:0] _mesh_15_15_io_out_a_0;
	wire [31:0] _mesh_15_15_io_out_c_0;
	wire [31:0] _mesh_15_15_io_out_b_0;
	wire _mesh_15_15_io_out_control_0_dataflow;
	wire _mesh_15_15_io_out_control_0_propagate;
	wire [4:0] _mesh_15_15_io_out_control_0_shift;
	wire [2:0] _mesh_15_15_io_out_id_0;
	wire _mesh_15_15_io_out_last_0;
	wire _mesh_15_15_io_out_valid_0;
	wire [31:0] _mesh_15_14_io_out_a_0;
	wire [31:0] _mesh_15_14_io_out_c_0;
	wire [31:0] _mesh_15_14_io_out_b_0;
	wire _mesh_15_14_io_out_control_0_dataflow;
	wire _mesh_15_14_io_out_control_0_propagate;
	wire [4:0] _mesh_15_14_io_out_control_0_shift;
	wire [2:0] _mesh_15_14_io_out_id_0;
	wire _mesh_15_14_io_out_last_0;
	wire _mesh_15_14_io_out_valid_0;
	wire [31:0] _mesh_15_13_io_out_a_0;
	wire [31:0] _mesh_15_13_io_out_c_0;
	wire [31:0] _mesh_15_13_io_out_b_0;
	wire _mesh_15_13_io_out_control_0_dataflow;
	wire _mesh_15_13_io_out_control_0_propagate;
	wire [4:0] _mesh_15_13_io_out_control_0_shift;
	wire [2:0] _mesh_15_13_io_out_id_0;
	wire _mesh_15_13_io_out_last_0;
	wire _mesh_15_13_io_out_valid_0;
	wire [31:0] _mesh_15_12_io_out_a_0;
	wire [31:0] _mesh_15_12_io_out_c_0;
	wire [31:0] _mesh_15_12_io_out_b_0;
	wire _mesh_15_12_io_out_control_0_dataflow;
	wire _mesh_15_12_io_out_control_0_propagate;
	wire [4:0] _mesh_15_12_io_out_control_0_shift;
	wire [2:0] _mesh_15_12_io_out_id_0;
	wire _mesh_15_12_io_out_last_0;
	wire _mesh_15_12_io_out_valid_0;
	wire [31:0] _mesh_15_11_io_out_a_0;
	wire [31:0] _mesh_15_11_io_out_c_0;
	wire [31:0] _mesh_15_11_io_out_b_0;
	wire _mesh_15_11_io_out_control_0_dataflow;
	wire _mesh_15_11_io_out_control_0_propagate;
	wire [4:0] _mesh_15_11_io_out_control_0_shift;
	wire [2:0] _mesh_15_11_io_out_id_0;
	wire _mesh_15_11_io_out_last_0;
	wire _mesh_15_11_io_out_valid_0;
	wire [31:0] _mesh_15_10_io_out_a_0;
	wire [31:0] _mesh_15_10_io_out_c_0;
	wire [31:0] _mesh_15_10_io_out_b_0;
	wire _mesh_15_10_io_out_control_0_dataflow;
	wire _mesh_15_10_io_out_control_0_propagate;
	wire [4:0] _mesh_15_10_io_out_control_0_shift;
	wire [2:0] _mesh_15_10_io_out_id_0;
	wire _mesh_15_10_io_out_last_0;
	wire _mesh_15_10_io_out_valid_0;
	wire [31:0] _mesh_15_9_io_out_a_0;
	wire [31:0] _mesh_15_9_io_out_c_0;
	wire [31:0] _mesh_15_9_io_out_b_0;
	wire _mesh_15_9_io_out_control_0_dataflow;
	wire _mesh_15_9_io_out_control_0_propagate;
	wire [4:0] _mesh_15_9_io_out_control_0_shift;
	wire [2:0] _mesh_15_9_io_out_id_0;
	wire _mesh_15_9_io_out_last_0;
	wire _mesh_15_9_io_out_valid_0;
	wire [31:0] _mesh_15_8_io_out_a_0;
	wire [31:0] _mesh_15_8_io_out_c_0;
	wire [31:0] _mesh_15_8_io_out_b_0;
	wire _mesh_15_8_io_out_control_0_dataflow;
	wire _mesh_15_8_io_out_control_0_propagate;
	wire [4:0] _mesh_15_8_io_out_control_0_shift;
	wire [2:0] _mesh_15_8_io_out_id_0;
	wire _mesh_15_8_io_out_last_0;
	wire _mesh_15_8_io_out_valid_0;
	wire [31:0] _mesh_15_7_io_out_a_0;
	wire [31:0] _mesh_15_7_io_out_c_0;
	wire [31:0] _mesh_15_7_io_out_b_0;
	wire _mesh_15_7_io_out_control_0_dataflow;
	wire _mesh_15_7_io_out_control_0_propagate;
	wire [4:0] _mesh_15_7_io_out_control_0_shift;
	wire [2:0] _mesh_15_7_io_out_id_0;
	wire _mesh_15_7_io_out_last_0;
	wire _mesh_15_7_io_out_valid_0;
	wire [31:0] _mesh_15_6_io_out_a_0;
	wire [31:0] _mesh_15_6_io_out_c_0;
	wire [31:0] _mesh_15_6_io_out_b_0;
	wire _mesh_15_6_io_out_control_0_dataflow;
	wire _mesh_15_6_io_out_control_0_propagate;
	wire [4:0] _mesh_15_6_io_out_control_0_shift;
	wire [2:0] _mesh_15_6_io_out_id_0;
	wire _mesh_15_6_io_out_last_0;
	wire _mesh_15_6_io_out_valid_0;
	wire [31:0] _mesh_15_5_io_out_a_0;
	wire [31:0] _mesh_15_5_io_out_c_0;
	wire [31:0] _mesh_15_5_io_out_b_0;
	wire _mesh_15_5_io_out_control_0_dataflow;
	wire _mesh_15_5_io_out_control_0_propagate;
	wire [4:0] _mesh_15_5_io_out_control_0_shift;
	wire [2:0] _mesh_15_5_io_out_id_0;
	wire _mesh_15_5_io_out_last_0;
	wire _mesh_15_5_io_out_valid_0;
	wire [31:0] _mesh_15_4_io_out_a_0;
	wire [31:0] _mesh_15_4_io_out_c_0;
	wire [31:0] _mesh_15_4_io_out_b_0;
	wire _mesh_15_4_io_out_control_0_dataflow;
	wire _mesh_15_4_io_out_control_0_propagate;
	wire [4:0] _mesh_15_4_io_out_control_0_shift;
	wire [2:0] _mesh_15_4_io_out_id_0;
	wire _mesh_15_4_io_out_last_0;
	wire _mesh_15_4_io_out_valid_0;
	wire [31:0] _mesh_15_3_io_out_a_0;
	wire [31:0] _mesh_15_3_io_out_c_0;
	wire [31:0] _mesh_15_3_io_out_b_0;
	wire _mesh_15_3_io_out_control_0_dataflow;
	wire _mesh_15_3_io_out_control_0_propagate;
	wire [4:0] _mesh_15_3_io_out_control_0_shift;
	wire [2:0] _mesh_15_3_io_out_id_0;
	wire _mesh_15_3_io_out_last_0;
	wire _mesh_15_3_io_out_valid_0;
	wire [31:0] _mesh_15_2_io_out_a_0;
	wire [31:0] _mesh_15_2_io_out_c_0;
	wire [31:0] _mesh_15_2_io_out_b_0;
	wire _mesh_15_2_io_out_control_0_dataflow;
	wire _mesh_15_2_io_out_control_0_propagate;
	wire [4:0] _mesh_15_2_io_out_control_0_shift;
	wire [2:0] _mesh_15_2_io_out_id_0;
	wire _mesh_15_2_io_out_last_0;
	wire _mesh_15_2_io_out_valid_0;
	wire [31:0] _mesh_15_1_io_out_a_0;
	wire [31:0] _mesh_15_1_io_out_c_0;
	wire [31:0] _mesh_15_1_io_out_b_0;
	wire _mesh_15_1_io_out_control_0_dataflow;
	wire _mesh_15_1_io_out_control_0_propagate;
	wire [4:0] _mesh_15_1_io_out_control_0_shift;
	wire [2:0] _mesh_15_1_io_out_id_0;
	wire _mesh_15_1_io_out_last_0;
	wire _mesh_15_1_io_out_valid_0;
	wire [31:0] _mesh_15_0_io_out_a_0;
	wire [31:0] _mesh_15_0_io_out_c_0;
	wire [31:0] _mesh_15_0_io_out_b_0;
	wire _mesh_15_0_io_out_control_0_dataflow;
	wire _mesh_15_0_io_out_control_0_propagate;
	wire [4:0] _mesh_15_0_io_out_control_0_shift;
	wire [2:0] _mesh_15_0_io_out_id_0;
	wire _mesh_15_0_io_out_last_0;
	wire _mesh_15_0_io_out_valid_0;
	wire [31:0] _mesh_14_31_io_out_a_0;
	wire [31:0] _mesh_14_31_io_out_c_0;
	wire [31:0] _mesh_14_31_io_out_b_0;
	wire _mesh_14_31_io_out_control_0_dataflow;
	wire _mesh_14_31_io_out_control_0_propagate;
	wire [4:0] _mesh_14_31_io_out_control_0_shift;
	wire [2:0] _mesh_14_31_io_out_id_0;
	wire _mesh_14_31_io_out_last_0;
	wire _mesh_14_31_io_out_valid_0;
	wire [31:0] _mesh_14_30_io_out_a_0;
	wire [31:0] _mesh_14_30_io_out_c_0;
	wire [31:0] _mesh_14_30_io_out_b_0;
	wire _mesh_14_30_io_out_control_0_dataflow;
	wire _mesh_14_30_io_out_control_0_propagate;
	wire [4:0] _mesh_14_30_io_out_control_0_shift;
	wire [2:0] _mesh_14_30_io_out_id_0;
	wire _mesh_14_30_io_out_last_0;
	wire _mesh_14_30_io_out_valid_0;
	wire [31:0] _mesh_14_29_io_out_a_0;
	wire [31:0] _mesh_14_29_io_out_c_0;
	wire [31:0] _mesh_14_29_io_out_b_0;
	wire _mesh_14_29_io_out_control_0_dataflow;
	wire _mesh_14_29_io_out_control_0_propagate;
	wire [4:0] _mesh_14_29_io_out_control_0_shift;
	wire [2:0] _mesh_14_29_io_out_id_0;
	wire _mesh_14_29_io_out_last_0;
	wire _mesh_14_29_io_out_valid_0;
	wire [31:0] _mesh_14_28_io_out_a_0;
	wire [31:0] _mesh_14_28_io_out_c_0;
	wire [31:0] _mesh_14_28_io_out_b_0;
	wire _mesh_14_28_io_out_control_0_dataflow;
	wire _mesh_14_28_io_out_control_0_propagate;
	wire [4:0] _mesh_14_28_io_out_control_0_shift;
	wire [2:0] _mesh_14_28_io_out_id_0;
	wire _mesh_14_28_io_out_last_0;
	wire _mesh_14_28_io_out_valid_0;
	wire [31:0] _mesh_14_27_io_out_a_0;
	wire [31:0] _mesh_14_27_io_out_c_0;
	wire [31:0] _mesh_14_27_io_out_b_0;
	wire _mesh_14_27_io_out_control_0_dataflow;
	wire _mesh_14_27_io_out_control_0_propagate;
	wire [4:0] _mesh_14_27_io_out_control_0_shift;
	wire [2:0] _mesh_14_27_io_out_id_0;
	wire _mesh_14_27_io_out_last_0;
	wire _mesh_14_27_io_out_valid_0;
	wire [31:0] _mesh_14_26_io_out_a_0;
	wire [31:0] _mesh_14_26_io_out_c_0;
	wire [31:0] _mesh_14_26_io_out_b_0;
	wire _mesh_14_26_io_out_control_0_dataflow;
	wire _mesh_14_26_io_out_control_0_propagate;
	wire [4:0] _mesh_14_26_io_out_control_0_shift;
	wire [2:0] _mesh_14_26_io_out_id_0;
	wire _mesh_14_26_io_out_last_0;
	wire _mesh_14_26_io_out_valid_0;
	wire [31:0] _mesh_14_25_io_out_a_0;
	wire [31:0] _mesh_14_25_io_out_c_0;
	wire [31:0] _mesh_14_25_io_out_b_0;
	wire _mesh_14_25_io_out_control_0_dataflow;
	wire _mesh_14_25_io_out_control_0_propagate;
	wire [4:0] _mesh_14_25_io_out_control_0_shift;
	wire [2:0] _mesh_14_25_io_out_id_0;
	wire _mesh_14_25_io_out_last_0;
	wire _mesh_14_25_io_out_valid_0;
	wire [31:0] _mesh_14_24_io_out_a_0;
	wire [31:0] _mesh_14_24_io_out_c_0;
	wire [31:0] _mesh_14_24_io_out_b_0;
	wire _mesh_14_24_io_out_control_0_dataflow;
	wire _mesh_14_24_io_out_control_0_propagate;
	wire [4:0] _mesh_14_24_io_out_control_0_shift;
	wire [2:0] _mesh_14_24_io_out_id_0;
	wire _mesh_14_24_io_out_last_0;
	wire _mesh_14_24_io_out_valid_0;
	wire [31:0] _mesh_14_23_io_out_a_0;
	wire [31:0] _mesh_14_23_io_out_c_0;
	wire [31:0] _mesh_14_23_io_out_b_0;
	wire _mesh_14_23_io_out_control_0_dataflow;
	wire _mesh_14_23_io_out_control_0_propagate;
	wire [4:0] _mesh_14_23_io_out_control_0_shift;
	wire [2:0] _mesh_14_23_io_out_id_0;
	wire _mesh_14_23_io_out_last_0;
	wire _mesh_14_23_io_out_valid_0;
	wire [31:0] _mesh_14_22_io_out_a_0;
	wire [31:0] _mesh_14_22_io_out_c_0;
	wire [31:0] _mesh_14_22_io_out_b_0;
	wire _mesh_14_22_io_out_control_0_dataflow;
	wire _mesh_14_22_io_out_control_0_propagate;
	wire [4:0] _mesh_14_22_io_out_control_0_shift;
	wire [2:0] _mesh_14_22_io_out_id_0;
	wire _mesh_14_22_io_out_last_0;
	wire _mesh_14_22_io_out_valid_0;
	wire [31:0] _mesh_14_21_io_out_a_0;
	wire [31:0] _mesh_14_21_io_out_c_0;
	wire [31:0] _mesh_14_21_io_out_b_0;
	wire _mesh_14_21_io_out_control_0_dataflow;
	wire _mesh_14_21_io_out_control_0_propagate;
	wire [4:0] _mesh_14_21_io_out_control_0_shift;
	wire [2:0] _mesh_14_21_io_out_id_0;
	wire _mesh_14_21_io_out_last_0;
	wire _mesh_14_21_io_out_valid_0;
	wire [31:0] _mesh_14_20_io_out_a_0;
	wire [31:0] _mesh_14_20_io_out_c_0;
	wire [31:0] _mesh_14_20_io_out_b_0;
	wire _mesh_14_20_io_out_control_0_dataflow;
	wire _mesh_14_20_io_out_control_0_propagate;
	wire [4:0] _mesh_14_20_io_out_control_0_shift;
	wire [2:0] _mesh_14_20_io_out_id_0;
	wire _mesh_14_20_io_out_last_0;
	wire _mesh_14_20_io_out_valid_0;
	wire [31:0] _mesh_14_19_io_out_a_0;
	wire [31:0] _mesh_14_19_io_out_c_0;
	wire [31:0] _mesh_14_19_io_out_b_0;
	wire _mesh_14_19_io_out_control_0_dataflow;
	wire _mesh_14_19_io_out_control_0_propagate;
	wire [4:0] _mesh_14_19_io_out_control_0_shift;
	wire [2:0] _mesh_14_19_io_out_id_0;
	wire _mesh_14_19_io_out_last_0;
	wire _mesh_14_19_io_out_valid_0;
	wire [31:0] _mesh_14_18_io_out_a_0;
	wire [31:0] _mesh_14_18_io_out_c_0;
	wire [31:0] _mesh_14_18_io_out_b_0;
	wire _mesh_14_18_io_out_control_0_dataflow;
	wire _mesh_14_18_io_out_control_0_propagate;
	wire [4:0] _mesh_14_18_io_out_control_0_shift;
	wire [2:0] _mesh_14_18_io_out_id_0;
	wire _mesh_14_18_io_out_last_0;
	wire _mesh_14_18_io_out_valid_0;
	wire [31:0] _mesh_14_17_io_out_a_0;
	wire [31:0] _mesh_14_17_io_out_c_0;
	wire [31:0] _mesh_14_17_io_out_b_0;
	wire _mesh_14_17_io_out_control_0_dataflow;
	wire _mesh_14_17_io_out_control_0_propagate;
	wire [4:0] _mesh_14_17_io_out_control_0_shift;
	wire [2:0] _mesh_14_17_io_out_id_0;
	wire _mesh_14_17_io_out_last_0;
	wire _mesh_14_17_io_out_valid_0;
	wire [31:0] _mesh_14_16_io_out_a_0;
	wire [31:0] _mesh_14_16_io_out_c_0;
	wire [31:0] _mesh_14_16_io_out_b_0;
	wire _mesh_14_16_io_out_control_0_dataflow;
	wire _mesh_14_16_io_out_control_0_propagate;
	wire [4:0] _mesh_14_16_io_out_control_0_shift;
	wire [2:0] _mesh_14_16_io_out_id_0;
	wire _mesh_14_16_io_out_last_0;
	wire _mesh_14_16_io_out_valid_0;
	wire [31:0] _mesh_14_15_io_out_a_0;
	wire [31:0] _mesh_14_15_io_out_c_0;
	wire [31:0] _mesh_14_15_io_out_b_0;
	wire _mesh_14_15_io_out_control_0_dataflow;
	wire _mesh_14_15_io_out_control_0_propagate;
	wire [4:0] _mesh_14_15_io_out_control_0_shift;
	wire [2:0] _mesh_14_15_io_out_id_0;
	wire _mesh_14_15_io_out_last_0;
	wire _mesh_14_15_io_out_valid_0;
	wire [31:0] _mesh_14_14_io_out_a_0;
	wire [31:0] _mesh_14_14_io_out_c_0;
	wire [31:0] _mesh_14_14_io_out_b_0;
	wire _mesh_14_14_io_out_control_0_dataflow;
	wire _mesh_14_14_io_out_control_0_propagate;
	wire [4:0] _mesh_14_14_io_out_control_0_shift;
	wire [2:0] _mesh_14_14_io_out_id_0;
	wire _mesh_14_14_io_out_last_0;
	wire _mesh_14_14_io_out_valid_0;
	wire [31:0] _mesh_14_13_io_out_a_0;
	wire [31:0] _mesh_14_13_io_out_c_0;
	wire [31:0] _mesh_14_13_io_out_b_0;
	wire _mesh_14_13_io_out_control_0_dataflow;
	wire _mesh_14_13_io_out_control_0_propagate;
	wire [4:0] _mesh_14_13_io_out_control_0_shift;
	wire [2:0] _mesh_14_13_io_out_id_0;
	wire _mesh_14_13_io_out_last_0;
	wire _mesh_14_13_io_out_valid_0;
	wire [31:0] _mesh_14_12_io_out_a_0;
	wire [31:0] _mesh_14_12_io_out_c_0;
	wire [31:0] _mesh_14_12_io_out_b_0;
	wire _mesh_14_12_io_out_control_0_dataflow;
	wire _mesh_14_12_io_out_control_0_propagate;
	wire [4:0] _mesh_14_12_io_out_control_0_shift;
	wire [2:0] _mesh_14_12_io_out_id_0;
	wire _mesh_14_12_io_out_last_0;
	wire _mesh_14_12_io_out_valid_0;
	wire [31:0] _mesh_14_11_io_out_a_0;
	wire [31:0] _mesh_14_11_io_out_c_0;
	wire [31:0] _mesh_14_11_io_out_b_0;
	wire _mesh_14_11_io_out_control_0_dataflow;
	wire _mesh_14_11_io_out_control_0_propagate;
	wire [4:0] _mesh_14_11_io_out_control_0_shift;
	wire [2:0] _mesh_14_11_io_out_id_0;
	wire _mesh_14_11_io_out_last_0;
	wire _mesh_14_11_io_out_valid_0;
	wire [31:0] _mesh_14_10_io_out_a_0;
	wire [31:0] _mesh_14_10_io_out_c_0;
	wire [31:0] _mesh_14_10_io_out_b_0;
	wire _mesh_14_10_io_out_control_0_dataflow;
	wire _mesh_14_10_io_out_control_0_propagate;
	wire [4:0] _mesh_14_10_io_out_control_0_shift;
	wire [2:0] _mesh_14_10_io_out_id_0;
	wire _mesh_14_10_io_out_last_0;
	wire _mesh_14_10_io_out_valid_0;
	wire [31:0] _mesh_14_9_io_out_a_0;
	wire [31:0] _mesh_14_9_io_out_c_0;
	wire [31:0] _mesh_14_9_io_out_b_0;
	wire _mesh_14_9_io_out_control_0_dataflow;
	wire _mesh_14_9_io_out_control_0_propagate;
	wire [4:0] _mesh_14_9_io_out_control_0_shift;
	wire [2:0] _mesh_14_9_io_out_id_0;
	wire _mesh_14_9_io_out_last_0;
	wire _mesh_14_9_io_out_valid_0;
	wire [31:0] _mesh_14_8_io_out_a_0;
	wire [31:0] _mesh_14_8_io_out_c_0;
	wire [31:0] _mesh_14_8_io_out_b_0;
	wire _mesh_14_8_io_out_control_0_dataflow;
	wire _mesh_14_8_io_out_control_0_propagate;
	wire [4:0] _mesh_14_8_io_out_control_0_shift;
	wire [2:0] _mesh_14_8_io_out_id_0;
	wire _mesh_14_8_io_out_last_0;
	wire _mesh_14_8_io_out_valid_0;
	wire [31:0] _mesh_14_7_io_out_a_0;
	wire [31:0] _mesh_14_7_io_out_c_0;
	wire [31:0] _mesh_14_7_io_out_b_0;
	wire _mesh_14_7_io_out_control_0_dataflow;
	wire _mesh_14_7_io_out_control_0_propagate;
	wire [4:0] _mesh_14_7_io_out_control_0_shift;
	wire [2:0] _mesh_14_7_io_out_id_0;
	wire _mesh_14_7_io_out_last_0;
	wire _mesh_14_7_io_out_valid_0;
	wire [31:0] _mesh_14_6_io_out_a_0;
	wire [31:0] _mesh_14_6_io_out_c_0;
	wire [31:0] _mesh_14_6_io_out_b_0;
	wire _mesh_14_6_io_out_control_0_dataflow;
	wire _mesh_14_6_io_out_control_0_propagate;
	wire [4:0] _mesh_14_6_io_out_control_0_shift;
	wire [2:0] _mesh_14_6_io_out_id_0;
	wire _mesh_14_6_io_out_last_0;
	wire _mesh_14_6_io_out_valid_0;
	wire [31:0] _mesh_14_5_io_out_a_0;
	wire [31:0] _mesh_14_5_io_out_c_0;
	wire [31:0] _mesh_14_5_io_out_b_0;
	wire _mesh_14_5_io_out_control_0_dataflow;
	wire _mesh_14_5_io_out_control_0_propagate;
	wire [4:0] _mesh_14_5_io_out_control_0_shift;
	wire [2:0] _mesh_14_5_io_out_id_0;
	wire _mesh_14_5_io_out_last_0;
	wire _mesh_14_5_io_out_valid_0;
	wire [31:0] _mesh_14_4_io_out_a_0;
	wire [31:0] _mesh_14_4_io_out_c_0;
	wire [31:0] _mesh_14_4_io_out_b_0;
	wire _mesh_14_4_io_out_control_0_dataflow;
	wire _mesh_14_4_io_out_control_0_propagate;
	wire [4:0] _mesh_14_4_io_out_control_0_shift;
	wire [2:0] _mesh_14_4_io_out_id_0;
	wire _mesh_14_4_io_out_last_0;
	wire _mesh_14_4_io_out_valid_0;
	wire [31:0] _mesh_14_3_io_out_a_0;
	wire [31:0] _mesh_14_3_io_out_c_0;
	wire [31:0] _mesh_14_3_io_out_b_0;
	wire _mesh_14_3_io_out_control_0_dataflow;
	wire _mesh_14_3_io_out_control_0_propagate;
	wire [4:0] _mesh_14_3_io_out_control_0_shift;
	wire [2:0] _mesh_14_3_io_out_id_0;
	wire _mesh_14_3_io_out_last_0;
	wire _mesh_14_3_io_out_valid_0;
	wire [31:0] _mesh_14_2_io_out_a_0;
	wire [31:0] _mesh_14_2_io_out_c_0;
	wire [31:0] _mesh_14_2_io_out_b_0;
	wire _mesh_14_2_io_out_control_0_dataflow;
	wire _mesh_14_2_io_out_control_0_propagate;
	wire [4:0] _mesh_14_2_io_out_control_0_shift;
	wire [2:0] _mesh_14_2_io_out_id_0;
	wire _mesh_14_2_io_out_last_0;
	wire _mesh_14_2_io_out_valid_0;
	wire [31:0] _mesh_14_1_io_out_a_0;
	wire [31:0] _mesh_14_1_io_out_c_0;
	wire [31:0] _mesh_14_1_io_out_b_0;
	wire _mesh_14_1_io_out_control_0_dataflow;
	wire _mesh_14_1_io_out_control_0_propagate;
	wire [4:0] _mesh_14_1_io_out_control_0_shift;
	wire [2:0] _mesh_14_1_io_out_id_0;
	wire _mesh_14_1_io_out_last_0;
	wire _mesh_14_1_io_out_valid_0;
	wire [31:0] _mesh_14_0_io_out_a_0;
	wire [31:0] _mesh_14_0_io_out_c_0;
	wire [31:0] _mesh_14_0_io_out_b_0;
	wire _mesh_14_0_io_out_control_0_dataflow;
	wire _mesh_14_0_io_out_control_0_propagate;
	wire [4:0] _mesh_14_0_io_out_control_0_shift;
	wire [2:0] _mesh_14_0_io_out_id_0;
	wire _mesh_14_0_io_out_last_0;
	wire _mesh_14_0_io_out_valid_0;
	wire [31:0] _mesh_13_31_io_out_a_0;
	wire [31:0] _mesh_13_31_io_out_c_0;
	wire [31:0] _mesh_13_31_io_out_b_0;
	wire _mesh_13_31_io_out_control_0_dataflow;
	wire _mesh_13_31_io_out_control_0_propagate;
	wire [4:0] _mesh_13_31_io_out_control_0_shift;
	wire [2:0] _mesh_13_31_io_out_id_0;
	wire _mesh_13_31_io_out_last_0;
	wire _mesh_13_31_io_out_valid_0;
	wire [31:0] _mesh_13_30_io_out_a_0;
	wire [31:0] _mesh_13_30_io_out_c_0;
	wire [31:0] _mesh_13_30_io_out_b_0;
	wire _mesh_13_30_io_out_control_0_dataflow;
	wire _mesh_13_30_io_out_control_0_propagate;
	wire [4:0] _mesh_13_30_io_out_control_0_shift;
	wire [2:0] _mesh_13_30_io_out_id_0;
	wire _mesh_13_30_io_out_last_0;
	wire _mesh_13_30_io_out_valid_0;
	wire [31:0] _mesh_13_29_io_out_a_0;
	wire [31:0] _mesh_13_29_io_out_c_0;
	wire [31:0] _mesh_13_29_io_out_b_0;
	wire _mesh_13_29_io_out_control_0_dataflow;
	wire _mesh_13_29_io_out_control_0_propagate;
	wire [4:0] _mesh_13_29_io_out_control_0_shift;
	wire [2:0] _mesh_13_29_io_out_id_0;
	wire _mesh_13_29_io_out_last_0;
	wire _mesh_13_29_io_out_valid_0;
	wire [31:0] _mesh_13_28_io_out_a_0;
	wire [31:0] _mesh_13_28_io_out_c_0;
	wire [31:0] _mesh_13_28_io_out_b_0;
	wire _mesh_13_28_io_out_control_0_dataflow;
	wire _mesh_13_28_io_out_control_0_propagate;
	wire [4:0] _mesh_13_28_io_out_control_0_shift;
	wire [2:0] _mesh_13_28_io_out_id_0;
	wire _mesh_13_28_io_out_last_0;
	wire _mesh_13_28_io_out_valid_0;
	wire [31:0] _mesh_13_27_io_out_a_0;
	wire [31:0] _mesh_13_27_io_out_c_0;
	wire [31:0] _mesh_13_27_io_out_b_0;
	wire _mesh_13_27_io_out_control_0_dataflow;
	wire _mesh_13_27_io_out_control_0_propagate;
	wire [4:0] _mesh_13_27_io_out_control_0_shift;
	wire [2:0] _mesh_13_27_io_out_id_0;
	wire _mesh_13_27_io_out_last_0;
	wire _mesh_13_27_io_out_valid_0;
	wire [31:0] _mesh_13_26_io_out_a_0;
	wire [31:0] _mesh_13_26_io_out_c_0;
	wire [31:0] _mesh_13_26_io_out_b_0;
	wire _mesh_13_26_io_out_control_0_dataflow;
	wire _mesh_13_26_io_out_control_0_propagate;
	wire [4:0] _mesh_13_26_io_out_control_0_shift;
	wire [2:0] _mesh_13_26_io_out_id_0;
	wire _mesh_13_26_io_out_last_0;
	wire _mesh_13_26_io_out_valid_0;
	wire [31:0] _mesh_13_25_io_out_a_0;
	wire [31:0] _mesh_13_25_io_out_c_0;
	wire [31:0] _mesh_13_25_io_out_b_0;
	wire _mesh_13_25_io_out_control_0_dataflow;
	wire _mesh_13_25_io_out_control_0_propagate;
	wire [4:0] _mesh_13_25_io_out_control_0_shift;
	wire [2:0] _mesh_13_25_io_out_id_0;
	wire _mesh_13_25_io_out_last_0;
	wire _mesh_13_25_io_out_valid_0;
	wire [31:0] _mesh_13_24_io_out_a_0;
	wire [31:0] _mesh_13_24_io_out_c_0;
	wire [31:0] _mesh_13_24_io_out_b_0;
	wire _mesh_13_24_io_out_control_0_dataflow;
	wire _mesh_13_24_io_out_control_0_propagate;
	wire [4:0] _mesh_13_24_io_out_control_0_shift;
	wire [2:0] _mesh_13_24_io_out_id_0;
	wire _mesh_13_24_io_out_last_0;
	wire _mesh_13_24_io_out_valid_0;
	wire [31:0] _mesh_13_23_io_out_a_0;
	wire [31:0] _mesh_13_23_io_out_c_0;
	wire [31:0] _mesh_13_23_io_out_b_0;
	wire _mesh_13_23_io_out_control_0_dataflow;
	wire _mesh_13_23_io_out_control_0_propagate;
	wire [4:0] _mesh_13_23_io_out_control_0_shift;
	wire [2:0] _mesh_13_23_io_out_id_0;
	wire _mesh_13_23_io_out_last_0;
	wire _mesh_13_23_io_out_valid_0;
	wire [31:0] _mesh_13_22_io_out_a_0;
	wire [31:0] _mesh_13_22_io_out_c_0;
	wire [31:0] _mesh_13_22_io_out_b_0;
	wire _mesh_13_22_io_out_control_0_dataflow;
	wire _mesh_13_22_io_out_control_0_propagate;
	wire [4:0] _mesh_13_22_io_out_control_0_shift;
	wire [2:0] _mesh_13_22_io_out_id_0;
	wire _mesh_13_22_io_out_last_0;
	wire _mesh_13_22_io_out_valid_0;
	wire [31:0] _mesh_13_21_io_out_a_0;
	wire [31:0] _mesh_13_21_io_out_c_0;
	wire [31:0] _mesh_13_21_io_out_b_0;
	wire _mesh_13_21_io_out_control_0_dataflow;
	wire _mesh_13_21_io_out_control_0_propagate;
	wire [4:0] _mesh_13_21_io_out_control_0_shift;
	wire [2:0] _mesh_13_21_io_out_id_0;
	wire _mesh_13_21_io_out_last_0;
	wire _mesh_13_21_io_out_valid_0;
	wire [31:0] _mesh_13_20_io_out_a_0;
	wire [31:0] _mesh_13_20_io_out_c_0;
	wire [31:0] _mesh_13_20_io_out_b_0;
	wire _mesh_13_20_io_out_control_0_dataflow;
	wire _mesh_13_20_io_out_control_0_propagate;
	wire [4:0] _mesh_13_20_io_out_control_0_shift;
	wire [2:0] _mesh_13_20_io_out_id_0;
	wire _mesh_13_20_io_out_last_0;
	wire _mesh_13_20_io_out_valid_0;
	wire [31:0] _mesh_13_19_io_out_a_0;
	wire [31:0] _mesh_13_19_io_out_c_0;
	wire [31:0] _mesh_13_19_io_out_b_0;
	wire _mesh_13_19_io_out_control_0_dataflow;
	wire _mesh_13_19_io_out_control_0_propagate;
	wire [4:0] _mesh_13_19_io_out_control_0_shift;
	wire [2:0] _mesh_13_19_io_out_id_0;
	wire _mesh_13_19_io_out_last_0;
	wire _mesh_13_19_io_out_valid_0;
	wire [31:0] _mesh_13_18_io_out_a_0;
	wire [31:0] _mesh_13_18_io_out_c_0;
	wire [31:0] _mesh_13_18_io_out_b_0;
	wire _mesh_13_18_io_out_control_0_dataflow;
	wire _mesh_13_18_io_out_control_0_propagate;
	wire [4:0] _mesh_13_18_io_out_control_0_shift;
	wire [2:0] _mesh_13_18_io_out_id_0;
	wire _mesh_13_18_io_out_last_0;
	wire _mesh_13_18_io_out_valid_0;
	wire [31:0] _mesh_13_17_io_out_a_0;
	wire [31:0] _mesh_13_17_io_out_c_0;
	wire [31:0] _mesh_13_17_io_out_b_0;
	wire _mesh_13_17_io_out_control_0_dataflow;
	wire _mesh_13_17_io_out_control_0_propagate;
	wire [4:0] _mesh_13_17_io_out_control_0_shift;
	wire [2:0] _mesh_13_17_io_out_id_0;
	wire _mesh_13_17_io_out_last_0;
	wire _mesh_13_17_io_out_valid_0;
	wire [31:0] _mesh_13_16_io_out_a_0;
	wire [31:0] _mesh_13_16_io_out_c_0;
	wire [31:0] _mesh_13_16_io_out_b_0;
	wire _mesh_13_16_io_out_control_0_dataflow;
	wire _mesh_13_16_io_out_control_0_propagate;
	wire [4:0] _mesh_13_16_io_out_control_0_shift;
	wire [2:0] _mesh_13_16_io_out_id_0;
	wire _mesh_13_16_io_out_last_0;
	wire _mesh_13_16_io_out_valid_0;
	wire [31:0] _mesh_13_15_io_out_a_0;
	wire [31:0] _mesh_13_15_io_out_c_0;
	wire [31:0] _mesh_13_15_io_out_b_0;
	wire _mesh_13_15_io_out_control_0_dataflow;
	wire _mesh_13_15_io_out_control_0_propagate;
	wire [4:0] _mesh_13_15_io_out_control_0_shift;
	wire [2:0] _mesh_13_15_io_out_id_0;
	wire _mesh_13_15_io_out_last_0;
	wire _mesh_13_15_io_out_valid_0;
	wire [31:0] _mesh_13_14_io_out_a_0;
	wire [31:0] _mesh_13_14_io_out_c_0;
	wire [31:0] _mesh_13_14_io_out_b_0;
	wire _mesh_13_14_io_out_control_0_dataflow;
	wire _mesh_13_14_io_out_control_0_propagate;
	wire [4:0] _mesh_13_14_io_out_control_0_shift;
	wire [2:0] _mesh_13_14_io_out_id_0;
	wire _mesh_13_14_io_out_last_0;
	wire _mesh_13_14_io_out_valid_0;
	wire [31:0] _mesh_13_13_io_out_a_0;
	wire [31:0] _mesh_13_13_io_out_c_0;
	wire [31:0] _mesh_13_13_io_out_b_0;
	wire _mesh_13_13_io_out_control_0_dataflow;
	wire _mesh_13_13_io_out_control_0_propagate;
	wire [4:0] _mesh_13_13_io_out_control_0_shift;
	wire [2:0] _mesh_13_13_io_out_id_0;
	wire _mesh_13_13_io_out_last_0;
	wire _mesh_13_13_io_out_valid_0;
	wire [31:0] _mesh_13_12_io_out_a_0;
	wire [31:0] _mesh_13_12_io_out_c_0;
	wire [31:0] _mesh_13_12_io_out_b_0;
	wire _mesh_13_12_io_out_control_0_dataflow;
	wire _mesh_13_12_io_out_control_0_propagate;
	wire [4:0] _mesh_13_12_io_out_control_0_shift;
	wire [2:0] _mesh_13_12_io_out_id_0;
	wire _mesh_13_12_io_out_last_0;
	wire _mesh_13_12_io_out_valid_0;
	wire [31:0] _mesh_13_11_io_out_a_0;
	wire [31:0] _mesh_13_11_io_out_c_0;
	wire [31:0] _mesh_13_11_io_out_b_0;
	wire _mesh_13_11_io_out_control_0_dataflow;
	wire _mesh_13_11_io_out_control_0_propagate;
	wire [4:0] _mesh_13_11_io_out_control_0_shift;
	wire [2:0] _mesh_13_11_io_out_id_0;
	wire _mesh_13_11_io_out_last_0;
	wire _mesh_13_11_io_out_valid_0;
	wire [31:0] _mesh_13_10_io_out_a_0;
	wire [31:0] _mesh_13_10_io_out_c_0;
	wire [31:0] _mesh_13_10_io_out_b_0;
	wire _mesh_13_10_io_out_control_0_dataflow;
	wire _mesh_13_10_io_out_control_0_propagate;
	wire [4:0] _mesh_13_10_io_out_control_0_shift;
	wire [2:0] _mesh_13_10_io_out_id_0;
	wire _mesh_13_10_io_out_last_0;
	wire _mesh_13_10_io_out_valid_0;
	wire [31:0] _mesh_13_9_io_out_a_0;
	wire [31:0] _mesh_13_9_io_out_c_0;
	wire [31:0] _mesh_13_9_io_out_b_0;
	wire _mesh_13_9_io_out_control_0_dataflow;
	wire _mesh_13_9_io_out_control_0_propagate;
	wire [4:0] _mesh_13_9_io_out_control_0_shift;
	wire [2:0] _mesh_13_9_io_out_id_0;
	wire _mesh_13_9_io_out_last_0;
	wire _mesh_13_9_io_out_valid_0;
	wire [31:0] _mesh_13_8_io_out_a_0;
	wire [31:0] _mesh_13_8_io_out_c_0;
	wire [31:0] _mesh_13_8_io_out_b_0;
	wire _mesh_13_8_io_out_control_0_dataflow;
	wire _mesh_13_8_io_out_control_0_propagate;
	wire [4:0] _mesh_13_8_io_out_control_0_shift;
	wire [2:0] _mesh_13_8_io_out_id_0;
	wire _mesh_13_8_io_out_last_0;
	wire _mesh_13_8_io_out_valid_0;
	wire [31:0] _mesh_13_7_io_out_a_0;
	wire [31:0] _mesh_13_7_io_out_c_0;
	wire [31:0] _mesh_13_7_io_out_b_0;
	wire _mesh_13_7_io_out_control_0_dataflow;
	wire _mesh_13_7_io_out_control_0_propagate;
	wire [4:0] _mesh_13_7_io_out_control_0_shift;
	wire [2:0] _mesh_13_7_io_out_id_0;
	wire _mesh_13_7_io_out_last_0;
	wire _mesh_13_7_io_out_valid_0;
	wire [31:0] _mesh_13_6_io_out_a_0;
	wire [31:0] _mesh_13_6_io_out_c_0;
	wire [31:0] _mesh_13_6_io_out_b_0;
	wire _mesh_13_6_io_out_control_0_dataflow;
	wire _mesh_13_6_io_out_control_0_propagate;
	wire [4:0] _mesh_13_6_io_out_control_0_shift;
	wire [2:0] _mesh_13_6_io_out_id_0;
	wire _mesh_13_6_io_out_last_0;
	wire _mesh_13_6_io_out_valid_0;
	wire [31:0] _mesh_13_5_io_out_a_0;
	wire [31:0] _mesh_13_5_io_out_c_0;
	wire [31:0] _mesh_13_5_io_out_b_0;
	wire _mesh_13_5_io_out_control_0_dataflow;
	wire _mesh_13_5_io_out_control_0_propagate;
	wire [4:0] _mesh_13_5_io_out_control_0_shift;
	wire [2:0] _mesh_13_5_io_out_id_0;
	wire _mesh_13_5_io_out_last_0;
	wire _mesh_13_5_io_out_valid_0;
	wire [31:0] _mesh_13_4_io_out_a_0;
	wire [31:0] _mesh_13_4_io_out_c_0;
	wire [31:0] _mesh_13_4_io_out_b_0;
	wire _mesh_13_4_io_out_control_0_dataflow;
	wire _mesh_13_4_io_out_control_0_propagate;
	wire [4:0] _mesh_13_4_io_out_control_0_shift;
	wire [2:0] _mesh_13_4_io_out_id_0;
	wire _mesh_13_4_io_out_last_0;
	wire _mesh_13_4_io_out_valid_0;
	wire [31:0] _mesh_13_3_io_out_a_0;
	wire [31:0] _mesh_13_3_io_out_c_0;
	wire [31:0] _mesh_13_3_io_out_b_0;
	wire _mesh_13_3_io_out_control_0_dataflow;
	wire _mesh_13_3_io_out_control_0_propagate;
	wire [4:0] _mesh_13_3_io_out_control_0_shift;
	wire [2:0] _mesh_13_3_io_out_id_0;
	wire _mesh_13_3_io_out_last_0;
	wire _mesh_13_3_io_out_valid_0;
	wire [31:0] _mesh_13_2_io_out_a_0;
	wire [31:0] _mesh_13_2_io_out_c_0;
	wire [31:0] _mesh_13_2_io_out_b_0;
	wire _mesh_13_2_io_out_control_0_dataflow;
	wire _mesh_13_2_io_out_control_0_propagate;
	wire [4:0] _mesh_13_2_io_out_control_0_shift;
	wire [2:0] _mesh_13_2_io_out_id_0;
	wire _mesh_13_2_io_out_last_0;
	wire _mesh_13_2_io_out_valid_0;
	wire [31:0] _mesh_13_1_io_out_a_0;
	wire [31:0] _mesh_13_1_io_out_c_0;
	wire [31:0] _mesh_13_1_io_out_b_0;
	wire _mesh_13_1_io_out_control_0_dataflow;
	wire _mesh_13_1_io_out_control_0_propagate;
	wire [4:0] _mesh_13_1_io_out_control_0_shift;
	wire [2:0] _mesh_13_1_io_out_id_0;
	wire _mesh_13_1_io_out_last_0;
	wire _mesh_13_1_io_out_valid_0;
	wire [31:0] _mesh_13_0_io_out_a_0;
	wire [31:0] _mesh_13_0_io_out_c_0;
	wire [31:0] _mesh_13_0_io_out_b_0;
	wire _mesh_13_0_io_out_control_0_dataflow;
	wire _mesh_13_0_io_out_control_0_propagate;
	wire [4:0] _mesh_13_0_io_out_control_0_shift;
	wire [2:0] _mesh_13_0_io_out_id_0;
	wire _mesh_13_0_io_out_last_0;
	wire _mesh_13_0_io_out_valid_0;
	wire [31:0] _mesh_12_31_io_out_a_0;
	wire [31:0] _mesh_12_31_io_out_c_0;
	wire [31:0] _mesh_12_31_io_out_b_0;
	wire _mesh_12_31_io_out_control_0_dataflow;
	wire _mesh_12_31_io_out_control_0_propagate;
	wire [4:0] _mesh_12_31_io_out_control_0_shift;
	wire [2:0] _mesh_12_31_io_out_id_0;
	wire _mesh_12_31_io_out_last_0;
	wire _mesh_12_31_io_out_valid_0;
	wire [31:0] _mesh_12_30_io_out_a_0;
	wire [31:0] _mesh_12_30_io_out_c_0;
	wire [31:0] _mesh_12_30_io_out_b_0;
	wire _mesh_12_30_io_out_control_0_dataflow;
	wire _mesh_12_30_io_out_control_0_propagate;
	wire [4:0] _mesh_12_30_io_out_control_0_shift;
	wire [2:0] _mesh_12_30_io_out_id_0;
	wire _mesh_12_30_io_out_last_0;
	wire _mesh_12_30_io_out_valid_0;
	wire [31:0] _mesh_12_29_io_out_a_0;
	wire [31:0] _mesh_12_29_io_out_c_0;
	wire [31:0] _mesh_12_29_io_out_b_0;
	wire _mesh_12_29_io_out_control_0_dataflow;
	wire _mesh_12_29_io_out_control_0_propagate;
	wire [4:0] _mesh_12_29_io_out_control_0_shift;
	wire [2:0] _mesh_12_29_io_out_id_0;
	wire _mesh_12_29_io_out_last_0;
	wire _mesh_12_29_io_out_valid_0;
	wire [31:0] _mesh_12_28_io_out_a_0;
	wire [31:0] _mesh_12_28_io_out_c_0;
	wire [31:0] _mesh_12_28_io_out_b_0;
	wire _mesh_12_28_io_out_control_0_dataflow;
	wire _mesh_12_28_io_out_control_0_propagate;
	wire [4:0] _mesh_12_28_io_out_control_0_shift;
	wire [2:0] _mesh_12_28_io_out_id_0;
	wire _mesh_12_28_io_out_last_0;
	wire _mesh_12_28_io_out_valid_0;
	wire [31:0] _mesh_12_27_io_out_a_0;
	wire [31:0] _mesh_12_27_io_out_c_0;
	wire [31:0] _mesh_12_27_io_out_b_0;
	wire _mesh_12_27_io_out_control_0_dataflow;
	wire _mesh_12_27_io_out_control_0_propagate;
	wire [4:0] _mesh_12_27_io_out_control_0_shift;
	wire [2:0] _mesh_12_27_io_out_id_0;
	wire _mesh_12_27_io_out_last_0;
	wire _mesh_12_27_io_out_valid_0;
	wire [31:0] _mesh_12_26_io_out_a_0;
	wire [31:0] _mesh_12_26_io_out_c_0;
	wire [31:0] _mesh_12_26_io_out_b_0;
	wire _mesh_12_26_io_out_control_0_dataflow;
	wire _mesh_12_26_io_out_control_0_propagate;
	wire [4:0] _mesh_12_26_io_out_control_0_shift;
	wire [2:0] _mesh_12_26_io_out_id_0;
	wire _mesh_12_26_io_out_last_0;
	wire _mesh_12_26_io_out_valid_0;
	wire [31:0] _mesh_12_25_io_out_a_0;
	wire [31:0] _mesh_12_25_io_out_c_0;
	wire [31:0] _mesh_12_25_io_out_b_0;
	wire _mesh_12_25_io_out_control_0_dataflow;
	wire _mesh_12_25_io_out_control_0_propagate;
	wire [4:0] _mesh_12_25_io_out_control_0_shift;
	wire [2:0] _mesh_12_25_io_out_id_0;
	wire _mesh_12_25_io_out_last_0;
	wire _mesh_12_25_io_out_valid_0;
	wire [31:0] _mesh_12_24_io_out_a_0;
	wire [31:0] _mesh_12_24_io_out_c_0;
	wire [31:0] _mesh_12_24_io_out_b_0;
	wire _mesh_12_24_io_out_control_0_dataflow;
	wire _mesh_12_24_io_out_control_0_propagate;
	wire [4:0] _mesh_12_24_io_out_control_0_shift;
	wire [2:0] _mesh_12_24_io_out_id_0;
	wire _mesh_12_24_io_out_last_0;
	wire _mesh_12_24_io_out_valid_0;
	wire [31:0] _mesh_12_23_io_out_a_0;
	wire [31:0] _mesh_12_23_io_out_c_0;
	wire [31:0] _mesh_12_23_io_out_b_0;
	wire _mesh_12_23_io_out_control_0_dataflow;
	wire _mesh_12_23_io_out_control_0_propagate;
	wire [4:0] _mesh_12_23_io_out_control_0_shift;
	wire [2:0] _mesh_12_23_io_out_id_0;
	wire _mesh_12_23_io_out_last_0;
	wire _mesh_12_23_io_out_valid_0;
	wire [31:0] _mesh_12_22_io_out_a_0;
	wire [31:0] _mesh_12_22_io_out_c_0;
	wire [31:0] _mesh_12_22_io_out_b_0;
	wire _mesh_12_22_io_out_control_0_dataflow;
	wire _mesh_12_22_io_out_control_0_propagate;
	wire [4:0] _mesh_12_22_io_out_control_0_shift;
	wire [2:0] _mesh_12_22_io_out_id_0;
	wire _mesh_12_22_io_out_last_0;
	wire _mesh_12_22_io_out_valid_0;
	wire [31:0] _mesh_12_21_io_out_a_0;
	wire [31:0] _mesh_12_21_io_out_c_0;
	wire [31:0] _mesh_12_21_io_out_b_0;
	wire _mesh_12_21_io_out_control_0_dataflow;
	wire _mesh_12_21_io_out_control_0_propagate;
	wire [4:0] _mesh_12_21_io_out_control_0_shift;
	wire [2:0] _mesh_12_21_io_out_id_0;
	wire _mesh_12_21_io_out_last_0;
	wire _mesh_12_21_io_out_valid_0;
	wire [31:0] _mesh_12_20_io_out_a_0;
	wire [31:0] _mesh_12_20_io_out_c_0;
	wire [31:0] _mesh_12_20_io_out_b_0;
	wire _mesh_12_20_io_out_control_0_dataflow;
	wire _mesh_12_20_io_out_control_0_propagate;
	wire [4:0] _mesh_12_20_io_out_control_0_shift;
	wire [2:0] _mesh_12_20_io_out_id_0;
	wire _mesh_12_20_io_out_last_0;
	wire _mesh_12_20_io_out_valid_0;
	wire [31:0] _mesh_12_19_io_out_a_0;
	wire [31:0] _mesh_12_19_io_out_c_0;
	wire [31:0] _mesh_12_19_io_out_b_0;
	wire _mesh_12_19_io_out_control_0_dataflow;
	wire _mesh_12_19_io_out_control_0_propagate;
	wire [4:0] _mesh_12_19_io_out_control_0_shift;
	wire [2:0] _mesh_12_19_io_out_id_0;
	wire _mesh_12_19_io_out_last_0;
	wire _mesh_12_19_io_out_valid_0;
	wire [31:0] _mesh_12_18_io_out_a_0;
	wire [31:0] _mesh_12_18_io_out_c_0;
	wire [31:0] _mesh_12_18_io_out_b_0;
	wire _mesh_12_18_io_out_control_0_dataflow;
	wire _mesh_12_18_io_out_control_0_propagate;
	wire [4:0] _mesh_12_18_io_out_control_0_shift;
	wire [2:0] _mesh_12_18_io_out_id_0;
	wire _mesh_12_18_io_out_last_0;
	wire _mesh_12_18_io_out_valid_0;
	wire [31:0] _mesh_12_17_io_out_a_0;
	wire [31:0] _mesh_12_17_io_out_c_0;
	wire [31:0] _mesh_12_17_io_out_b_0;
	wire _mesh_12_17_io_out_control_0_dataflow;
	wire _mesh_12_17_io_out_control_0_propagate;
	wire [4:0] _mesh_12_17_io_out_control_0_shift;
	wire [2:0] _mesh_12_17_io_out_id_0;
	wire _mesh_12_17_io_out_last_0;
	wire _mesh_12_17_io_out_valid_0;
	wire [31:0] _mesh_12_16_io_out_a_0;
	wire [31:0] _mesh_12_16_io_out_c_0;
	wire [31:0] _mesh_12_16_io_out_b_0;
	wire _mesh_12_16_io_out_control_0_dataflow;
	wire _mesh_12_16_io_out_control_0_propagate;
	wire [4:0] _mesh_12_16_io_out_control_0_shift;
	wire [2:0] _mesh_12_16_io_out_id_0;
	wire _mesh_12_16_io_out_last_0;
	wire _mesh_12_16_io_out_valid_0;
	wire [31:0] _mesh_12_15_io_out_a_0;
	wire [31:0] _mesh_12_15_io_out_c_0;
	wire [31:0] _mesh_12_15_io_out_b_0;
	wire _mesh_12_15_io_out_control_0_dataflow;
	wire _mesh_12_15_io_out_control_0_propagate;
	wire [4:0] _mesh_12_15_io_out_control_0_shift;
	wire [2:0] _mesh_12_15_io_out_id_0;
	wire _mesh_12_15_io_out_last_0;
	wire _mesh_12_15_io_out_valid_0;
	wire [31:0] _mesh_12_14_io_out_a_0;
	wire [31:0] _mesh_12_14_io_out_c_0;
	wire [31:0] _mesh_12_14_io_out_b_0;
	wire _mesh_12_14_io_out_control_0_dataflow;
	wire _mesh_12_14_io_out_control_0_propagate;
	wire [4:0] _mesh_12_14_io_out_control_0_shift;
	wire [2:0] _mesh_12_14_io_out_id_0;
	wire _mesh_12_14_io_out_last_0;
	wire _mesh_12_14_io_out_valid_0;
	wire [31:0] _mesh_12_13_io_out_a_0;
	wire [31:0] _mesh_12_13_io_out_c_0;
	wire [31:0] _mesh_12_13_io_out_b_0;
	wire _mesh_12_13_io_out_control_0_dataflow;
	wire _mesh_12_13_io_out_control_0_propagate;
	wire [4:0] _mesh_12_13_io_out_control_0_shift;
	wire [2:0] _mesh_12_13_io_out_id_0;
	wire _mesh_12_13_io_out_last_0;
	wire _mesh_12_13_io_out_valid_0;
	wire [31:0] _mesh_12_12_io_out_a_0;
	wire [31:0] _mesh_12_12_io_out_c_0;
	wire [31:0] _mesh_12_12_io_out_b_0;
	wire _mesh_12_12_io_out_control_0_dataflow;
	wire _mesh_12_12_io_out_control_0_propagate;
	wire [4:0] _mesh_12_12_io_out_control_0_shift;
	wire [2:0] _mesh_12_12_io_out_id_0;
	wire _mesh_12_12_io_out_last_0;
	wire _mesh_12_12_io_out_valid_0;
	wire [31:0] _mesh_12_11_io_out_a_0;
	wire [31:0] _mesh_12_11_io_out_c_0;
	wire [31:0] _mesh_12_11_io_out_b_0;
	wire _mesh_12_11_io_out_control_0_dataflow;
	wire _mesh_12_11_io_out_control_0_propagate;
	wire [4:0] _mesh_12_11_io_out_control_0_shift;
	wire [2:0] _mesh_12_11_io_out_id_0;
	wire _mesh_12_11_io_out_last_0;
	wire _mesh_12_11_io_out_valid_0;
	wire [31:0] _mesh_12_10_io_out_a_0;
	wire [31:0] _mesh_12_10_io_out_c_0;
	wire [31:0] _mesh_12_10_io_out_b_0;
	wire _mesh_12_10_io_out_control_0_dataflow;
	wire _mesh_12_10_io_out_control_0_propagate;
	wire [4:0] _mesh_12_10_io_out_control_0_shift;
	wire [2:0] _mesh_12_10_io_out_id_0;
	wire _mesh_12_10_io_out_last_0;
	wire _mesh_12_10_io_out_valid_0;
	wire [31:0] _mesh_12_9_io_out_a_0;
	wire [31:0] _mesh_12_9_io_out_c_0;
	wire [31:0] _mesh_12_9_io_out_b_0;
	wire _mesh_12_9_io_out_control_0_dataflow;
	wire _mesh_12_9_io_out_control_0_propagate;
	wire [4:0] _mesh_12_9_io_out_control_0_shift;
	wire [2:0] _mesh_12_9_io_out_id_0;
	wire _mesh_12_9_io_out_last_0;
	wire _mesh_12_9_io_out_valid_0;
	wire [31:0] _mesh_12_8_io_out_a_0;
	wire [31:0] _mesh_12_8_io_out_c_0;
	wire [31:0] _mesh_12_8_io_out_b_0;
	wire _mesh_12_8_io_out_control_0_dataflow;
	wire _mesh_12_8_io_out_control_0_propagate;
	wire [4:0] _mesh_12_8_io_out_control_0_shift;
	wire [2:0] _mesh_12_8_io_out_id_0;
	wire _mesh_12_8_io_out_last_0;
	wire _mesh_12_8_io_out_valid_0;
	wire [31:0] _mesh_12_7_io_out_a_0;
	wire [31:0] _mesh_12_7_io_out_c_0;
	wire [31:0] _mesh_12_7_io_out_b_0;
	wire _mesh_12_7_io_out_control_0_dataflow;
	wire _mesh_12_7_io_out_control_0_propagate;
	wire [4:0] _mesh_12_7_io_out_control_0_shift;
	wire [2:0] _mesh_12_7_io_out_id_0;
	wire _mesh_12_7_io_out_last_0;
	wire _mesh_12_7_io_out_valid_0;
	wire [31:0] _mesh_12_6_io_out_a_0;
	wire [31:0] _mesh_12_6_io_out_c_0;
	wire [31:0] _mesh_12_6_io_out_b_0;
	wire _mesh_12_6_io_out_control_0_dataflow;
	wire _mesh_12_6_io_out_control_0_propagate;
	wire [4:0] _mesh_12_6_io_out_control_0_shift;
	wire [2:0] _mesh_12_6_io_out_id_0;
	wire _mesh_12_6_io_out_last_0;
	wire _mesh_12_6_io_out_valid_0;
	wire [31:0] _mesh_12_5_io_out_a_0;
	wire [31:0] _mesh_12_5_io_out_c_0;
	wire [31:0] _mesh_12_5_io_out_b_0;
	wire _mesh_12_5_io_out_control_0_dataflow;
	wire _mesh_12_5_io_out_control_0_propagate;
	wire [4:0] _mesh_12_5_io_out_control_0_shift;
	wire [2:0] _mesh_12_5_io_out_id_0;
	wire _mesh_12_5_io_out_last_0;
	wire _mesh_12_5_io_out_valid_0;
	wire [31:0] _mesh_12_4_io_out_a_0;
	wire [31:0] _mesh_12_4_io_out_c_0;
	wire [31:0] _mesh_12_4_io_out_b_0;
	wire _mesh_12_4_io_out_control_0_dataflow;
	wire _mesh_12_4_io_out_control_0_propagate;
	wire [4:0] _mesh_12_4_io_out_control_0_shift;
	wire [2:0] _mesh_12_4_io_out_id_0;
	wire _mesh_12_4_io_out_last_0;
	wire _mesh_12_4_io_out_valid_0;
	wire [31:0] _mesh_12_3_io_out_a_0;
	wire [31:0] _mesh_12_3_io_out_c_0;
	wire [31:0] _mesh_12_3_io_out_b_0;
	wire _mesh_12_3_io_out_control_0_dataflow;
	wire _mesh_12_3_io_out_control_0_propagate;
	wire [4:0] _mesh_12_3_io_out_control_0_shift;
	wire [2:0] _mesh_12_3_io_out_id_0;
	wire _mesh_12_3_io_out_last_0;
	wire _mesh_12_3_io_out_valid_0;
	wire [31:0] _mesh_12_2_io_out_a_0;
	wire [31:0] _mesh_12_2_io_out_c_0;
	wire [31:0] _mesh_12_2_io_out_b_0;
	wire _mesh_12_2_io_out_control_0_dataflow;
	wire _mesh_12_2_io_out_control_0_propagate;
	wire [4:0] _mesh_12_2_io_out_control_0_shift;
	wire [2:0] _mesh_12_2_io_out_id_0;
	wire _mesh_12_2_io_out_last_0;
	wire _mesh_12_2_io_out_valid_0;
	wire [31:0] _mesh_12_1_io_out_a_0;
	wire [31:0] _mesh_12_1_io_out_c_0;
	wire [31:0] _mesh_12_1_io_out_b_0;
	wire _mesh_12_1_io_out_control_0_dataflow;
	wire _mesh_12_1_io_out_control_0_propagate;
	wire [4:0] _mesh_12_1_io_out_control_0_shift;
	wire [2:0] _mesh_12_1_io_out_id_0;
	wire _mesh_12_1_io_out_last_0;
	wire _mesh_12_1_io_out_valid_0;
	wire [31:0] _mesh_12_0_io_out_a_0;
	wire [31:0] _mesh_12_0_io_out_c_0;
	wire [31:0] _mesh_12_0_io_out_b_0;
	wire _mesh_12_0_io_out_control_0_dataflow;
	wire _mesh_12_0_io_out_control_0_propagate;
	wire [4:0] _mesh_12_0_io_out_control_0_shift;
	wire [2:0] _mesh_12_0_io_out_id_0;
	wire _mesh_12_0_io_out_last_0;
	wire _mesh_12_0_io_out_valid_0;
	wire [31:0] _mesh_11_31_io_out_a_0;
	wire [31:0] _mesh_11_31_io_out_c_0;
	wire [31:0] _mesh_11_31_io_out_b_0;
	wire _mesh_11_31_io_out_control_0_dataflow;
	wire _mesh_11_31_io_out_control_0_propagate;
	wire [4:0] _mesh_11_31_io_out_control_0_shift;
	wire [2:0] _mesh_11_31_io_out_id_0;
	wire _mesh_11_31_io_out_last_0;
	wire _mesh_11_31_io_out_valid_0;
	wire [31:0] _mesh_11_30_io_out_a_0;
	wire [31:0] _mesh_11_30_io_out_c_0;
	wire [31:0] _mesh_11_30_io_out_b_0;
	wire _mesh_11_30_io_out_control_0_dataflow;
	wire _mesh_11_30_io_out_control_0_propagate;
	wire [4:0] _mesh_11_30_io_out_control_0_shift;
	wire [2:0] _mesh_11_30_io_out_id_0;
	wire _mesh_11_30_io_out_last_0;
	wire _mesh_11_30_io_out_valid_0;
	wire [31:0] _mesh_11_29_io_out_a_0;
	wire [31:0] _mesh_11_29_io_out_c_0;
	wire [31:0] _mesh_11_29_io_out_b_0;
	wire _mesh_11_29_io_out_control_0_dataflow;
	wire _mesh_11_29_io_out_control_0_propagate;
	wire [4:0] _mesh_11_29_io_out_control_0_shift;
	wire [2:0] _mesh_11_29_io_out_id_0;
	wire _mesh_11_29_io_out_last_0;
	wire _mesh_11_29_io_out_valid_0;
	wire [31:0] _mesh_11_28_io_out_a_0;
	wire [31:0] _mesh_11_28_io_out_c_0;
	wire [31:0] _mesh_11_28_io_out_b_0;
	wire _mesh_11_28_io_out_control_0_dataflow;
	wire _mesh_11_28_io_out_control_0_propagate;
	wire [4:0] _mesh_11_28_io_out_control_0_shift;
	wire [2:0] _mesh_11_28_io_out_id_0;
	wire _mesh_11_28_io_out_last_0;
	wire _mesh_11_28_io_out_valid_0;
	wire [31:0] _mesh_11_27_io_out_a_0;
	wire [31:0] _mesh_11_27_io_out_c_0;
	wire [31:0] _mesh_11_27_io_out_b_0;
	wire _mesh_11_27_io_out_control_0_dataflow;
	wire _mesh_11_27_io_out_control_0_propagate;
	wire [4:0] _mesh_11_27_io_out_control_0_shift;
	wire [2:0] _mesh_11_27_io_out_id_0;
	wire _mesh_11_27_io_out_last_0;
	wire _mesh_11_27_io_out_valid_0;
	wire [31:0] _mesh_11_26_io_out_a_0;
	wire [31:0] _mesh_11_26_io_out_c_0;
	wire [31:0] _mesh_11_26_io_out_b_0;
	wire _mesh_11_26_io_out_control_0_dataflow;
	wire _mesh_11_26_io_out_control_0_propagate;
	wire [4:0] _mesh_11_26_io_out_control_0_shift;
	wire [2:0] _mesh_11_26_io_out_id_0;
	wire _mesh_11_26_io_out_last_0;
	wire _mesh_11_26_io_out_valid_0;
	wire [31:0] _mesh_11_25_io_out_a_0;
	wire [31:0] _mesh_11_25_io_out_c_0;
	wire [31:0] _mesh_11_25_io_out_b_0;
	wire _mesh_11_25_io_out_control_0_dataflow;
	wire _mesh_11_25_io_out_control_0_propagate;
	wire [4:0] _mesh_11_25_io_out_control_0_shift;
	wire [2:0] _mesh_11_25_io_out_id_0;
	wire _mesh_11_25_io_out_last_0;
	wire _mesh_11_25_io_out_valid_0;
	wire [31:0] _mesh_11_24_io_out_a_0;
	wire [31:0] _mesh_11_24_io_out_c_0;
	wire [31:0] _mesh_11_24_io_out_b_0;
	wire _mesh_11_24_io_out_control_0_dataflow;
	wire _mesh_11_24_io_out_control_0_propagate;
	wire [4:0] _mesh_11_24_io_out_control_0_shift;
	wire [2:0] _mesh_11_24_io_out_id_0;
	wire _mesh_11_24_io_out_last_0;
	wire _mesh_11_24_io_out_valid_0;
	wire [31:0] _mesh_11_23_io_out_a_0;
	wire [31:0] _mesh_11_23_io_out_c_0;
	wire [31:0] _mesh_11_23_io_out_b_0;
	wire _mesh_11_23_io_out_control_0_dataflow;
	wire _mesh_11_23_io_out_control_0_propagate;
	wire [4:0] _mesh_11_23_io_out_control_0_shift;
	wire [2:0] _mesh_11_23_io_out_id_0;
	wire _mesh_11_23_io_out_last_0;
	wire _mesh_11_23_io_out_valid_0;
	wire [31:0] _mesh_11_22_io_out_a_0;
	wire [31:0] _mesh_11_22_io_out_c_0;
	wire [31:0] _mesh_11_22_io_out_b_0;
	wire _mesh_11_22_io_out_control_0_dataflow;
	wire _mesh_11_22_io_out_control_0_propagate;
	wire [4:0] _mesh_11_22_io_out_control_0_shift;
	wire [2:0] _mesh_11_22_io_out_id_0;
	wire _mesh_11_22_io_out_last_0;
	wire _mesh_11_22_io_out_valid_0;
	wire [31:0] _mesh_11_21_io_out_a_0;
	wire [31:0] _mesh_11_21_io_out_c_0;
	wire [31:0] _mesh_11_21_io_out_b_0;
	wire _mesh_11_21_io_out_control_0_dataflow;
	wire _mesh_11_21_io_out_control_0_propagate;
	wire [4:0] _mesh_11_21_io_out_control_0_shift;
	wire [2:0] _mesh_11_21_io_out_id_0;
	wire _mesh_11_21_io_out_last_0;
	wire _mesh_11_21_io_out_valid_0;
	wire [31:0] _mesh_11_20_io_out_a_0;
	wire [31:0] _mesh_11_20_io_out_c_0;
	wire [31:0] _mesh_11_20_io_out_b_0;
	wire _mesh_11_20_io_out_control_0_dataflow;
	wire _mesh_11_20_io_out_control_0_propagate;
	wire [4:0] _mesh_11_20_io_out_control_0_shift;
	wire [2:0] _mesh_11_20_io_out_id_0;
	wire _mesh_11_20_io_out_last_0;
	wire _mesh_11_20_io_out_valid_0;
	wire [31:0] _mesh_11_19_io_out_a_0;
	wire [31:0] _mesh_11_19_io_out_c_0;
	wire [31:0] _mesh_11_19_io_out_b_0;
	wire _mesh_11_19_io_out_control_0_dataflow;
	wire _mesh_11_19_io_out_control_0_propagate;
	wire [4:0] _mesh_11_19_io_out_control_0_shift;
	wire [2:0] _mesh_11_19_io_out_id_0;
	wire _mesh_11_19_io_out_last_0;
	wire _mesh_11_19_io_out_valid_0;
	wire [31:0] _mesh_11_18_io_out_a_0;
	wire [31:0] _mesh_11_18_io_out_c_0;
	wire [31:0] _mesh_11_18_io_out_b_0;
	wire _mesh_11_18_io_out_control_0_dataflow;
	wire _mesh_11_18_io_out_control_0_propagate;
	wire [4:0] _mesh_11_18_io_out_control_0_shift;
	wire [2:0] _mesh_11_18_io_out_id_0;
	wire _mesh_11_18_io_out_last_0;
	wire _mesh_11_18_io_out_valid_0;
	wire [31:0] _mesh_11_17_io_out_a_0;
	wire [31:0] _mesh_11_17_io_out_c_0;
	wire [31:0] _mesh_11_17_io_out_b_0;
	wire _mesh_11_17_io_out_control_0_dataflow;
	wire _mesh_11_17_io_out_control_0_propagate;
	wire [4:0] _mesh_11_17_io_out_control_0_shift;
	wire [2:0] _mesh_11_17_io_out_id_0;
	wire _mesh_11_17_io_out_last_0;
	wire _mesh_11_17_io_out_valid_0;
	wire [31:0] _mesh_11_16_io_out_a_0;
	wire [31:0] _mesh_11_16_io_out_c_0;
	wire [31:0] _mesh_11_16_io_out_b_0;
	wire _mesh_11_16_io_out_control_0_dataflow;
	wire _mesh_11_16_io_out_control_0_propagate;
	wire [4:0] _mesh_11_16_io_out_control_0_shift;
	wire [2:0] _mesh_11_16_io_out_id_0;
	wire _mesh_11_16_io_out_last_0;
	wire _mesh_11_16_io_out_valid_0;
	wire [31:0] _mesh_11_15_io_out_a_0;
	wire [31:0] _mesh_11_15_io_out_c_0;
	wire [31:0] _mesh_11_15_io_out_b_0;
	wire _mesh_11_15_io_out_control_0_dataflow;
	wire _mesh_11_15_io_out_control_0_propagate;
	wire [4:0] _mesh_11_15_io_out_control_0_shift;
	wire [2:0] _mesh_11_15_io_out_id_0;
	wire _mesh_11_15_io_out_last_0;
	wire _mesh_11_15_io_out_valid_0;
	wire [31:0] _mesh_11_14_io_out_a_0;
	wire [31:0] _mesh_11_14_io_out_c_0;
	wire [31:0] _mesh_11_14_io_out_b_0;
	wire _mesh_11_14_io_out_control_0_dataflow;
	wire _mesh_11_14_io_out_control_0_propagate;
	wire [4:0] _mesh_11_14_io_out_control_0_shift;
	wire [2:0] _mesh_11_14_io_out_id_0;
	wire _mesh_11_14_io_out_last_0;
	wire _mesh_11_14_io_out_valid_0;
	wire [31:0] _mesh_11_13_io_out_a_0;
	wire [31:0] _mesh_11_13_io_out_c_0;
	wire [31:0] _mesh_11_13_io_out_b_0;
	wire _mesh_11_13_io_out_control_0_dataflow;
	wire _mesh_11_13_io_out_control_0_propagate;
	wire [4:0] _mesh_11_13_io_out_control_0_shift;
	wire [2:0] _mesh_11_13_io_out_id_0;
	wire _mesh_11_13_io_out_last_0;
	wire _mesh_11_13_io_out_valid_0;
	wire [31:0] _mesh_11_12_io_out_a_0;
	wire [31:0] _mesh_11_12_io_out_c_0;
	wire [31:0] _mesh_11_12_io_out_b_0;
	wire _mesh_11_12_io_out_control_0_dataflow;
	wire _mesh_11_12_io_out_control_0_propagate;
	wire [4:0] _mesh_11_12_io_out_control_0_shift;
	wire [2:0] _mesh_11_12_io_out_id_0;
	wire _mesh_11_12_io_out_last_0;
	wire _mesh_11_12_io_out_valid_0;
	wire [31:0] _mesh_11_11_io_out_a_0;
	wire [31:0] _mesh_11_11_io_out_c_0;
	wire [31:0] _mesh_11_11_io_out_b_0;
	wire _mesh_11_11_io_out_control_0_dataflow;
	wire _mesh_11_11_io_out_control_0_propagate;
	wire [4:0] _mesh_11_11_io_out_control_0_shift;
	wire [2:0] _mesh_11_11_io_out_id_0;
	wire _mesh_11_11_io_out_last_0;
	wire _mesh_11_11_io_out_valid_0;
	wire [31:0] _mesh_11_10_io_out_a_0;
	wire [31:0] _mesh_11_10_io_out_c_0;
	wire [31:0] _mesh_11_10_io_out_b_0;
	wire _mesh_11_10_io_out_control_0_dataflow;
	wire _mesh_11_10_io_out_control_0_propagate;
	wire [4:0] _mesh_11_10_io_out_control_0_shift;
	wire [2:0] _mesh_11_10_io_out_id_0;
	wire _mesh_11_10_io_out_last_0;
	wire _mesh_11_10_io_out_valid_0;
	wire [31:0] _mesh_11_9_io_out_a_0;
	wire [31:0] _mesh_11_9_io_out_c_0;
	wire [31:0] _mesh_11_9_io_out_b_0;
	wire _mesh_11_9_io_out_control_0_dataflow;
	wire _mesh_11_9_io_out_control_0_propagate;
	wire [4:0] _mesh_11_9_io_out_control_0_shift;
	wire [2:0] _mesh_11_9_io_out_id_0;
	wire _mesh_11_9_io_out_last_0;
	wire _mesh_11_9_io_out_valid_0;
	wire [31:0] _mesh_11_8_io_out_a_0;
	wire [31:0] _mesh_11_8_io_out_c_0;
	wire [31:0] _mesh_11_8_io_out_b_0;
	wire _mesh_11_8_io_out_control_0_dataflow;
	wire _mesh_11_8_io_out_control_0_propagate;
	wire [4:0] _mesh_11_8_io_out_control_0_shift;
	wire [2:0] _mesh_11_8_io_out_id_0;
	wire _mesh_11_8_io_out_last_0;
	wire _mesh_11_8_io_out_valid_0;
	wire [31:0] _mesh_11_7_io_out_a_0;
	wire [31:0] _mesh_11_7_io_out_c_0;
	wire [31:0] _mesh_11_7_io_out_b_0;
	wire _mesh_11_7_io_out_control_0_dataflow;
	wire _mesh_11_7_io_out_control_0_propagate;
	wire [4:0] _mesh_11_7_io_out_control_0_shift;
	wire [2:0] _mesh_11_7_io_out_id_0;
	wire _mesh_11_7_io_out_last_0;
	wire _mesh_11_7_io_out_valid_0;
	wire [31:0] _mesh_11_6_io_out_a_0;
	wire [31:0] _mesh_11_6_io_out_c_0;
	wire [31:0] _mesh_11_6_io_out_b_0;
	wire _mesh_11_6_io_out_control_0_dataflow;
	wire _mesh_11_6_io_out_control_0_propagate;
	wire [4:0] _mesh_11_6_io_out_control_0_shift;
	wire [2:0] _mesh_11_6_io_out_id_0;
	wire _mesh_11_6_io_out_last_0;
	wire _mesh_11_6_io_out_valid_0;
	wire [31:0] _mesh_11_5_io_out_a_0;
	wire [31:0] _mesh_11_5_io_out_c_0;
	wire [31:0] _mesh_11_5_io_out_b_0;
	wire _mesh_11_5_io_out_control_0_dataflow;
	wire _mesh_11_5_io_out_control_0_propagate;
	wire [4:0] _mesh_11_5_io_out_control_0_shift;
	wire [2:0] _mesh_11_5_io_out_id_0;
	wire _mesh_11_5_io_out_last_0;
	wire _mesh_11_5_io_out_valid_0;
	wire [31:0] _mesh_11_4_io_out_a_0;
	wire [31:0] _mesh_11_4_io_out_c_0;
	wire [31:0] _mesh_11_4_io_out_b_0;
	wire _mesh_11_4_io_out_control_0_dataflow;
	wire _mesh_11_4_io_out_control_0_propagate;
	wire [4:0] _mesh_11_4_io_out_control_0_shift;
	wire [2:0] _mesh_11_4_io_out_id_0;
	wire _mesh_11_4_io_out_last_0;
	wire _mesh_11_4_io_out_valid_0;
	wire [31:0] _mesh_11_3_io_out_a_0;
	wire [31:0] _mesh_11_3_io_out_c_0;
	wire [31:0] _mesh_11_3_io_out_b_0;
	wire _mesh_11_3_io_out_control_0_dataflow;
	wire _mesh_11_3_io_out_control_0_propagate;
	wire [4:0] _mesh_11_3_io_out_control_0_shift;
	wire [2:0] _mesh_11_3_io_out_id_0;
	wire _mesh_11_3_io_out_last_0;
	wire _mesh_11_3_io_out_valid_0;
	wire [31:0] _mesh_11_2_io_out_a_0;
	wire [31:0] _mesh_11_2_io_out_c_0;
	wire [31:0] _mesh_11_2_io_out_b_0;
	wire _mesh_11_2_io_out_control_0_dataflow;
	wire _mesh_11_2_io_out_control_0_propagate;
	wire [4:0] _mesh_11_2_io_out_control_0_shift;
	wire [2:0] _mesh_11_2_io_out_id_0;
	wire _mesh_11_2_io_out_last_0;
	wire _mesh_11_2_io_out_valid_0;
	wire [31:0] _mesh_11_1_io_out_a_0;
	wire [31:0] _mesh_11_1_io_out_c_0;
	wire [31:0] _mesh_11_1_io_out_b_0;
	wire _mesh_11_1_io_out_control_0_dataflow;
	wire _mesh_11_1_io_out_control_0_propagate;
	wire [4:0] _mesh_11_1_io_out_control_0_shift;
	wire [2:0] _mesh_11_1_io_out_id_0;
	wire _mesh_11_1_io_out_last_0;
	wire _mesh_11_1_io_out_valid_0;
	wire [31:0] _mesh_11_0_io_out_a_0;
	wire [31:0] _mesh_11_0_io_out_c_0;
	wire [31:0] _mesh_11_0_io_out_b_0;
	wire _mesh_11_0_io_out_control_0_dataflow;
	wire _mesh_11_0_io_out_control_0_propagate;
	wire [4:0] _mesh_11_0_io_out_control_0_shift;
	wire [2:0] _mesh_11_0_io_out_id_0;
	wire _mesh_11_0_io_out_last_0;
	wire _mesh_11_0_io_out_valid_0;
	wire [31:0] _mesh_10_31_io_out_a_0;
	wire [31:0] _mesh_10_31_io_out_c_0;
	wire [31:0] _mesh_10_31_io_out_b_0;
	wire _mesh_10_31_io_out_control_0_dataflow;
	wire _mesh_10_31_io_out_control_0_propagate;
	wire [4:0] _mesh_10_31_io_out_control_0_shift;
	wire [2:0] _mesh_10_31_io_out_id_0;
	wire _mesh_10_31_io_out_last_0;
	wire _mesh_10_31_io_out_valid_0;
	wire [31:0] _mesh_10_30_io_out_a_0;
	wire [31:0] _mesh_10_30_io_out_c_0;
	wire [31:0] _mesh_10_30_io_out_b_0;
	wire _mesh_10_30_io_out_control_0_dataflow;
	wire _mesh_10_30_io_out_control_0_propagate;
	wire [4:0] _mesh_10_30_io_out_control_0_shift;
	wire [2:0] _mesh_10_30_io_out_id_0;
	wire _mesh_10_30_io_out_last_0;
	wire _mesh_10_30_io_out_valid_0;
	wire [31:0] _mesh_10_29_io_out_a_0;
	wire [31:0] _mesh_10_29_io_out_c_0;
	wire [31:0] _mesh_10_29_io_out_b_0;
	wire _mesh_10_29_io_out_control_0_dataflow;
	wire _mesh_10_29_io_out_control_0_propagate;
	wire [4:0] _mesh_10_29_io_out_control_0_shift;
	wire [2:0] _mesh_10_29_io_out_id_0;
	wire _mesh_10_29_io_out_last_0;
	wire _mesh_10_29_io_out_valid_0;
	wire [31:0] _mesh_10_28_io_out_a_0;
	wire [31:0] _mesh_10_28_io_out_c_0;
	wire [31:0] _mesh_10_28_io_out_b_0;
	wire _mesh_10_28_io_out_control_0_dataflow;
	wire _mesh_10_28_io_out_control_0_propagate;
	wire [4:0] _mesh_10_28_io_out_control_0_shift;
	wire [2:0] _mesh_10_28_io_out_id_0;
	wire _mesh_10_28_io_out_last_0;
	wire _mesh_10_28_io_out_valid_0;
	wire [31:0] _mesh_10_27_io_out_a_0;
	wire [31:0] _mesh_10_27_io_out_c_0;
	wire [31:0] _mesh_10_27_io_out_b_0;
	wire _mesh_10_27_io_out_control_0_dataflow;
	wire _mesh_10_27_io_out_control_0_propagate;
	wire [4:0] _mesh_10_27_io_out_control_0_shift;
	wire [2:0] _mesh_10_27_io_out_id_0;
	wire _mesh_10_27_io_out_last_0;
	wire _mesh_10_27_io_out_valid_0;
	wire [31:0] _mesh_10_26_io_out_a_0;
	wire [31:0] _mesh_10_26_io_out_c_0;
	wire [31:0] _mesh_10_26_io_out_b_0;
	wire _mesh_10_26_io_out_control_0_dataflow;
	wire _mesh_10_26_io_out_control_0_propagate;
	wire [4:0] _mesh_10_26_io_out_control_0_shift;
	wire [2:0] _mesh_10_26_io_out_id_0;
	wire _mesh_10_26_io_out_last_0;
	wire _mesh_10_26_io_out_valid_0;
	wire [31:0] _mesh_10_25_io_out_a_0;
	wire [31:0] _mesh_10_25_io_out_c_0;
	wire [31:0] _mesh_10_25_io_out_b_0;
	wire _mesh_10_25_io_out_control_0_dataflow;
	wire _mesh_10_25_io_out_control_0_propagate;
	wire [4:0] _mesh_10_25_io_out_control_0_shift;
	wire [2:0] _mesh_10_25_io_out_id_0;
	wire _mesh_10_25_io_out_last_0;
	wire _mesh_10_25_io_out_valid_0;
	wire [31:0] _mesh_10_24_io_out_a_0;
	wire [31:0] _mesh_10_24_io_out_c_0;
	wire [31:0] _mesh_10_24_io_out_b_0;
	wire _mesh_10_24_io_out_control_0_dataflow;
	wire _mesh_10_24_io_out_control_0_propagate;
	wire [4:0] _mesh_10_24_io_out_control_0_shift;
	wire [2:0] _mesh_10_24_io_out_id_0;
	wire _mesh_10_24_io_out_last_0;
	wire _mesh_10_24_io_out_valid_0;
	wire [31:0] _mesh_10_23_io_out_a_0;
	wire [31:0] _mesh_10_23_io_out_c_0;
	wire [31:0] _mesh_10_23_io_out_b_0;
	wire _mesh_10_23_io_out_control_0_dataflow;
	wire _mesh_10_23_io_out_control_0_propagate;
	wire [4:0] _mesh_10_23_io_out_control_0_shift;
	wire [2:0] _mesh_10_23_io_out_id_0;
	wire _mesh_10_23_io_out_last_0;
	wire _mesh_10_23_io_out_valid_0;
	wire [31:0] _mesh_10_22_io_out_a_0;
	wire [31:0] _mesh_10_22_io_out_c_0;
	wire [31:0] _mesh_10_22_io_out_b_0;
	wire _mesh_10_22_io_out_control_0_dataflow;
	wire _mesh_10_22_io_out_control_0_propagate;
	wire [4:0] _mesh_10_22_io_out_control_0_shift;
	wire [2:0] _mesh_10_22_io_out_id_0;
	wire _mesh_10_22_io_out_last_0;
	wire _mesh_10_22_io_out_valid_0;
	wire [31:0] _mesh_10_21_io_out_a_0;
	wire [31:0] _mesh_10_21_io_out_c_0;
	wire [31:0] _mesh_10_21_io_out_b_0;
	wire _mesh_10_21_io_out_control_0_dataflow;
	wire _mesh_10_21_io_out_control_0_propagate;
	wire [4:0] _mesh_10_21_io_out_control_0_shift;
	wire [2:0] _mesh_10_21_io_out_id_0;
	wire _mesh_10_21_io_out_last_0;
	wire _mesh_10_21_io_out_valid_0;
	wire [31:0] _mesh_10_20_io_out_a_0;
	wire [31:0] _mesh_10_20_io_out_c_0;
	wire [31:0] _mesh_10_20_io_out_b_0;
	wire _mesh_10_20_io_out_control_0_dataflow;
	wire _mesh_10_20_io_out_control_0_propagate;
	wire [4:0] _mesh_10_20_io_out_control_0_shift;
	wire [2:0] _mesh_10_20_io_out_id_0;
	wire _mesh_10_20_io_out_last_0;
	wire _mesh_10_20_io_out_valid_0;
	wire [31:0] _mesh_10_19_io_out_a_0;
	wire [31:0] _mesh_10_19_io_out_c_0;
	wire [31:0] _mesh_10_19_io_out_b_0;
	wire _mesh_10_19_io_out_control_0_dataflow;
	wire _mesh_10_19_io_out_control_0_propagate;
	wire [4:0] _mesh_10_19_io_out_control_0_shift;
	wire [2:0] _mesh_10_19_io_out_id_0;
	wire _mesh_10_19_io_out_last_0;
	wire _mesh_10_19_io_out_valid_0;
	wire [31:0] _mesh_10_18_io_out_a_0;
	wire [31:0] _mesh_10_18_io_out_c_0;
	wire [31:0] _mesh_10_18_io_out_b_0;
	wire _mesh_10_18_io_out_control_0_dataflow;
	wire _mesh_10_18_io_out_control_0_propagate;
	wire [4:0] _mesh_10_18_io_out_control_0_shift;
	wire [2:0] _mesh_10_18_io_out_id_0;
	wire _mesh_10_18_io_out_last_0;
	wire _mesh_10_18_io_out_valid_0;
	wire [31:0] _mesh_10_17_io_out_a_0;
	wire [31:0] _mesh_10_17_io_out_c_0;
	wire [31:0] _mesh_10_17_io_out_b_0;
	wire _mesh_10_17_io_out_control_0_dataflow;
	wire _mesh_10_17_io_out_control_0_propagate;
	wire [4:0] _mesh_10_17_io_out_control_0_shift;
	wire [2:0] _mesh_10_17_io_out_id_0;
	wire _mesh_10_17_io_out_last_0;
	wire _mesh_10_17_io_out_valid_0;
	wire [31:0] _mesh_10_16_io_out_a_0;
	wire [31:0] _mesh_10_16_io_out_c_0;
	wire [31:0] _mesh_10_16_io_out_b_0;
	wire _mesh_10_16_io_out_control_0_dataflow;
	wire _mesh_10_16_io_out_control_0_propagate;
	wire [4:0] _mesh_10_16_io_out_control_0_shift;
	wire [2:0] _mesh_10_16_io_out_id_0;
	wire _mesh_10_16_io_out_last_0;
	wire _mesh_10_16_io_out_valid_0;
	wire [31:0] _mesh_10_15_io_out_a_0;
	wire [31:0] _mesh_10_15_io_out_c_0;
	wire [31:0] _mesh_10_15_io_out_b_0;
	wire _mesh_10_15_io_out_control_0_dataflow;
	wire _mesh_10_15_io_out_control_0_propagate;
	wire [4:0] _mesh_10_15_io_out_control_0_shift;
	wire [2:0] _mesh_10_15_io_out_id_0;
	wire _mesh_10_15_io_out_last_0;
	wire _mesh_10_15_io_out_valid_0;
	wire [31:0] _mesh_10_14_io_out_a_0;
	wire [31:0] _mesh_10_14_io_out_c_0;
	wire [31:0] _mesh_10_14_io_out_b_0;
	wire _mesh_10_14_io_out_control_0_dataflow;
	wire _mesh_10_14_io_out_control_0_propagate;
	wire [4:0] _mesh_10_14_io_out_control_0_shift;
	wire [2:0] _mesh_10_14_io_out_id_0;
	wire _mesh_10_14_io_out_last_0;
	wire _mesh_10_14_io_out_valid_0;
	wire [31:0] _mesh_10_13_io_out_a_0;
	wire [31:0] _mesh_10_13_io_out_c_0;
	wire [31:0] _mesh_10_13_io_out_b_0;
	wire _mesh_10_13_io_out_control_0_dataflow;
	wire _mesh_10_13_io_out_control_0_propagate;
	wire [4:0] _mesh_10_13_io_out_control_0_shift;
	wire [2:0] _mesh_10_13_io_out_id_0;
	wire _mesh_10_13_io_out_last_0;
	wire _mesh_10_13_io_out_valid_0;
	wire [31:0] _mesh_10_12_io_out_a_0;
	wire [31:0] _mesh_10_12_io_out_c_0;
	wire [31:0] _mesh_10_12_io_out_b_0;
	wire _mesh_10_12_io_out_control_0_dataflow;
	wire _mesh_10_12_io_out_control_0_propagate;
	wire [4:0] _mesh_10_12_io_out_control_0_shift;
	wire [2:0] _mesh_10_12_io_out_id_0;
	wire _mesh_10_12_io_out_last_0;
	wire _mesh_10_12_io_out_valid_0;
	wire [31:0] _mesh_10_11_io_out_a_0;
	wire [31:0] _mesh_10_11_io_out_c_0;
	wire [31:0] _mesh_10_11_io_out_b_0;
	wire _mesh_10_11_io_out_control_0_dataflow;
	wire _mesh_10_11_io_out_control_0_propagate;
	wire [4:0] _mesh_10_11_io_out_control_0_shift;
	wire [2:0] _mesh_10_11_io_out_id_0;
	wire _mesh_10_11_io_out_last_0;
	wire _mesh_10_11_io_out_valid_0;
	wire [31:0] _mesh_10_10_io_out_a_0;
	wire [31:0] _mesh_10_10_io_out_c_0;
	wire [31:0] _mesh_10_10_io_out_b_0;
	wire _mesh_10_10_io_out_control_0_dataflow;
	wire _mesh_10_10_io_out_control_0_propagate;
	wire [4:0] _mesh_10_10_io_out_control_0_shift;
	wire [2:0] _mesh_10_10_io_out_id_0;
	wire _mesh_10_10_io_out_last_0;
	wire _mesh_10_10_io_out_valid_0;
	wire [31:0] _mesh_10_9_io_out_a_0;
	wire [31:0] _mesh_10_9_io_out_c_0;
	wire [31:0] _mesh_10_9_io_out_b_0;
	wire _mesh_10_9_io_out_control_0_dataflow;
	wire _mesh_10_9_io_out_control_0_propagate;
	wire [4:0] _mesh_10_9_io_out_control_0_shift;
	wire [2:0] _mesh_10_9_io_out_id_0;
	wire _mesh_10_9_io_out_last_0;
	wire _mesh_10_9_io_out_valid_0;
	wire [31:0] _mesh_10_8_io_out_a_0;
	wire [31:0] _mesh_10_8_io_out_c_0;
	wire [31:0] _mesh_10_8_io_out_b_0;
	wire _mesh_10_8_io_out_control_0_dataflow;
	wire _mesh_10_8_io_out_control_0_propagate;
	wire [4:0] _mesh_10_8_io_out_control_0_shift;
	wire [2:0] _mesh_10_8_io_out_id_0;
	wire _mesh_10_8_io_out_last_0;
	wire _mesh_10_8_io_out_valid_0;
	wire [31:0] _mesh_10_7_io_out_a_0;
	wire [31:0] _mesh_10_7_io_out_c_0;
	wire [31:0] _mesh_10_7_io_out_b_0;
	wire _mesh_10_7_io_out_control_0_dataflow;
	wire _mesh_10_7_io_out_control_0_propagate;
	wire [4:0] _mesh_10_7_io_out_control_0_shift;
	wire [2:0] _mesh_10_7_io_out_id_0;
	wire _mesh_10_7_io_out_last_0;
	wire _mesh_10_7_io_out_valid_0;
	wire [31:0] _mesh_10_6_io_out_a_0;
	wire [31:0] _mesh_10_6_io_out_c_0;
	wire [31:0] _mesh_10_6_io_out_b_0;
	wire _mesh_10_6_io_out_control_0_dataflow;
	wire _mesh_10_6_io_out_control_0_propagate;
	wire [4:0] _mesh_10_6_io_out_control_0_shift;
	wire [2:0] _mesh_10_6_io_out_id_0;
	wire _mesh_10_6_io_out_last_0;
	wire _mesh_10_6_io_out_valid_0;
	wire [31:0] _mesh_10_5_io_out_a_0;
	wire [31:0] _mesh_10_5_io_out_c_0;
	wire [31:0] _mesh_10_5_io_out_b_0;
	wire _mesh_10_5_io_out_control_0_dataflow;
	wire _mesh_10_5_io_out_control_0_propagate;
	wire [4:0] _mesh_10_5_io_out_control_0_shift;
	wire [2:0] _mesh_10_5_io_out_id_0;
	wire _mesh_10_5_io_out_last_0;
	wire _mesh_10_5_io_out_valid_0;
	wire [31:0] _mesh_10_4_io_out_a_0;
	wire [31:0] _mesh_10_4_io_out_c_0;
	wire [31:0] _mesh_10_4_io_out_b_0;
	wire _mesh_10_4_io_out_control_0_dataflow;
	wire _mesh_10_4_io_out_control_0_propagate;
	wire [4:0] _mesh_10_4_io_out_control_0_shift;
	wire [2:0] _mesh_10_4_io_out_id_0;
	wire _mesh_10_4_io_out_last_0;
	wire _mesh_10_4_io_out_valid_0;
	wire [31:0] _mesh_10_3_io_out_a_0;
	wire [31:0] _mesh_10_3_io_out_c_0;
	wire [31:0] _mesh_10_3_io_out_b_0;
	wire _mesh_10_3_io_out_control_0_dataflow;
	wire _mesh_10_3_io_out_control_0_propagate;
	wire [4:0] _mesh_10_3_io_out_control_0_shift;
	wire [2:0] _mesh_10_3_io_out_id_0;
	wire _mesh_10_3_io_out_last_0;
	wire _mesh_10_3_io_out_valid_0;
	wire [31:0] _mesh_10_2_io_out_a_0;
	wire [31:0] _mesh_10_2_io_out_c_0;
	wire [31:0] _mesh_10_2_io_out_b_0;
	wire _mesh_10_2_io_out_control_0_dataflow;
	wire _mesh_10_2_io_out_control_0_propagate;
	wire [4:0] _mesh_10_2_io_out_control_0_shift;
	wire [2:0] _mesh_10_2_io_out_id_0;
	wire _mesh_10_2_io_out_last_0;
	wire _mesh_10_2_io_out_valid_0;
	wire [31:0] _mesh_10_1_io_out_a_0;
	wire [31:0] _mesh_10_1_io_out_c_0;
	wire [31:0] _mesh_10_1_io_out_b_0;
	wire _mesh_10_1_io_out_control_0_dataflow;
	wire _mesh_10_1_io_out_control_0_propagate;
	wire [4:0] _mesh_10_1_io_out_control_0_shift;
	wire [2:0] _mesh_10_1_io_out_id_0;
	wire _mesh_10_1_io_out_last_0;
	wire _mesh_10_1_io_out_valid_0;
	wire [31:0] _mesh_10_0_io_out_a_0;
	wire [31:0] _mesh_10_0_io_out_c_0;
	wire [31:0] _mesh_10_0_io_out_b_0;
	wire _mesh_10_0_io_out_control_0_dataflow;
	wire _mesh_10_0_io_out_control_0_propagate;
	wire [4:0] _mesh_10_0_io_out_control_0_shift;
	wire [2:0] _mesh_10_0_io_out_id_0;
	wire _mesh_10_0_io_out_last_0;
	wire _mesh_10_0_io_out_valid_0;
	wire [31:0] _mesh_9_31_io_out_a_0;
	wire [31:0] _mesh_9_31_io_out_c_0;
	wire [31:0] _mesh_9_31_io_out_b_0;
	wire _mesh_9_31_io_out_control_0_dataflow;
	wire _mesh_9_31_io_out_control_0_propagate;
	wire [4:0] _mesh_9_31_io_out_control_0_shift;
	wire [2:0] _mesh_9_31_io_out_id_0;
	wire _mesh_9_31_io_out_last_0;
	wire _mesh_9_31_io_out_valid_0;
	wire [31:0] _mesh_9_30_io_out_a_0;
	wire [31:0] _mesh_9_30_io_out_c_0;
	wire [31:0] _mesh_9_30_io_out_b_0;
	wire _mesh_9_30_io_out_control_0_dataflow;
	wire _mesh_9_30_io_out_control_0_propagate;
	wire [4:0] _mesh_9_30_io_out_control_0_shift;
	wire [2:0] _mesh_9_30_io_out_id_0;
	wire _mesh_9_30_io_out_last_0;
	wire _mesh_9_30_io_out_valid_0;
	wire [31:0] _mesh_9_29_io_out_a_0;
	wire [31:0] _mesh_9_29_io_out_c_0;
	wire [31:0] _mesh_9_29_io_out_b_0;
	wire _mesh_9_29_io_out_control_0_dataflow;
	wire _mesh_9_29_io_out_control_0_propagate;
	wire [4:0] _mesh_9_29_io_out_control_0_shift;
	wire [2:0] _mesh_9_29_io_out_id_0;
	wire _mesh_9_29_io_out_last_0;
	wire _mesh_9_29_io_out_valid_0;
	wire [31:0] _mesh_9_28_io_out_a_0;
	wire [31:0] _mesh_9_28_io_out_c_0;
	wire [31:0] _mesh_9_28_io_out_b_0;
	wire _mesh_9_28_io_out_control_0_dataflow;
	wire _mesh_9_28_io_out_control_0_propagate;
	wire [4:0] _mesh_9_28_io_out_control_0_shift;
	wire [2:0] _mesh_9_28_io_out_id_0;
	wire _mesh_9_28_io_out_last_0;
	wire _mesh_9_28_io_out_valid_0;
	wire [31:0] _mesh_9_27_io_out_a_0;
	wire [31:0] _mesh_9_27_io_out_c_0;
	wire [31:0] _mesh_9_27_io_out_b_0;
	wire _mesh_9_27_io_out_control_0_dataflow;
	wire _mesh_9_27_io_out_control_0_propagate;
	wire [4:0] _mesh_9_27_io_out_control_0_shift;
	wire [2:0] _mesh_9_27_io_out_id_0;
	wire _mesh_9_27_io_out_last_0;
	wire _mesh_9_27_io_out_valid_0;
	wire [31:0] _mesh_9_26_io_out_a_0;
	wire [31:0] _mesh_9_26_io_out_c_0;
	wire [31:0] _mesh_9_26_io_out_b_0;
	wire _mesh_9_26_io_out_control_0_dataflow;
	wire _mesh_9_26_io_out_control_0_propagate;
	wire [4:0] _mesh_9_26_io_out_control_0_shift;
	wire [2:0] _mesh_9_26_io_out_id_0;
	wire _mesh_9_26_io_out_last_0;
	wire _mesh_9_26_io_out_valid_0;
	wire [31:0] _mesh_9_25_io_out_a_0;
	wire [31:0] _mesh_9_25_io_out_c_0;
	wire [31:0] _mesh_9_25_io_out_b_0;
	wire _mesh_9_25_io_out_control_0_dataflow;
	wire _mesh_9_25_io_out_control_0_propagate;
	wire [4:0] _mesh_9_25_io_out_control_0_shift;
	wire [2:0] _mesh_9_25_io_out_id_0;
	wire _mesh_9_25_io_out_last_0;
	wire _mesh_9_25_io_out_valid_0;
	wire [31:0] _mesh_9_24_io_out_a_0;
	wire [31:0] _mesh_9_24_io_out_c_0;
	wire [31:0] _mesh_9_24_io_out_b_0;
	wire _mesh_9_24_io_out_control_0_dataflow;
	wire _mesh_9_24_io_out_control_0_propagate;
	wire [4:0] _mesh_9_24_io_out_control_0_shift;
	wire [2:0] _mesh_9_24_io_out_id_0;
	wire _mesh_9_24_io_out_last_0;
	wire _mesh_9_24_io_out_valid_0;
	wire [31:0] _mesh_9_23_io_out_a_0;
	wire [31:0] _mesh_9_23_io_out_c_0;
	wire [31:0] _mesh_9_23_io_out_b_0;
	wire _mesh_9_23_io_out_control_0_dataflow;
	wire _mesh_9_23_io_out_control_0_propagate;
	wire [4:0] _mesh_9_23_io_out_control_0_shift;
	wire [2:0] _mesh_9_23_io_out_id_0;
	wire _mesh_9_23_io_out_last_0;
	wire _mesh_9_23_io_out_valid_0;
	wire [31:0] _mesh_9_22_io_out_a_0;
	wire [31:0] _mesh_9_22_io_out_c_0;
	wire [31:0] _mesh_9_22_io_out_b_0;
	wire _mesh_9_22_io_out_control_0_dataflow;
	wire _mesh_9_22_io_out_control_0_propagate;
	wire [4:0] _mesh_9_22_io_out_control_0_shift;
	wire [2:0] _mesh_9_22_io_out_id_0;
	wire _mesh_9_22_io_out_last_0;
	wire _mesh_9_22_io_out_valid_0;
	wire [31:0] _mesh_9_21_io_out_a_0;
	wire [31:0] _mesh_9_21_io_out_c_0;
	wire [31:0] _mesh_9_21_io_out_b_0;
	wire _mesh_9_21_io_out_control_0_dataflow;
	wire _mesh_9_21_io_out_control_0_propagate;
	wire [4:0] _mesh_9_21_io_out_control_0_shift;
	wire [2:0] _mesh_9_21_io_out_id_0;
	wire _mesh_9_21_io_out_last_0;
	wire _mesh_9_21_io_out_valid_0;
	wire [31:0] _mesh_9_20_io_out_a_0;
	wire [31:0] _mesh_9_20_io_out_c_0;
	wire [31:0] _mesh_9_20_io_out_b_0;
	wire _mesh_9_20_io_out_control_0_dataflow;
	wire _mesh_9_20_io_out_control_0_propagate;
	wire [4:0] _mesh_9_20_io_out_control_0_shift;
	wire [2:0] _mesh_9_20_io_out_id_0;
	wire _mesh_9_20_io_out_last_0;
	wire _mesh_9_20_io_out_valid_0;
	wire [31:0] _mesh_9_19_io_out_a_0;
	wire [31:0] _mesh_9_19_io_out_c_0;
	wire [31:0] _mesh_9_19_io_out_b_0;
	wire _mesh_9_19_io_out_control_0_dataflow;
	wire _mesh_9_19_io_out_control_0_propagate;
	wire [4:0] _mesh_9_19_io_out_control_0_shift;
	wire [2:0] _mesh_9_19_io_out_id_0;
	wire _mesh_9_19_io_out_last_0;
	wire _mesh_9_19_io_out_valid_0;
	wire [31:0] _mesh_9_18_io_out_a_0;
	wire [31:0] _mesh_9_18_io_out_c_0;
	wire [31:0] _mesh_9_18_io_out_b_0;
	wire _mesh_9_18_io_out_control_0_dataflow;
	wire _mesh_9_18_io_out_control_0_propagate;
	wire [4:0] _mesh_9_18_io_out_control_0_shift;
	wire [2:0] _mesh_9_18_io_out_id_0;
	wire _mesh_9_18_io_out_last_0;
	wire _mesh_9_18_io_out_valid_0;
	wire [31:0] _mesh_9_17_io_out_a_0;
	wire [31:0] _mesh_9_17_io_out_c_0;
	wire [31:0] _mesh_9_17_io_out_b_0;
	wire _mesh_9_17_io_out_control_0_dataflow;
	wire _mesh_9_17_io_out_control_0_propagate;
	wire [4:0] _mesh_9_17_io_out_control_0_shift;
	wire [2:0] _mesh_9_17_io_out_id_0;
	wire _mesh_9_17_io_out_last_0;
	wire _mesh_9_17_io_out_valid_0;
	wire [31:0] _mesh_9_16_io_out_a_0;
	wire [31:0] _mesh_9_16_io_out_c_0;
	wire [31:0] _mesh_9_16_io_out_b_0;
	wire _mesh_9_16_io_out_control_0_dataflow;
	wire _mesh_9_16_io_out_control_0_propagate;
	wire [4:0] _mesh_9_16_io_out_control_0_shift;
	wire [2:0] _mesh_9_16_io_out_id_0;
	wire _mesh_9_16_io_out_last_0;
	wire _mesh_9_16_io_out_valid_0;
	wire [31:0] _mesh_9_15_io_out_a_0;
	wire [31:0] _mesh_9_15_io_out_c_0;
	wire [31:0] _mesh_9_15_io_out_b_0;
	wire _mesh_9_15_io_out_control_0_dataflow;
	wire _mesh_9_15_io_out_control_0_propagate;
	wire [4:0] _mesh_9_15_io_out_control_0_shift;
	wire [2:0] _mesh_9_15_io_out_id_0;
	wire _mesh_9_15_io_out_last_0;
	wire _mesh_9_15_io_out_valid_0;
	wire [31:0] _mesh_9_14_io_out_a_0;
	wire [31:0] _mesh_9_14_io_out_c_0;
	wire [31:0] _mesh_9_14_io_out_b_0;
	wire _mesh_9_14_io_out_control_0_dataflow;
	wire _mesh_9_14_io_out_control_0_propagate;
	wire [4:0] _mesh_9_14_io_out_control_0_shift;
	wire [2:0] _mesh_9_14_io_out_id_0;
	wire _mesh_9_14_io_out_last_0;
	wire _mesh_9_14_io_out_valid_0;
	wire [31:0] _mesh_9_13_io_out_a_0;
	wire [31:0] _mesh_9_13_io_out_c_0;
	wire [31:0] _mesh_9_13_io_out_b_0;
	wire _mesh_9_13_io_out_control_0_dataflow;
	wire _mesh_9_13_io_out_control_0_propagate;
	wire [4:0] _mesh_9_13_io_out_control_0_shift;
	wire [2:0] _mesh_9_13_io_out_id_0;
	wire _mesh_9_13_io_out_last_0;
	wire _mesh_9_13_io_out_valid_0;
	wire [31:0] _mesh_9_12_io_out_a_0;
	wire [31:0] _mesh_9_12_io_out_c_0;
	wire [31:0] _mesh_9_12_io_out_b_0;
	wire _mesh_9_12_io_out_control_0_dataflow;
	wire _mesh_9_12_io_out_control_0_propagate;
	wire [4:0] _mesh_9_12_io_out_control_0_shift;
	wire [2:0] _mesh_9_12_io_out_id_0;
	wire _mesh_9_12_io_out_last_0;
	wire _mesh_9_12_io_out_valid_0;
	wire [31:0] _mesh_9_11_io_out_a_0;
	wire [31:0] _mesh_9_11_io_out_c_0;
	wire [31:0] _mesh_9_11_io_out_b_0;
	wire _mesh_9_11_io_out_control_0_dataflow;
	wire _mesh_9_11_io_out_control_0_propagate;
	wire [4:0] _mesh_9_11_io_out_control_0_shift;
	wire [2:0] _mesh_9_11_io_out_id_0;
	wire _mesh_9_11_io_out_last_0;
	wire _mesh_9_11_io_out_valid_0;
	wire [31:0] _mesh_9_10_io_out_a_0;
	wire [31:0] _mesh_9_10_io_out_c_0;
	wire [31:0] _mesh_9_10_io_out_b_0;
	wire _mesh_9_10_io_out_control_0_dataflow;
	wire _mesh_9_10_io_out_control_0_propagate;
	wire [4:0] _mesh_9_10_io_out_control_0_shift;
	wire [2:0] _mesh_9_10_io_out_id_0;
	wire _mesh_9_10_io_out_last_0;
	wire _mesh_9_10_io_out_valid_0;
	wire [31:0] _mesh_9_9_io_out_a_0;
	wire [31:0] _mesh_9_9_io_out_c_0;
	wire [31:0] _mesh_9_9_io_out_b_0;
	wire _mesh_9_9_io_out_control_0_dataflow;
	wire _mesh_9_9_io_out_control_0_propagate;
	wire [4:0] _mesh_9_9_io_out_control_0_shift;
	wire [2:0] _mesh_9_9_io_out_id_0;
	wire _mesh_9_9_io_out_last_0;
	wire _mesh_9_9_io_out_valid_0;
	wire [31:0] _mesh_9_8_io_out_a_0;
	wire [31:0] _mesh_9_8_io_out_c_0;
	wire [31:0] _mesh_9_8_io_out_b_0;
	wire _mesh_9_8_io_out_control_0_dataflow;
	wire _mesh_9_8_io_out_control_0_propagate;
	wire [4:0] _mesh_9_8_io_out_control_0_shift;
	wire [2:0] _mesh_9_8_io_out_id_0;
	wire _mesh_9_8_io_out_last_0;
	wire _mesh_9_8_io_out_valid_0;
	wire [31:0] _mesh_9_7_io_out_a_0;
	wire [31:0] _mesh_9_7_io_out_c_0;
	wire [31:0] _mesh_9_7_io_out_b_0;
	wire _mesh_9_7_io_out_control_0_dataflow;
	wire _mesh_9_7_io_out_control_0_propagate;
	wire [4:0] _mesh_9_7_io_out_control_0_shift;
	wire [2:0] _mesh_9_7_io_out_id_0;
	wire _mesh_9_7_io_out_last_0;
	wire _mesh_9_7_io_out_valid_0;
	wire [31:0] _mesh_9_6_io_out_a_0;
	wire [31:0] _mesh_9_6_io_out_c_0;
	wire [31:0] _mesh_9_6_io_out_b_0;
	wire _mesh_9_6_io_out_control_0_dataflow;
	wire _mesh_9_6_io_out_control_0_propagate;
	wire [4:0] _mesh_9_6_io_out_control_0_shift;
	wire [2:0] _mesh_9_6_io_out_id_0;
	wire _mesh_9_6_io_out_last_0;
	wire _mesh_9_6_io_out_valid_0;
	wire [31:0] _mesh_9_5_io_out_a_0;
	wire [31:0] _mesh_9_5_io_out_c_0;
	wire [31:0] _mesh_9_5_io_out_b_0;
	wire _mesh_9_5_io_out_control_0_dataflow;
	wire _mesh_9_5_io_out_control_0_propagate;
	wire [4:0] _mesh_9_5_io_out_control_0_shift;
	wire [2:0] _mesh_9_5_io_out_id_0;
	wire _mesh_9_5_io_out_last_0;
	wire _mesh_9_5_io_out_valid_0;
	wire [31:0] _mesh_9_4_io_out_a_0;
	wire [31:0] _mesh_9_4_io_out_c_0;
	wire [31:0] _mesh_9_4_io_out_b_0;
	wire _mesh_9_4_io_out_control_0_dataflow;
	wire _mesh_9_4_io_out_control_0_propagate;
	wire [4:0] _mesh_9_4_io_out_control_0_shift;
	wire [2:0] _mesh_9_4_io_out_id_0;
	wire _mesh_9_4_io_out_last_0;
	wire _mesh_9_4_io_out_valid_0;
	wire [31:0] _mesh_9_3_io_out_a_0;
	wire [31:0] _mesh_9_3_io_out_c_0;
	wire [31:0] _mesh_9_3_io_out_b_0;
	wire _mesh_9_3_io_out_control_0_dataflow;
	wire _mesh_9_3_io_out_control_0_propagate;
	wire [4:0] _mesh_9_3_io_out_control_0_shift;
	wire [2:0] _mesh_9_3_io_out_id_0;
	wire _mesh_9_3_io_out_last_0;
	wire _mesh_9_3_io_out_valid_0;
	wire [31:0] _mesh_9_2_io_out_a_0;
	wire [31:0] _mesh_9_2_io_out_c_0;
	wire [31:0] _mesh_9_2_io_out_b_0;
	wire _mesh_9_2_io_out_control_0_dataflow;
	wire _mesh_9_2_io_out_control_0_propagate;
	wire [4:0] _mesh_9_2_io_out_control_0_shift;
	wire [2:0] _mesh_9_2_io_out_id_0;
	wire _mesh_9_2_io_out_last_0;
	wire _mesh_9_2_io_out_valid_0;
	wire [31:0] _mesh_9_1_io_out_a_0;
	wire [31:0] _mesh_9_1_io_out_c_0;
	wire [31:0] _mesh_9_1_io_out_b_0;
	wire _mesh_9_1_io_out_control_0_dataflow;
	wire _mesh_9_1_io_out_control_0_propagate;
	wire [4:0] _mesh_9_1_io_out_control_0_shift;
	wire [2:0] _mesh_9_1_io_out_id_0;
	wire _mesh_9_1_io_out_last_0;
	wire _mesh_9_1_io_out_valid_0;
	wire [31:0] _mesh_9_0_io_out_a_0;
	wire [31:0] _mesh_9_0_io_out_c_0;
	wire [31:0] _mesh_9_0_io_out_b_0;
	wire _mesh_9_0_io_out_control_0_dataflow;
	wire _mesh_9_0_io_out_control_0_propagate;
	wire [4:0] _mesh_9_0_io_out_control_0_shift;
	wire [2:0] _mesh_9_0_io_out_id_0;
	wire _mesh_9_0_io_out_last_0;
	wire _mesh_9_0_io_out_valid_0;
	wire [31:0] _mesh_8_31_io_out_a_0;
	wire [31:0] _mesh_8_31_io_out_c_0;
	wire [31:0] _mesh_8_31_io_out_b_0;
	wire _mesh_8_31_io_out_control_0_dataflow;
	wire _mesh_8_31_io_out_control_0_propagate;
	wire [4:0] _mesh_8_31_io_out_control_0_shift;
	wire [2:0] _mesh_8_31_io_out_id_0;
	wire _mesh_8_31_io_out_last_0;
	wire _mesh_8_31_io_out_valid_0;
	wire [31:0] _mesh_8_30_io_out_a_0;
	wire [31:0] _mesh_8_30_io_out_c_0;
	wire [31:0] _mesh_8_30_io_out_b_0;
	wire _mesh_8_30_io_out_control_0_dataflow;
	wire _mesh_8_30_io_out_control_0_propagate;
	wire [4:0] _mesh_8_30_io_out_control_0_shift;
	wire [2:0] _mesh_8_30_io_out_id_0;
	wire _mesh_8_30_io_out_last_0;
	wire _mesh_8_30_io_out_valid_0;
	wire [31:0] _mesh_8_29_io_out_a_0;
	wire [31:0] _mesh_8_29_io_out_c_0;
	wire [31:0] _mesh_8_29_io_out_b_0;
	wire _mesh_8_29_io_out_control_0_dataflow;
	wire _mesh_8_29_io_out_control_0_propagate;
	wire [4:0] _mesh_8_29_io_out_control_0_shift;
	wire [2:0] _mesh_8_29_io_out_id_0;
	wire _mesh_8_29_io_out_last_0;
	wire _mesh_8_29_io_out_valid_0;
	wire [31:0] _mesh_8_28_io_out_a_0;
	wire [31:0] _mesh_8_28_io_out_c_0;
	wire [31:0] _mesh_8_28_io_out_b_0;
	wire _mesh_8_28_io_out_control_0_dataflow;
	wire _mesh_8_28_io_out_control_0_propagate;
	wire [4:0] _mesh_8_28_io_out_control_0_shift;
	wire [2:0] _mesh_8_28_io_out_id_0;
	wire _mesh_8_28_io_out_last_0;
	wire _mesh_8_28_io_out_valid_0;
	wire [31:0] _mesh_8_27_io_out_a_0;
	wire [31:0] _mesh_8_27_io_out_c_0;
	wire [31:0] _mesh_8_27_io_out_b_0;
	wire _mesh_8_27_io_out_control_0_dataflow;
	wire _mesh_8_27_io_out_control_0_propagate;
	wire [4:0] _mesh_8_27_io_out_control_0_shift;
	wire [2:0] _mesh_8_27_io_out_id_0;
	wire _mesh_8_27_io_out_last_0;
	wire _mesh_8_27_io_out_valid_0;
	wire [31:0] _mesh_8_26_io_out_a_0;
	wire [31:0] _mesh_8_26_io_out_c_0;
	wire [31:0] _mesh_8_26_io_out_b_0;
	wire _mesh_8_26_io_out_control_0_dataflow;
	wire _mesh_8_26_io_out_control_0_propagate;
	wire [4:0] _mesh_8_26_io_out_control_0_shift;
	wire [2:0] _mesh_8_26_io_out_id_0;
	wire _mesh_8_26_io_out_last_0;
	wire _mesh_8_26_io_out_valid_0;
	wire [31:0] _mesh_8_25_io_out_a_0;
	wire [31:0] _mesh_8_25_io_out_c_0;
	wire [31:0] _mesh_8_25_io_out_b_0;
	wire _mesh_8_25_io_out_control_0_dataflow;
	wire _mesh_8_25_io_out_control_0_propagate;
	wire [4:0] _mesh_8_25_io_out_control_0_shift;
	wire [2:0] _mesh_8_25_io_out_id_0;
	wire _mesh_8_25_io_out_last_0;
	wire _mesh_8_25_io_out_valid_0;
	wire [31:0] _mesh_8_24_io_out_a_0;
	wire [31:0] _mesh_8_24_io_out_c_0;
	wire [31:0] _mesh_8_24_io_out_b_0;
	wire _mesh_8_24_io_out_control_0_dataflow;
	wire _mesh_8_24_io_out_control_0_propagate;
	wire [4:0] _mesh_8_24_io_out_control_0_shift;
	wire [2:0] _mesh_8_24_io_out_id_0;
	wire _mesh_8_24_io_out_last_0;
	wire _mesh_8_24_io_out_valid_0;
	wire [31:0] _mesh_8_23_io_out_a_0;
	wire [31:0] _mesh_8_23_io_out_c_0;
	wire [31:0] _mesh_8_23_io_out_b_0;
	wire _mesh_8_23_io_out_control_0_dataflow;
	wire _mesh_8_23_io_out_control_0_propagate;
	wire [4:0] _mesh_8_23_io_out_control_0_shift;
	wire [2:0] _mesh_8_23_io_out_id_0;
	wire _mesh_8_23_io_out_last_0;
	wire _mesh_8_23_io_out_valid_0;
	wire [31:0] _mesh_8_22_io_out_a_0;
	wire [31:0] _mesh_8_22_io_out_c_0;
	wire [31:0] _mesh_8_22_io_out_b_0;
	wire _mesh_8_22_io_out_control_0_dataflow;
	wire _mesh_8_22_io_out_control_0_propagate;
	wire [4:0] _mesh_8_22_io_out_control_0_shift;
	wire [2:0] _mesh_8_22_io_out_id_0;
	wire _mesh_8_22_io_out_last_0;
	wire _mesh_8_22_io_out_valid_0;
	wire [31:0] _mesh_8_21_io_out_a_0;
	wire [31:0] _mesh_8_21_io_out_c_0;
	wire [31:0] _mesh_8_21_io_out_b_0;
	wire _mesh_8_21_io_out_control_0_dataflow;
	wire _mesh_8_21_io_out_control_0_propagate;
	wire [4:0] _mesh_8_21_io_out_control_0_shift;
	wire [2:0] _mesh_8_21_io_out_id_0;
	wire _mesh_8_21_io_out_last_0;
	wire _mesh_8_21_io_out_valid_0;
	wire [31:0] _mesh_8_20_io_out_a_0;
	wire [31:0] _mesh_8_20_io_out_c_0;
	wire [31:0] _mesh_8_20_io_out_b_0;
	wire _mesh_8_20_io_out_control_0_dataflow;
	wire _mesh_8_20_io_out_control_0_propagate;
	wire [4:0] _mesh_8_20_io_out_control_0_shift;
	wire [2:0] _mesh_8_20_io_out_id_0;
	wire _mesh_8_20_io_out_last_0;
	wire _mesh_8_20_io_out_valid_0;
	wire [31:0] _mesh_8_19_io_out_a_0;
	wire [31:0] _mesh_8_19_io_out_c_0;
	wire [31:0] _mesh_8_19_io_out_b_0;
	wire _mesh_8_19_io_out_control_0_dataflow;
	wire _mesh_8_19_io_out_control_0_propagate;
	wire [4:0] _mesh_8_19_io_out_control_0_shift;
	wire [2:0] _mesh_8_19_io_out_id_0;
	wire _mesh_8_19_io_out_last_0;
	wire _mesh_8_19_io_out_valid_0;
	wire [31:0] _mesh_8_18_io_out_a_0;
	wire [31:0] _mesh_8_18_io_out_c_0;
	wire [31:0] _mesh_8_18_io_out_b_0;
	wire _mesh_8_18_io_out_control_0_dataflow;
	wire _mesh_8_18_io_out_control_0_propagate;
	wire [4:0] _mesh_8_18_io_out_control_0_shift;
	wire [2:0] _mesh_8_18_io_out_id_0;
	wire _mesh_8_18_io_out_last_0;
	wire _mesh_8_18_io_out_valid_0;
	wire [31:0] _mesh_8_17_io_out_a_0;
	wire [31:0] _mesh_8_17_io_out_c_0;
	wire [31:0] _mesh_8_17_io_out_b_0;
	wire _mesh_8_17_io_out_control_0_dataflow;
	wire _mesh_8_17_io_out_control_0_propagate;
	wire [4:0] _mesh_8_17_io_out_control_0_shift;
	wire [2:0] _mesh_8_17_io_out_id_0;
	wire _mesh_8_17_io_out_last_0;
	wire _mesh_8_17_io_out_valid_0;
	wire [31:0] _mesh_8_16_io_out_a_0;
	wire [31:0] _mesh_8_16_io_out_c_0;
	wire [31:0] _mesh_8_16_io_out_b_0;
	wire _mesh_8_16_io_out_control_0_dataflow;
	wire _mesh_8_16_io_out_control_0_propagate;
	wire [4:0] _mesh_8_16_io_out_control_0_shift;
	wire [2:0] _mesh_8_16_io_out_id_0;
	wire _mesh_8_16_io_out_last_0;
	wire _mesh_8_16_io_out_valid_0;
	wire [31:0] _mesh_8_15_io_out_a_0;
	wire [31:0] _mesh_8_15_io_out_c_0;
	wire [31:0] _mesh_8_15_io_out_b_0;
	wire _mesh_8_15_io_out_control_0_dataflow;
	wire _mesh_8_15_io_out_control_0_propagate;
	wire [4:0] _mesh_8_15_io_out_control_0_shift;
	wire [2:0] _mesh_8_15_io_out_id_0;
	wire _mesh_8_15_io_out_last_0;
	wire _mesh_8_15_io_out_valid_0;
	wire [31:0] _mesh_8_14_io_out_a_0;
	wire [31:0] _mesh_8_14_io_out_c_0;
	wire [31:0] _mesh_8_14_io_out_b_0;
	wire _mesh_8_14_io_out_control_0_dataflow;
	wire _mesh_8_14_io_out_control_0_propagate;
	wire [4:0] _mesh_8_14_io_out_control_0_shift;
	wire [2:0] _mesh_8_14_io_out_id_0;
	wire _mesh_8_14_io_out_last_0;
	wire _mesh_8_14_io_out_valid_0;
	wire [31:0] _mesh_8_13_io_out_a_0;
	wire [31:0] _mesh_8_13_io_out_c_0;
	wire [31:0] _mesh_8_13_io_out_b_0;
	wire _mesh_8_13_io_out_control_0_dataflow;
	wire _mesh_8_13_io_out_control_0_propagate;
	wire [4:0] _mesh_8_13_io_out_control_0_shift;
	wire [2:0] _mesh_8_13_io_out_id_0;
	wire _mesh_8_13_io_out_last_0;
	wire _mesh_8_13_io_out_valid_0;
	wire [31:0] _mesh_8_12_io_out_a_0;
	wire [31:0] _mesh_8_12_io_out_c_0;
	wire [31:0] _mesh_8_12_io_out_b_0;
	wire _mesh_8_12_io_out_control_0_dataflow;
	wire _mesh_8_12_io_out_control_0_propagate;
	wire [4:0] _mesh_8_12_io_out_control_0_shift;
	wire [2:0] _mesh_8_12_io_out_id_0;
	wire _mesh_8_12_io_out_last_0;
	wire _mesh_8_12_io_out_valid_0;
	wire [31:0] _mesh_8_11_io_out_a_0;
	wire [31:0] _mesh_8_11_io_out_c_0;
	wire [31:0] _mesh_8_11_io_out_b_0;
	wire _mesh_8_11_io_out_control_0_dataflow;
	wire _mesh_8_11_io_out_control_0_propagate;
	wire [4:0] _mesh_8_11_io_out_control_0_shift;
	wire [2:0] _mesh_8_11_io_out_id_0;
	wire _mesh_8_11_io_out_last_0;
	wire _mesh_8_11_io_out_valid_0;
	wire [31:0] _mesh_8_10_io_out_a_0;
	wire [31:0] _mesh_8_10_io_out_c_0;
	wire [31:0] _mesh_8_10_io_out_b_0;
	wire _mesh_8_10_io_out_control_0_dataflow;
	wire _mesh_8_10_io_out_control_0_propagate;
	wire [4:0] _mesh_8_10_io_out_control_0_shift;
	wire [2:0] _mesh_8_10_io_out_id_0;
	wire _mesh_8_10_io_out_last_0;
	wire _mesh_8_10_io_out_valid_0;
	wire [31:0] _mesh_8_9_io_out_a_0;
	wire [31:0] _mesh_8_9_io_out_c_0;
	wire [31:0] _mesh_8_9_io_out_b_0;
	wire _mesh_8_9_io_out_control_0_dataflow;
	wire _mesh_8_9_io_out_control_0_propagate;
	wire [4:0] _mesh_8_9_io_out_control_0_shift;
	wire [2:0] _mesh_8_9_io_out_id_0;
	wire _mesh_8_9_io_out_last_0;
	wire _mesh_8_9_io_out_valid_0;
	wire [31:0] _mesh_8_8_io_out_a_0;
	wire [31:0] _mesh_8_8_io_out_c_0;
	wire [31:0] _mesh_8_8_io_out_b_0;
	wire _mesh_8_8_io_out_control_0_dataflow;
	wire _mesh_8_8_io_out_control_0_propagate;
	wire [4:0] _mesh_8_8_io_out_control_0_shift;
	wire [2:0] _mesh_8_8_io_out_id_0;
	wire _mesh_8_8_io_out_last_0;
	wire _mesh_8_8_io_out_valid_0;
	wire [31:0] _mesh_8_7_io_out_a_0;
	wire [31:0] _mesh_8_7_io_out_c_0;
	wire [31:0] _mesh_8_7_io_out_b_0;
	wire _mesh_8_7_io_out_control_0_dataflow;
	wire _mesh_8_7_io_out_control_0_propagate;
	wire [4:0] _mesh_8_7_io_out_control_0_shift;
	wire [2:0] _mesh_8_7_io_out_id_0;
	wire _mesh_8_7_io_out_last_0;
	wire _mesh_8_7_io_out_valid_0;
	wire [31:0] _mesh_8_6_io_out_a_0;
	wire [31:0] _mesh_8_6_io_out_c_0;
	wire [31:0] _mesh_8_6_io_out_b_0;
	wire _mesh_8_6_io_out_control_0_dataflow;
	wire _mesh_8_6_io_out_control_0_propagate;
	wire [4:0] _mesh_8_6_io_out_control_0_shift;
	wire [2:0] _mesh_8_6_io_out_id_0;
	wire _mesh_8_6_io_out_last_0;
	wire _mesh_8_6_io_out_valid_0;
	wire [31:0] _mesh_8_5_io_out_a_0;
	wire [31:0] _mesh_8_5_io_out_c_0;
	wire [31:0] _mesh_8_5_io_out_b_0;
	wire _mesh_8_5_io_out_control_0_dataflow;
	wire _mesh_8_5_io_out_control_0_propagate;
	wire [4:0] _mesh_8_5_io_out_control_0_shift;
	wire [2:0] _mesh_8_5_io_out_id_0;
	wire _mesh_8_5_io_out_last_0;
	wire _mesh_8_5_io_out_valid_0;
	wire [31:0] _mesh_8_4_io_out_a_0;
	wire [31:0] _mesh_8_4_io_out_c_0;
	wire [31:0] _mesh_8_4_io_out_b_0;
	wire _mesh_8_4_io_out_control_0_dataflow;
	wire _mesh_8_4_io_out_control_0_propagate;
	wire [4:0] _mesh_8_4_io_out_control_0_shift;
	wire [2:0] _mesh_8_4_io_out_id_0;
	wire _mesh_8_4_io_out_last_0;
	wire _mesh_8_4_io_out_valid_0;
	wire [31:0] _mesh_8_3_io_out_a_0;
	wire [31:0] _mesh_8_3_io_out_c_0;
	wire [31:0] _mesh_8_3_io_out_b_0;
	wire _mesh_8_3_io_out_control_0_dataflow;
	wire _mesh_8_3_io_out_control_0_propagate;
	wire [4:0] _mesh_8_3_io_out_control_0_shift;
	wire [2:0] _mesh_8_3_io_out_id_0;
	wire _mesh_8_3_io_out_last_0;
	wire _mesh_8_3_io_out_valid_0;
	wire [31:0] _mesh_8_2_io_out_a_0;
	wire [31:0] _mesh_8_2_io_out_c_0;
	wire [31:0] _mesh_8_2_io_out_b_0;
	wire _mesh_8_2_io_out_control_0_dataflow;
	wire _mesh_8_2_io_out_control_0_propagate;
	wire [4:0] _mesh_8_2_io_out_control_0_shift;
	wire [2:0] _mesh_8_2_io_out_id_0;
	wire _mesh_8_2_io_out_last_0;
	wire _mesh_8_2_io_out_valid_0;
	wire [31:0] _mesh_8_1_io_out_a_0;
	wire [31:0] _mesh_8_1_io_out_c_0;
	wire [31:0] _mesh_8_1_io_out_b_0;
	wire _mesh_8_1_io_out_control_0_dataflow;
	wire _mesh_8_1_io_out_control_0_propagate;
	wire [4:0] _mesh_8_1_io_out_control_0_shift;
	wire [2:0] _mesh_8_1_io_out_id_0;
	wire _mesh_8_1_io_out_last_0;
	wire _mesh_8_1_io_out_valid_0;
	wire [31:0] _mesh_8_0_io_out_a_0;
	wire [31:0] _mesh_8_0_io_out_c_0;
	wire [31:0] _mesh_8_0_io_out_b_0;
	wire _mesh_8_0_io_out_control_0_dataflow;
	wire _mesh_8_0_io_out_control_0_propagate;
	wire [4:0] _mesh_8_0_io_out_control_0_shift;
	wire [2:0] _mesh_8_0_io_out_id_0;
	wire _mesh_8_0_io_out_last_0;
	wire _mesh_8_0_io_out_valid_0;
	wire [31:0] _mesh_7_31_io_out_a_0;
	wire [31:0] _mesh_7_31_io_out_c_0;
	wire [31:0] _mesh_7_31_io_out_b_0;
	wire _mesh_7_31_io_out_control_0_dataflow;
	wire _mesh_7_31_io_out_control_0_propagate;
	wire [4:0] _mesh_7_31_io_out_control_0_shift;
	wire [2:0] _mesh_7_31_io_out_id_0;
	wire _mesh_7_31_io_out_last_0;
	wire _mesh_7_31_io_out_valid_0;
	wire [31:0] _mesh_7_30_io_out_a_0;
	wire [31:0] _mesh_7_30_io_out_c_0;
	wire [31:0] _mesh_7_30_io_out_b_0;
	wire _mesh_7_30_io_out_control_0_dataflow;
	wire _mesh_7_30_io_out_control_0_propagate;
	wire [4:0] _mesh_7_30_io_out_control_0_shift;
	wire [2:0] _mesh_7_30_io_out_id_0;
	wire _mesh_7_30_io_out_last_0;
	wire _mesh_7_30_io_out_valid_0;
	wire [31:0] _mesh_7_29_io_out_a_0;
	wire [31:0] _mesh_7_29_io_out_c_0;
	wire [31:0] _mesh_7_29_io_out_b_0;
	wire _mesh_7_29_io_out_control_0_dataflow;
	wire _mesh_7_29_io_out_control_0_propagate;
	wire [4:0] _mesh_7_29_io_out_control_0_shift;
	wire [2:0] _mesh_7_29_io_out_id_0;
	wire _mesh_7_29_io_out_last_0;
	wire _mesh_7_29_io_out_valid_0;
	wire [31:0] _mesh_7_28_io_out_a_0;
	wire [31:0] _mesh_7_28_io_out_c_0;
	wire [31:0] _mesh_7_28_io_out_b_0;
	wire _mesh_7_28_io_out_control_0_dataflow;
	wire _mesh_7_28_io_out_control_0_propagate;
	wire [4:0] _mesh_7_28_io_out_control_0_shift;
	wire [2:0] _mesh_7_28_io_out_id_0;
	wire _mesh_7_28_io_out_last_0;
	wire _mesh_7_28_io_out_valid_0;
	wire [31:0] _mesh_7_27_io_out_a_0;
	wire [31:0] _mesh_7_27_io_out_c_0;
	wire [31:0] _mesh_7_27_io_out_b_0;
	wire _mesh_7_27_io_out_control_0_dataflow;
	wire _mesh_7_27_io_out_control_0_propagate;
	wire [4:0] _mesh_7_27_io_out_control_0_shift;
	wire [2:0] _mesh_7_27_io_out_id_0;
	wire _mesh_7_27_io_out_last_0;
	wire _mesh_7_27_io_out_valid_0;
	wire [31:0] _mesh_7_26_io_out_a_0;
	wire [31:0] _mesh_7_26_io_out_c_0;
	wire [31:0] _mesh_7_26_io_out_b_0;
	wire _mesh_7_26_io_out_control_0_dataflow;
	wire _mesh_7_26_io_out_control_0_propagate;
	wire [4:0] _mesh_7_26_io_out_control_0_shift;
	wire [2:0] _mesh_7_26_io_out_id_0;
	wire _mesh_7_26_io_out_last_0;
	wire _mesh_7_26_io_out_valid_0;
	wire [31:0] _mesh_7_25_io_out_a_0;
	wire [31:0] _mesh_7_25_io_out_c_0;
	wire [31:0] _mesh_7_25_io_out_b_0;
	wire _mesh_7_25_io_out_control_0_dataflow;
	wire _mesh_7_25_io_out_control_0_propagate;
	wire [4:0] _mesh_7_25_io_out_control_0_shift;
	wire [2:0] _mesh_7_25_io_out_id_0;
	wire _mesh_7_25_io_out_last_0;
	wire _mesh_7_25_io_out_valid_0;
	wire [31:0] _mesh_7_24_io_out_a_0;
	wire [31:0] _mesh_7_24_io_out_c_0;
	wire [31:0] _mesh_7_24_io_out_b_0;
	wire _mesh_7_24_io_out_control_0_dataflow;
	wire _mesh_7_24_io_out_control_0_propagate;
	wire [4:0] _mesh_7_24_io_out_control_0_shift;
	wire [2:0] _mesh_7_24_io_out_id_0;
	wire _mesh_7_24_io_out_last_0;
	wire _mesh_7_24_io_out_valid_0;
	wire [31:0] _mesh_7_23_io_out_a_0;
	wire [31:0] _mesh_7_23_io_out_c_0;
	wire [31:0] _mesh_7_23_io_out_b_0;
	wire _mesh_7_23_io_out_control_0_dataflow;
	wire _mesh_7_23_io_out_control_0_propagate;
	wire [4:0] _mesh_7_23_io_out_control_0_shift;
	wire [2:0] _mesh_7_23_io_out_id_0;
	wire _mesh_7_23_io_out_last_0;
	wire _mesh_7_23_io_out_valid_0;
	wire [31:0] _mesh_7_22_io_out_a_0;
	wire [31:0] _mesh_7_22_io_out_c_0;
	wire [31:0] _mesh_7_22_io_out_b_0;
	wire _mesh_7_22_io_out_control_0_dataflow;
	wire _mesh_7_22_io_out_control_0_propagate;
	wire [4:0] _mesh_7_22_io_out_control_0_shift;
	wire [2:0] _mesh_7_22_io_out_id_0;
	wire _mesh_7_22_io_out_last_0;
	wire _mesh_7_22_io_out_valid_0;
	wire [31:0] _mesh_7_21_io_out_a_0;
	wire [31:0] _mesh_7_21_io_out_c_0;
	wire [31:0] _mesh_7_21_io_out_b_0;
	wire _mesh_7_21_io_out_control_0_dataflow;
	wire _mesh_7_21_io_out_control_0_propagate;
	wire [4:0] _mesh_7_21_io_out_control_0_shift;
	wire [2:0] _mesh_7_21_io_out_id_0;
	wire _mesh_7_21_io_out_last_0;
	wire _mesh_7_21_io_out_valid_0;
	wire [31:0] _mesh_7_20_io_out_a_0;
	wire [31:0] _mesh_7_20_io_out_c_0;
	wire [31:0] _mesh_7_20_io_out_b_0;
	wire _mesh_7_20_io_out_control_0_dataflow;
	wire _mesh_7_20_io_out_control_0_propagate;
	wire [4:0] _mesh_7_20_io_out_control_0_shift;
	wire [2:0] _mesh_7_20_io_out_id_0;
	wire _mesh_7_20_io_out_last_0;
	wire _mesh_7_20_io_out_valid_0;
	wire [31:0] _mesh_7_19_io_out_a_0;
	wire [31:0] _mesh_7_19_io_out_c_0;
	wire [31:0] _mesh_7_19_io_out_b_0;
	wire _mesh_7_19_io_out_control_0_dataflow;
	wire _mesh_7_19_io_out_control_0_propagate;
	wire [4:0] _mesh_7_19_io_out_control_0_shift;
	wire [2:0] _mesh_7_19_io_out_id_0;
	wire _mesh_7_19_io_out_last_0;
	wire _mesh_7_19_io_out_valid_0;
	wire [31:0] _mesh_7_18_io_out_a_0;
	wire [31:0] _mesh_7_18_io_out_c_0;
	wire [31:0] _mesh_7_18_io_out_b_0;
	wire _mesh_7_18_io_out_control_0_dataflow;
	wire _mesh_7_18_io_out_control_0_propagate;
	wire [4:0] _mesh_7_18_io_out_control_0_shift;
	wire [2:0] _mesh_7_18_io_out_id_0;
	wire _mesh_7_18_io_out_last_0;
	wire _mesh_7_18_io_out_valid_0;
	wire [31:0] _mesh_7_17_io_out_a_0;
	wire [31:0] _mesh_7_17_io_out_c_0;
	wire [31:0] _mesh_7_17_io_out_b_0;
	wire _mesh_7_17_io_out_control_0_dataflow;
	wire _mesh_7_17_io_out_control_0_propagate;
	wire [4:0] _mesh_7_17_io_out_control_0_shift;
	wire [2:0] _mesh_7_17_io_out_id_0;
	wire _mesh_7_17_io_out_last_0;
	wire _mesh_7_17_io_out_valid_0;
	wire [31:0] _mesh_7_16_io_out_a_0;
	wire [31:0] _mesh_7_16_io_out_c_0;
	wire [31:0] _mesh_7_16_io_out_b_0;
	wire _mesh_7_16_io_out_control_0_dataflow;
	wire _mesh_7_16_io_out_control_0_propagate;
	wire [4:0] _mesh_7_16_io_out_control_0_shift;
	wire [2:0] _mesh_7_16_io_out_id_0;
	wire _mesh_7_16_io_out_last_0;
	wire _mesh_7_16_io_out_valid_0;
	wire [31:0] _mesh_7_15_io_out_a_0;
	wire [31:0] _mesh_7_15_io_out_c_0;
	wire [31:0] _mesh_7_15_io_out_b_0;
	wire _mesh_7_15_io_out_control_0_dataflow;
	wire _mesh_7_15_io_out_control_0_propagate;
	wire [4:0] _mesh_7_15_io_out_control_0_shift;
	wire [2:0] _mesh_7_15_io_out_id_0;
	wire _mesh_7_15_io_out_last_0;
	wire _mesh_7_15_io_out_valid_0;
	wire [31:0] _mesh_7_14_io_out_a_0;
	wire [31:0] _mesh_7_14_io_out_c_0;
	wire [31:0] _mesh_7_14_io_out_b_0;
	wire _mesh_7_14_io_out_control_0_dataflow;
	wire _mesh_7_14_io_out_control_0_propagate;
	wire [4:0] _mesh_7_14_io_out_control_0_shift;
	wire [2:0] _mesh_7_14_io_out_id_0;
	wire _mesh_7_14_io_out_last_0;
	wire _mesh_7_14_io_out_valid_0;
	wire [31:0] _mesh_7_13_io_out_a_0;
	wire [31:0] _mesh_7_13_io_out_c_0;
	wire [31:0] _mesh_7_13_io_out_b_0;
	wire _mesh_7_13_io_out_control_0_dataflow;
	wire _mesh_7_13_io_out_control_0_propagate;
	wire [4:0] _mesh_7_13_io_out_control_0_shift;
	wire [2:0] _mesh_7_13_io_out_id_0;
	wire _mesh_7_13_io_out_last_0;
	wire _mesh_7_13_io_out_valid_0;
	wire [31:0] _mesh_7_12_io_out_a_0;
	wire [31:0] _mesh_7_12_io_out_c_0;
	wire [31:0] _mesh_7_12_io_out_b_0;
	wire _mesh_7_12_io_out_control_0_dataflow;
	wire _mesh_7_12_io_out_control_0_propagate;
	wire [4:0] _mesh_7_12_io_out_control_0_shift;
	wire [2:0] _mesh_7_12_io_out_id_0;
	wire _mesh_7_12_io_out_last_0;
	wire _mesh_7_12_io_out_valid_0;
	wire [31:0] _mesh_7_11_io_out_a_0;
	wire [31:0] _mesh_7_11_io_out_c_0;
	wire [31:0] _mesh_7_11_io_out_b_0;
	wire _mesh_7_11_io_out_control_0_dataflow;
	wire _mesh_7_11_io_out_control_0_propagate;
	wire [4:0] _mesh_7_11_io_out_control_0_shift;
	wire [2:0] _mesh_7_11_io_out_id_0;
	wire _mesh_7_11_io_out_last_0;
	wire _mesh_7_11_io_out_valid_0;
	wire [31:0] _mesh_7_10_io_out_a_0;
	wire [31:0] _mesh_7_10_io_out_c_0;
	wire [31:0] _mesh_7_10_io_out_b_0;
	wire _mesh_7_10_io_out_control_0_dataflow;
	wire _mesh_7_10_io_out_control_0_propagate;
	wire [4:0] _mesh_7_10_io_out_control_0_shift;
	wire [2:0] _mesh_7_10_io_out_id_0;
	wire _mesh_7_10_io_out_last_0;
	wire _mesh_7_10_io_out_valid_0;
	wire [31:0] _mesh_7_9_io_out_a_0;
	wire [31:0] _mesh_7_9_io_out_c_0;
	wire [31:0] _mesh_7_9_io_out_b_0;
	wire _mesh_7_9_io_out_control_0_dataflow;
	wire _mesh_7_9_io_out_control_0_propagate;
	wire [4:0] _mesh_7_9_io_out_control_0_shift;
	wire [2:0] _mesh_7_9_io_out_id_0;
	wire _mesh_7_9_io_out_last_0;
	wire _mesh_7_9_io_out_valid_0;
	wire [31:0] _mesh_7_8_io_out_a_0;
	wire [31:0] _mesh_7_8_io_out_c_0;
	wire [31:0] _mesh_7_8_io_out_b_0;
	wire _mesh_7_8_io_out_control_0_dataflow;
	wire _mesh_7_8_io_out_control_0_propagate;
	wire [4:0] _mesh_7_8_io_out_control_0_shift;
	wire [2:0] _mesh_7_8_io_out_id_0;
	wire _mesh_7_8_io_out_last_0;
	wire _mesh_7_8_io_out_valid_0;
	wire [31:0] _mesh_7_7_io_out_a_0;
	wire [31:0] _mesh_7_7_io_out_c_0;
	wire [31:0] _mesh_7_7_io_out_b_0;
	wire _mesh_7_7_io_out_control_0_dataflow;
	wire _mesh_7_7_io_out_control_0_propagate;
	wire [4:0] _mesh_7_7_io_out_control_0_shift;
	wire [2:0] _mesh_7_7_io_out_id_0;
	wire _mesh_7_7_io_out_last_0;
	wire _mesh_7_7_io_out_valid_0;
	wire [31:0] _mesh_7_6_io_out_a_0;
	wire [31:0] _mesh_7_6_io_out_c_0;
	wire [31:0] _mesh_7_6_io_out_b_0;
	wire _mesh_7_6_io_out_control_0_dataflow;
	wire _mesh_7_6_io_out_control_0_propagate;
	wire [4:0] _mesh_7_6_io_out_control_0_shift;
	wire [2:0] _mesh_7_6_io_out_id_0;
	wire _mesh_7_6_io_out_last_0;
	wire _mesh_7_6_io_out_valid_0;
	wire [31:0] _mesh_7_5_io_out_a_0;
	wire [31:0] _mesh_7_5_io_out_c_0;
	wire [31:0] _mesh_7_5_io_out_b_0;
	wire _mesh_7_5_io_out_control_0_dataflow;
	wire _mesh_7_5_io_out_control_0_propagate;
	wire [4:0] _mesh_7_5_io_out_control_0_shift;
	wire [2:0] _mesh_7_5_io_out_id_0;
	wire _mesh_7_5_io_out_last_0;
	wire _mesh_7_5_io_out_valid_0;
	wire [31:0] _mesh_7_4_io_out_a_0;
	wire [31:0] _mesh_7_4_io_out_c_0;
	wire [31:0] _mesh_7_4_io_out_b_0;
	wire _mesh_7_4_io_out_control_0_dataflow;
	wire _mesh_7_4_io_out_control_0_propagate;
	wire [4:0] _mesh_7_4_io_out_control_0_shift;
	wire [2:0] _mesh_7_4_io_out_id_0;
	wire _mesh_7_4_io_out_last_0;
	wire _mesh_7_4_io_out_valid_0;
	wire [31:0] _mesh_7_3_io_out_a_0;
	wire [31:0] _mesh_7_3_io_out_c_0;
	wire [31:0] _mesh_7_3_io_out_b_0;
	wire _mesh_7_3_io_out_control_0_dataflow;
	wire _mesh_7_3_io_out_control_0_propagate;
	wire [4:0] _mesh_7_3_io_out_control_0_shift;
	wire [2:0] _mesh_7_3_io_out_id_0;
	wire _mesh_7_3_io_out_last_0;
	wire _mesh_7_3_io_out_valid_0;
	wire [31:0] _mesh_7_2_io_out_a_0;
	wire [31:0] _mesh_7_2_io_out_c_0;
	wire [31:0] _mesh_7_2_io_out_b_0;
	wire _mesh_7_2_io_out_control_0_dataflow;
	wire _mesh_7_2_io_out_control_0_propagate;
	wire [4:0] _mesh_7_2_io_out_control_0_shift;
	wire [2:0] _mesh_7_2_io_out_id_0;
	wire _mesh_7_2_io_out_last_0;
	wire _mesh_7_2_io_out_valid_0;
	wire [31:0] _mesh_7_1_io_out_a_0;
	wire [31:0] _mesh_7_1_io_out_c_0;
	wire [31:0] _mesh_7_1_io_out_b_0;
	wire _mesh_7_1_io_out_control_0_dataflow;
	wire _mesh_7_1_io_out_control_0_propagate;
	wire [4:0] _mesh_7_1_io_out_control_0_shift;
	wire [2:0] _mesh_7_1_io_out_id_0;
	wire _mesh_7_1_io_out_last_0;
	wire _mesh_7_1_io_out_valid_0;
	wire [31:0] _mesh_7_0_io_out_a_0;
	wire [31:0] _mesh_7_0_io_out_c_0;
	wire [31:0] _mesh_7_0_io_out_b_0;
	wire _mesh_7_0_io_out_control_0_dataflow;
	wire _mesh_7_0_io_out_control_0_propagate;
	wire [4:0] _mesh_7_0_io_out_control_0_shift;
	wire [2:0] _mesh_7_0_io_out_id_0;
	wire _mesh_7_0_io_out_last_0;
	wire _mesh_7_0_io_out_valid_0;
	wire [31:0] _mesh_6_31_io_out_a_0;
	wire [31:0] _mesh_6_31_io_out_c_0;
	wire [31:0] _mesh_6_31_io_out_b_0;
	wire _mesh_6_31_io_out_control_0_dataflow;
	wire _mesh_6_31_io_out_control_0_propagate;
	wire [4:0] _mesh_6_31_io_out_control_0_shift;
	wire [2:0] _mesh_6_31_io_out_id_0;
	wire _mesh_6_31_io_out_last_0;
	wire _mesh_6_31_io_out_valid_0;
	wire [31:0] _mesh_6_30_io_out_a_0;
	wire [31:0] _mesh_6_30_io_out_c_0;
	wire [31:0] _mesh_6_30_io_out_b_0;
	wire _mesh_6_30_io_out_control_0_dataflow;
	wire _mesh_6_30_io_out_control_0_propagate;
	wire [4:0] _mesh_6_30_io_out_control_0_shift;
	wire [2:0] _mesh_6_30_io_out_id_0;
	wire _mesh_6_30_io_out_last_0;
	wire _mesh_6_30_io_out_valid_0;
	wire [31:0] _mesh_6_29_io_out_a_0;
	wire [31:0] _mesh_6_29_io_out_c_0;
	wire [31:0] _mesh_6_29_io_out_b_0;
	wire _mesh_6_29_io_out_control_0_dataflow;
	wire _mesh_6_29_io_out_control_0_propagate;
	wire [4:0] _mesh_6_29_io_out_control_0_shift;
	wire [2:0] _mesh_6_29_io_out_id_0;
	wire _mesh_6_29_io_out_last_0;
	wire _mesh_6_29_io_out_valid_0;
	wire [31:0] _mesh_6_28_io_out_a_0;
	wire [31:0] _mesh_6_28_io_out_c_0;
	wire [31:0] _mesh_6_28_io_out_b_0;
	wire _mesh_6_28_io_out_control_0_dataflow;
	wire _mesh_6_28_io_out_control_0_propagate;
	wire [4:0] _mesh_6_28_io_out_control_0_shift;
	wire [2:0] _mesh_6_28_io_out_id_0;
	wire _mesh_6_28_io_out_last_0;
	wire _mesh_6_28_io_out_valid_0;
	wire [31:0] _mesh_6_27_io_out_a_0;
	wire [31:0] _mesh_6_27_io_out_c_0;
	wire [31:0] _mesh_6_27_io_out_b_0;
	wire _mesh_6_27_io_out_control_0_dataflow;
	wire _mesh_6_27_io_out_control_0_propagate;
	wire [4:0] _mesh_6_27_io_out_control_0_shift;
	wire [2:0] _mesh_6_27_io_out_id_0;
	wire _mesh_6_27_io_out_last_0;
	wire _mesh_6_27_io_out_valid_0;
	wire [31:0] _mesh_6_26_io_out_a_0;
	wire [31:0] _mesh_6_26_io_out_c_0;
	wire [31:0] _mesh_6_26_io_out_b_0;
	wire _mesh_6_26_io_out_control_0_dataflow;
	wire _mesh_6_26_io_out_control_0_propagate;
	wire [4:0] _mesh_6_26_io_out_control_0_shift;
	wire [2:0] _mesh_6_26_io_out_id_0;
	wire _mesh_6_26_io_out_last_0;
	wire _mesh_6_26_io_out_valid_0;
	wire [31:0] _mesh_6_25_io_out_a_0;
	wire [31:0] _mesh_6_25_io_out_c_0;
	wire [31:0] _mesh_6_25_io_out_b_0;
	wire _mesh_6_25_io_out_control_0_dataflow;
	wire _mesh_6_25_io_out_control_0_propagate;
	wire [4:0] _mesh_6_25_io_out_control_0_shift;
	wire [2:0] _mesh_6_25_io_out_id_0;
	wire _mesh_6_25_io_out_last_0;
	wire _mesh_6_25_io_out_valid_0;
	wire [31:0] _mesh_6_24_io_out_a_0;
	wire [31:0] _mesh_6_24_io_out_c_0;
	wire [31:0] _mesh_6_24_io_out_b_0;
	wire _mesh_6_24_io_out_control_0_dataflow;
	wire _mesh_6_24_io_out_control_0_propagate;
	wire [4:0] _mesh_6_24_io_out_control_0_shift;
	wire [2:0] _mesh_6_24_io_out_id_0;
	wire _mesh_6_24_io_out_last_0;
	wire _mesh_6_24_io_out_valid_0;
	wire [31:0] _mesh_6_23_io_out_a_0;
	wire [31:0] _mesh_6_23_io_out_c_0;
	wire [31:0] _mesh_6_23_io_out_b_0;
	wire _mesh_6_23_io_out_control_0_dataflow;
	wire _mesh_6_23_io_out_control_0_propagate;
	wire [4:0] _mesh_6_23_io_out_control_0_shift;
	wire [2:0] _mesh_6_23_io_out_id_0;
	wire _mesh_6_23_io_out_last_0;
	wire _mesh_6_23_io_out_valid_0;
	wire [31:0] _mesh_6_22_io_out_a_0;
	wire [31:0] _mesh_6_22_io_out_c_0;
	wire [31:0] _mesh_6_22_io_out_b_0;
	wire _mesh_6_22_io_out_control_0_dataflow;
	wire _mesh_6_22_io_out_control_0_propagate;
	wire [4:0] _mesh_6_22_io_out_control_0_shift;
	wire [2:0] _mesh_6_22_io_out_id_0;
	wire _mesh_6_22_io_out_last_0;
	wire _mesh_6_22_io_out_valid_0;
	wire [31:0] _mesh_6_21_io_out_a_0;
	wire [31:0] _mesh_6_21_io_out_c_0;
	wire [31:0] _mesh_6_21_io_out_b_0;
	wire _mesh_6_21_io_out_control_0_dataflow;
	wire _mesh_6_21_io_out_control_0_propagate;
	wire [4:0] _mesh_6_21_io_out_control_0_shift;
	wire [2:0] _mesh_6_21_io_out_id_0;
	wire _mesh_6_21_io_out_last_0;
	wire _mesh_6_21_io_out_valid_0;
	wire [31:0] _mesh_6_20_io_out_a_0;
	wire [31:0] _mesh_6_20_io_out_c_0;
	wire [31:0] _mesh_6_20_io_out_b_0;
	wire _mesh_6_20_io_out_control_0_dataflow;
	wire _mesh_6_20_io_out_control_0_propagate;
	wire [4:0] _mesh_6_20_io_out_control_0_shift;
	wire [2:0] _mesh_6_20_io_out_id_0;
	wire _mesh_6_20_io_out_last_0;
	wire _mesh_6_20_io_out_valid_0;
	wire [31:0] _mesh_6_19_io_out_a_0;
	wire [31:0] _mesh_6_19_io_out_c_0;
	wire [31:0] _mesh_6_19_io_out_b_0;
	wire _mesh_6_19_io_out_control_0_dataflow;
	wire _mesh_6_19_io_out_control_0_propagate;
	wire [4:0] _mesh_6_19_io_out_control_0_shift;
	wire [2:0] _mesh_6_19_io_out_id_0;
	wire _mesh_6_19_io_out_last_0;
	wire _mesh_6_19_io_out_valid_0;
	wire [31:0] _mesh_6_18_io_out_a_0;
	wire [31:0] _mesh_6_18_io_out_c_0;
	wire [31:0] _mesh_6_18_io_out_b_0;
	wire _mesh_6_18_io_out_control_0_dataflow;
	wire _mesh_6_18_io_out_control_0_propagate;
	wire [4:0] _mesh_6_18_io_out_control_0_shift;
	wire [2:0] _mesh_6_18_io_out_id_0;
	wire _mesh_6_18_io_out_last_0;
	wire _mesh_6_18_io_out_valid_0;
	wire [31:0] _mesh_6_17_io_out_a_0;
	wire [31:0] _mesh_6_17_io_out_c_0;
	wire [31:0] _mesh_6_17_io_out_b_0;
	wire _mesh_6_17_io_out_control_0_dataflow;
	wire _mesh_6_17_io_out_control_0_propagate;
	wire [4:0] _mesh_6_17_io_out_control_0_shift;
	wire [2:0] _mesh_6_17_io_out_id_0;
	wire _mesh_6_17_io_out_last_0;
	wire _mesh_6_17_io_out_valid_0;
	wire [31:0] _mesh_6_16_io_out_a_0;
	wire [31:0] _mesh_6_16_io_out_c_0;
	wire [31:0] _mesh_6_16_io_out_b_0;
	wire _mesh_6_16_io_out_control_0_dataflow;
	wire _mesh_6_16_io_out_control_0_propagate;
	wire [4:0] _mesh_6_16_io_out_control_0_shift;
	wire [2:0] _mesh_6_16_io_out_id_0;
	wire _mesh_6_16_io_out_last_0;
	wire _mesh_6_16_io_out_valid_0;
	wire [31:0] _mesh_6_15_io_out_a_0;
	wire [31:0] _mesh_6_15_io_out_c_0;
	wire [31:0] _mesh_6_15_io_out_b_0;
	wire _mesh_6_15_io_out_control_0_dataflow;
	wire _mesh_6_15_io_out_control_0_propagate;
	wire [4:0] _mesh_6_15_io_out_control_0_shift;
	wire [2:0] _mesh_6_15_io_out_id_0;
	wire _mesh_6_15_io_out_last_0;
	wire _mesh_6_15_io_out_valid_0;
	wire [31:0] _mesh_6_14_io_out_a_0;
	wire [31:0] _mesh_6_14_io_out_c_0;
	wire [31:0] _mesh_6_14_io_out_b_0;
	wire _mesh_6_14_io_out_control_0_dataflow;
	wire _mesh_6_14_io_out_control_0_propagate;
	wire [4:0] _mesh_6_14_io_out_control_0_shift;
	wire [2:0] _mesh_6_14_io_out_id_0;
	wire _mesh_6_14_io_out_last_0;
	wire _mesh_6_14_io_out_valid_0;
	wire [31:0] _mesh_6_13_io_out_a_0;
	wire [31:0] _mesh_6_13_io_out_c_0;
	wire [31:0] _mesh_6_13_io_out_b_0;
	wire _mesh_6_13_io_out_control_0_dataflow;
	wire _mesh_6_13_io_out_control_0_propagate;
	wire [4:0] _mesh_6_13_io_out_control_0_shift;
	wire [2:0] _mesh_6_13_io_out_id_0;
	wire _mesh_6_13_io_out_last_0;
	wire _mesh_6_13_io_out_valid_0;
	wire [31:0] _mesh_6_12_io_out_a_0;
	wire [31:0] _mesh_6_12_io_out_c_0;
	wire [31:0] _mesh_6_12_io_out_b_0;
	wire _mesh_6_12_io_out_control_0_dataflow;
	wire _mesh_6_12_io_out_control_0_propagate;
	wire [4:0] _mesh_6_12_io_out_control_0_shift;
	wire [2:0] _mesh_6_12_io_out_id_0;
	wire _mesh_6_12_io_out_last_0;
	wire _mesh_6_12_io_out_valid_0;
	wire [31:0] _mesh_6_11_io_out_a_0;
	wire [31:0] _mesh_6_11_io_out_c_0;
	wire [31:0] _mesh_6_11_io_out_b_0;
	wire _mesh_6_11_io_out_control_0_dataflow;
	wire _mesh_6_11_io_out_control_0_propagate;
	wire [4:0] _mesh_6_11_io_out_control_0_shift;
	wire [2:0] _mesh_6_11_io_out_id_0;
	wire _mesh_6_11_io_out_last_0;
	wire _mesh_6_11_io_out_valid_0;
	wire [31:0] _mesh_6_10_io_out_a_0;
	wire [31:0] _mesh_6_10_io_out_c_0;
	wire [31:0] _mesh_6_10_io_out_b_0;
	wire _mesh_6_10_io_out_control_0_dataflow;
	wire _mesh_6_10_io_out_control_0_propagate;
	wire [4:0] _mesh_6_10_io_out_control_0_shift;
	wire [2:0] _mesh_6_10_io_out_id_0;
	wire _mesh_6_10_io_out_last_0;
	wire _mesh_6_10_io_out_valid_0;
	wire [31:0] _mesh_6_9_io_out_a_0;
	wire [31:0] _mesh_6_9_io_out_c_0;
	wire [31:0] _mesh_6_9_io_out_b_0;
	wire _mesh_6_9_io_out_control_0_dataflow;
	wire _mesh_6_9_io_out_control_0_propagate;
	wire [4:0] _mesh_6_9_io_out_control_0_shift;
	wire [2:0] _mesh_6_9_io_out_id_0;
	wire _mesh_6_9_io_out_last_0;
	wire _mesh_6_9_io_out_valid_0;
	wire [31:0] _mesh_6_8_io_out_a_0;
	wire [31:0] _mesh_6_8_io_out_c_0;
	wire [31:0] _mesh_6_8_io_out_b_0;
	wire _mesh_6_8_io_out_control_0_dataflow;
	wire _mesh_6_8_io_out_control_0_propagate;
	wire [4:0] _mesh_6_8_io_out_control_0_shift;
	wire [2:0] _mesh_6_8_io_out_id_0;
	wire _mesh_6_8_io_out_last_0;
	wire _mesh_6_8_io_out_valid_0;
	wire [31:0] _mesh_6_7_io_out_a_0;
	wire [31:0] _mesh_6_7_io_out_c_0;
	wire [31:0] _mesh_6_7_io_out_b_0;
	wire _mesh_6_7_io_out_control_0_dataflow;
	wire _mesh_6_7_io_out_control_0_propagate;
	wire [4:0] _mesh_6_7_io_out_control_0_shift;
	wire [2:0] _mesh_6_7_io_out_id_0;
	wire _mesh_6_7_io_out_last_0;
	wire _mesh_6_7_io_out_valid_0;
	wire [31:0] _mesh_6_6_io_out_a_0;
	wire [31:0] _mesh_6_6_io_out_c_0;
	wire [31:0] _mesh_6_6_io_out_b_0;
	wire _mesh_6_6_io_out_control_0_dataflow;
	wire _mesh_6_6_io_out_control_0_propagate;
	wire [4:0] _mesh_6_6_io_out_control_0_shift;
	wire [2:0] _mesh_6_6_io_out_id_0;
	wire _mesh_6_6_io_out_last_0;
	wire _mesh_6_6_io_out_valid_0;
	wire [31:0] _mesh_6_5_io_out_a_0;
	wire [31:0] _mesh_6_5_io_out_c_0;
	wire [31:0] _mesh_6_5_io_out_b_0;
	wire _mesh_6_5_io_out_control_0_dataflow;
	wire _mesh_6_5_io_out_control_0_propagate;
	wire [4:0] _mesh_6_5_io_out_control_0_shift;
	wire [2:0] _mesh_6_5_io_out_id_0;
	wire _mesh_6_5_io_out_last_0;
	wire _mesh_6_5_io_out_valid_0;
	wire [31:0] _mesh_6_4_io_out_a_0;
	wire [31:0] _mesh_6_4_io_out_c_0;
	wire [31:0] _mesh_6_4_io_out_b_0;
	wire _mesh_6_4_io_out_control_0_dataflow;
	wire _mesh_6_4_io_out_control_0_propagate;
	wire [4:0] _mesh_6_4_io_out_control_0_shift;
	wire [2:0] _mesh_6_4_io_out_id_0;
	wire _mesh_6_4_io_out_last_0;
	wire _mesh_6_4_io_out_valid_0;
	wire [31:0] _mesh_6_3_io_out_a_0;
	wire [31:0] _mesh_6_3_io_out_c_0;
	wire [31:0] _mesh_6_3_io_out_b_0;
	wire _mesh_6_3_io_out_control_0_dataflow;
	wire _mesh_6_3_io_out_control_0_propagate;
	wire [4:0] _mesh_6_3_io_out_control_0_shift;
	wire [2:0] _mesh_6_3_io_out_id_0;
	wire _mesh_6_3_io_out_last_0;
	wire _mesh_6_3_io_out_valid_0;
	wire [31:0] _mesh_6_2_io_out_a_0;
	wire [31:0] _mesh_6_2_io_out_c_0;
	wire [31:0] _mesh_6_2_io_out_b_0;
	wire _mesh_6_2_io_out_control_0_dataflow;
	wire _mesh_6_2_io_out_control_0_propagate;
	wire [4:0] _mesh_6_2_io_out_control_0_shift;
	wire [2:0] _mesh_6_2_io_out_id_0;
	wire _mesh_6_2_io_out_last_0;
	wire _mesh_6_2_io_out_valid_0;
	wire [31:0] _mesh_6_1_io_out_a_0;
	wire [31:0] _mesh_6_1_io_out_c_0;
	wire [31:0] _mesh_6_1_io_out_b_0;
	wire _mesh_6_1_io_out_control_0_dataflow;
	wire _mesh_6_1_io_out_control_0_propagate;
	wire [4:0] _mesh_6_1_io_out_control_0_shift;
	wire [2:0] _mesh_6_1_io_out_id_0;
	wire _mesh_6_1_io_out_last_0;
	wire _mesh_6_1_io_out_valid_0;
	wire [31:0] _mesh_6_0_io_out_a_0;
	wire [31:0] _mesh_6_0_io_out_c_0;
	wire [31:0] _mesh_6_0_io_out_b_0;
	wire _mesh_6_0_io_out_control_0_dataflow;
	wire _mesh_6_0_io_out_control_0_propagate;
	wire [4:0] _mesh_6_0_io_out_control_0_shift;
	wire [2:0] _mesh_6_0_io_out_id_0;
	wire _mesh_6_0_io_out_last_0;
	wire _mesh_6_0_io_out_valid_0;
	wire [31:0] _mesh_5_31_io_out_a_0;
	wire [31:0] _mesh_5_31_io_out_c_0;
	wire [31:0] _mesh_5_31_io_out_b_0;
	wire _mesh_5_31_io_out_control_0_dataflow;
	wire _mesh_5_31_io_out_control_0_propagate;
	wire [4:0] _mesh_5_31_io_out_control_0_shift;
	wire [2:0] _mesh_5_31_io_out_id_0;
	wire _mesh_5_31_io_out_last_0;
	wire _mesh_5_31_io_out_valid_0;
	wire [31:0] _mesh_5_30_io_out_a_0;
	wire [31:0] _mesh_5_30_io_out_c_0;
	wire [31:0] _mesh_5_30_io_out_b_0;
	wire _mesh_5_30_io_out_control_0_dataflow;
	wire _mesh_5_30_io_out_control_0_propagate;
	wire [4:0] _mesh_5_30_io_out_control_0_shift;
	wire [2:0] _mesh_5_30_io_out_id_0;
	wire _mesh_5_30_io_out_last_0;
	wire _mesh_5_30_io_out_valid_0;
	wire [31:0] _mesh_5_29_io_out_a_0;
	wire [31:0] _mesh_5_29_io_out_c_0;
	wire [31:0] _mesh_5_29_io_out_b_0;
	wire _mesh_5_29_io_out_control_0_dataflow;
	wire _mesh_5_29_io_out_control_0_propagate;
	wire [4:0] _mesh_5_29_io_out_control_0_shift;
	wire [2:0] _mesh_5_29_io_out_id_0;
	wire _mesh_5_29_io_out_last_0;
	wire _mesh_5_29_io_out_valid_0;
	wire [31:0] _mesh_5_28_io_out_a_0;
	wire [31:0] _mesh_5_28_io_out_c_0;
	wire [31:0] _mesh_5_28_io_out_b_0;
	wire _mesh_5_28_io_out_control_0_dataflow;
	wire _mesh_5_28_io_out_control_0_propagate;
	wire [4:0] _mesh_5_28_io_out_control_0_shift;
	wire [2:0] _mesh_5_28_io_out_id_0;
	wire _mesh_5_28_io_out_last_0;
	wire _mesh_5_28_io_out_valid_0;
	wire [31:0] _mesh_5_27_io_out_a_0;
	wire [31:0] _mesh_5_27_io_out_c_0;
	wire [31:0] _mesh_5_27_io_out_b_0;
	wire _mesh_5_27_io_out_control_0_dataflow;
	wire _mesh_5_27_io_out_control_0_propagate;
	wire [4:0] _mesh_5_27_io_out_control_0_shift;
	wire [2:0] _mesh_5_27_io_out_id_0;
	wire _mesh_5_27_io_out_last_0;
	wire _mesh_5_27_io_out_valid_0;
	wire [31:0] _mesh_5_26_io_out_a_0;
	wire [31:0] _mesh_5_26_io_out_c_0;
	wire [31:0] _mesh_5_26_io_out_b_0;
	wire _mesh_5_26_io_out_control_0_dataflow;
	wire _mesh_5_26_io_out_control_0_propagate;
	wire [4:0] _mesh_5_26_io_out_control_0_shift;
	wire [2:0] _mesh_5_26_io_out_id_0;
	wire _mesh_5_26_io_out_last_0;
	wire _mesh_5_26_io_out_valid_0;
	wire [31:0] _mesh_5_25_io_out_a_0;
	wire [31:0] _mesh_5_25_io_out_c_0;
	wire [31:0] _mesh_5_25_io_out_b_0;
	wire _mesh_5_25_io_out_control_0_dataflow;
	wire _mesh_5_25_io_out_control_0_propagate;
	wire [4:0] _mesh_5_25_io_out_control_0_shift;
	wire [2:0] _mesh_5_25_io_out_id_0;
	wire _mesh_5_25_io_out_last_0;
	wire _mesh_5_25_io_out_valid_0;
	wire [31:0] _mesh_5_24_io_out_a_0;
	wire [31:0] _mesh_5_24_io_out_c_0;
	wire [31:0] _mesh_5_24_io_out_b_0;
	wire _mesh_5_24_io_out_control_0_dataflow;
	wire _mesh_5_24_io_out_control_0_propagate;
	wire [4:0] _mesh_5_24_io_out_control_0_shift;
	wire [2:0] _mesh_5_24_io_out_id_0;
	wire _mesh_5_24_io_out_last_0;
	wire _mesh_5_24_io_out_valid_0;
	wire [31:0] _mesh_5_23_io_out_a_0;
	wire [31:0] _mesh_5_23_io_out_c_0;
	wire [31:0] _mesh_5_23_io_out_b_0;
	wire _mesh_5_23_io_out_control_0_dataflow;
	wire _mesh_5_23_io_out_control_0_propagate;
	wire [4:0] _mesh_5_23_io_out_control_0_shift;
	wire [2:0] _mesh_5_23_io_out_id_0;
	wire _mesh_5_23_io_out_last_0;
	wire _mesh_5_23_io_out_valid_0;
	wire [31:0] _mesh_5_22_io_out_a_0;
	wire [31:0] _mesh_5_22_io_out_c_0;
	wire [31:0] _mesh_5_22_io_out_b_0;
	wire _mesh_5_22_io_out_control_0_dataflow;
	wire _mesh_5_22_io_out_control_0_propagate;
	wire [4:0] _mesh_5_22_io_out_control_0_shift;
	wire [2:0] _mesh_5_22_io_out_id_0;
	wire _mesh_5_22_io_out_last_0;
	wire _mesh_5_22_io_out_valid_0;
	wire [31:0] _mesh_5_21_io_out_a_0;
	wire [31:0] _mesh_5_21_io_out_c_0;
	wire [31:0] _mesh_5_21_io_out_b_0;
	wire _mesh_5_21_io_out_control_0_dataflow;
	wire _mesh_5_21_io_out_control_0_propagate;
	wire [4:0] _mesh_5_21_io_out_control_0_shift;
	wire [2:0] _mesh_5_21_io_out_id_0;
	wire _mesh_5_21_io_out_last_0;
	wire _mesh_5_21_io_out_valid_0;
	wire [31:0] _mesh_5_20_io_out_a_0;
	wire [31:0] _mesh_5_20_io_out_c_0;
	wire [31:0] _mesh_5_20_io_out_b_0;
	wire _mesh_5_20_io_out_control_0_dataflow;
	wire _mesh_5_20_io_out_control_0_propagate;
	wire [4:0] _mesh_5_20_io_out_control_0_shift;
	wire [2:0] _mesh_5_20_io_out_id_0;
	wire _mesh_5_20_io_out_last_0;
	wire _mesh_5_20_io_out_valid_0;
	wire [31:0] _mesh_5_19_io_out_a_0;
	wire [31:0] _mesh_5_19_io_out_c_0;
	wire [31:0] _mesh_5_19_io_out_b_0;
	wire _mesh_5_19_io_out_control_0_dataflow;
	wire _mesh_5_19_io_out_control_0_propagate;
	wire [4:0] _mesh_5_19_io_out_control_0_shift;
	wire [2:0] _mesh_5_19_io_out_id_0;
	wire _mesh_5_19_io_out_last_0;
	wire _mesh_5_19_io_out_valid_0;
	wire [31:0] _mesh_5_18_io_out_a_0;
	wire [31:0] _mesh_5_18_io_out_c_0;
	wire [31:0] _mesh_5_18_io_out_b_0;
	wire _mesh_5_18_io_out_control_0_dataflow;
	wire _mesh_5_18_io_out_control_0_propagate;
	wire [4:0] _mesh_5_18_io_out_control_0_shift;
	wire [2:0] _mesh_5_18_io_out_id_0;
	wire _mesh_5_18_io_out_last_0;
	wire _mesh_5_18_io_out_valid_0;
	wire [31:0] _mesh_5_17_io_out_a_0;
	wire [31:0] _mesh_5_17_io_out_c_0;
	wire [31:0] _mesh_5_17_io_out_b_0;
	wire _mesh_5_17_io_out_control_0_dataflow;
	wire _mesh_5_17_io_out_control_0_propagate;
	wire [4:0] _mesh_5_17_io_out_control_0_shift;
	wire [2:0] _mesh_5_17_io_out_id_0;
	wire _mesh_5_17_io_out_last_0;
	wire _mesh_5_17_io_out_valid_0;
	wire [31:0] _mesh_5_16_io_out_a_0;
	wire [31:0] _mesh_5_16_io_out_c_0;
	wire [31:0] _mesh_5_16_io_out_b_0;
	wire _mesh_5_16_io_out_control_0_dataflow;
	wire _mesh_5_16_io_out_control_0_propagate;
	wire [4:0] _mesh_5_16_io_out_control_0_shift;
	wire [2:0] _mesh_5_16_io_out_id_0;
	wire _mesh_5_16_io_out_last_0;
	wire _mesh_5_16_io_out_valid_0;
	wire [31:0] _mesh_5_15_io_out_a_0;
	wire [31:0] _mesh_5_15_io_out_c_0;
	wire [31:0] _mesh_5_15_io_out_b_0;
	wire _mesh_5_15_io_out_control_0_dataflow;
	wire _mesh_5_15_io_out_control_0_propagate;
	wire [4:0] _mesh_5_15_io_out_control_0_shift;
	wire [2:0] _mesh_5_15_io_out_id_0;
	wire _mesh_5_15_io_out_last_0;
	wire _mesh_5_15_io_out_valid_0;
	wire [31:0] _mesh_5_14_io_out_a_0;
	wire [31:0] _mesh_5_14_io_out_c_0;
	wire [31:0] _mesh_5_14_io_out_b_0;
	wire _mesh_5_14_io_out_control_0_dataflow;
	wire _mesh_5_14_io_out_control_0_propagate;
	wire [4:0] _mesh_5_14_io_out_control_0_shift;
	wire [2:0] _mesh_5_14_io_out_id_0;
	wire _mesh_5_14_io_out_last_0;
	wire _mesh_5_14_io_out_valid_0;
	wire [31:0] _mesh_5_13_io_out_a_0;
	wire [31:0] _mesh_5_13_io_out_c_0;
	wire [31:0] _mesh_5_13_io_out_b_0;
	wire _mesh_5_13_io_out_control_0_dataflow;
	wire _mesh_5_13_io_out_control_0_propagate;
	wire [4:0] _mesh_5_13_io_out_control_0_shift;
	wire [2:0] _mesh_5_13_io_out_id_0;
	wire _mesh_5_13_io_out_last_0;
	wire _mesh_5_13_io_out_valid_0;
	wire [31:0] _mesh_5_12_io_out_a_0;
	wire [31:0] _mesh_5_12_io_out_c_0;
	wire [31:0] _mesh_5_12_io_out_b_0;
	wire _mesh_5_12_io_out_control_0_dataflow;
	wire _mesh_5_12_io_out_control_0_propagate;
	wire [4:0] _mesh_5_12_io_out_control_0_shift;
	wire [2:0] _mesh_5_12_io_out_id_0;
	wire _mesh_5_12_io_out_last_0;
	wire _mesh_5_12_io_out_valid_0;
	wire [31:0] _mesh_5_11_io_out_a_0;
	wire [31:0] _mesh_5_11_io_out_c_0;
	wire [31:0] _mesh_5_11_io_out_b_0;
	wire _mesh_5_11_io_out_control_0_dataflow;
	wire _mesh_5_11_io_out_control_0_propagate;
	wire [4:0] _mesh_5_11_io_out_control_0_shift;
	wire [2:0] _mesh_5_11_io_out_id_0;
	wire _mesh_5_11_io_out_last_0;
	wire _mesh_5_11_io_out_valid_0;
	wire [31:0] _mesh_5_10_io_out_a_0;
	wire [31:0] _mesh_5_10_io_out_c_0;
	wire [31:0] _mesh_5_10_io_out_b_0;
	wire _mesh_5_10_io_out_control_0_dataflow;
	wire _mesh_5_10_io_out_control_0_propagate;
	wire [4:0] _mesh_5_10_io_out_control_0_shift;
	wire [2:0] _mesh_5_10_io_out_id_0;
	wire _mesh_5_10_io_out_last_0;
	wire _mesh_5_10_io_out_valid_0;
	wire [31:0] _mesh_5_9_io_out_a_0;
	wire [31:0] _mesh_5_9_io_out_c_0;
	wire [31:0] _mesh_5_9_io_out_b_0;
	wire _mesh_5_9_io_out_control_0_dataflow;
	wire _mesh_5_9_io_out_control_0_propagate;
	wire [4:0] _mesh_5_9_io_out_control_0_shift;
	wire [2:0] _mesh_5_9_io_out_id_0;
	wire _mesh_5_9_io_out_last_0;
	wire _mesh_5_9_io_out_valid_0;
	wire [31:0] _mesh_5_8_io_out_a_0;
	wire [31:0] _mesh_5_8_io_out_c_0;
	wire [31:0] _mesh_5_8_io_out_b_0;
	wire _mesh_5_8_io_out_control_0_dataflow;
	wire _mesh_5_8_io_out_control_0_propagate;
	wire [4:0] _mesh_5_8_io_out_control_0_shift;
	wire [2:0] _mesh_5_8_io_out_id_0;
	wire _mesh_5_8_io_out_last_0;
	wire _mesh_5_8_io_out_valid_0;
	wire [31:0] _mesh_5_7_io_out_a_0;
	wire [31:0] _mesh_5_7_io_out_c_0;
	wire [31:0] _mesh_5_7_io_out_b_0;
	wire _mesh_5_7_io_out_control_0_dataflow;
	wire _mesh_5_7_io_out_control_0_propagate;
	wire [4:0] _mesh_5_7_io_out_control_0_shift;
	wire [2:0] _mesh_5_7_io_out_id_0;
	wire _mesh_5_7_io_out_last_0;
	wire _mesh_5_7_io_out_valid_0;
	wire [31:0] _mesh_5_6_io_out_a_0;
	wire [31:0] _mesh_5_6_io_out_c_0;
	wire [31:0] _mesh_5_6_io_out_b_0;
	wire _mesh_5_6_io_out_control_0_dataflow;
	wire _mesh_5_6_io_out_control_0_propagate;
	wire [4:0] _mesh_5_6_io_out_control_0_shift;
	wire [2:0] _mesh_5_6_io_out_id_0;
	wire _mesh_5_6_io_out_last_0;
	wire _mesh_5_6_io_out_valid_0;
	wire [31:0] _mesh_5_5_io_out_a_0;
	wire [31:0] _mesh_5_5_io_out_c_0;
	wire [31:0] _mesh_5_5_io_out_b_0;
	wire _mesh_5_5_io_out_control_0_dataflow;
	wire _mesh_5_5_io_out_control_0_propagate;
	wire [4:0] _mesh_5_5_io_out_control_0_shift;
	wire [2:0] _mesh_5_5_io_out_id_0;
	wire _mesh_5_5_io_out_last_0;
	wire _mesh_5_5_io_out_valid_0;
	wire [31:0] _mesh_5_4_io_out_a_0;
	wire [31:0] _mesh_5_4_io_out_c_0;
	wire [31:0] _mesh_5_4_io_out_b_0;
	wire _mesh_5_4_io_out_control_0_dataflow;
	wire _mesh_5_4_io_out_control_0_propagate;
	wire [4:0] _mesh_5_4_io_out_control_0_shift;
	wire [2:0] _mesh_5_4_io_out_id_0;
	wire _mesh_5_4_io_out_last_0;
	wire _mesh_5_4_io_out_valid_0;
	wire [31:0] _mesh_5_3_io_out_a_0;
	wire [31:0] _mesh_5_3_io_out_c_0;
	wire [31:0] _mesh_5_3_io_out_b_0;
	wire _mesh_5_3_io_out_control_0_dataflow;
	wire _mesh_5_3_io_out_control_0_propagate;
	wire [4:0] _mesh_5_3_io_out_control_0_shift;
	wire [2:0] _mesh_5_3_io_out_id_0;
	wire _mesh_5_3_io_out_last_0;
	wire _mesh_5_3_io_out_valid_0;
	wire [31:0] _mesh_5_2_io_out_a_0;
	wire [31:0] _mesh_5_2_io_out_c_0;
	wire [31:0] _mesh_5_2_io_out_b_0;
	wire _mesh_5_2_io_out_control_0_dataflow;
	wire _mesh_5_2_io_out_control_0_propagate;
	wire [4:0] _mesh_5_2_io_out_control_0_shift;
	wire [2:0] _mesh_5_2_io_out_id_0;
	wire _mesh_5_2_io_out_last_0;
	wire _mesh_5_2_io_out_valid_0;
	wire [31:0] _mesh_5_1_io_out_a_0;
	wire [31:0] _mesh_5_1_io_out_c_0;
	wire [31:0] _mesh_5_1_io_out_b_0;
	wire _mesh_5_1_io_out_control_0_dataflow;
	wire _mesh_5_1_io_out_control_0_propagate;
	wire [4:0] _mesh_5_1_io_out_control_0_shift;
	wire [2:0] _mesh_5_1_io_out_id_0;
	wire _mesh_5_1_io_out_last_0;
	wire _mesh_5_1_io_out_valid_0;
	wire [31:0] _mesh_5_0_io_out_a_0;
	wire [31:0] _mesh_5_0_io_out_c_0;
	wire [31:0] _mesh_5_0_io_out_b_0;
	wire _mesh_5_0_io_out_control_0_dataflow;
	wire _mesh_5_0_io_out_control_0_propagate;
	wire [4:0] _mesh_5_0_io_out_control_0_shift;
	wire [2:0] _mesh_5_0_io_out_id_0;
	wire _mesh_5_0_io_out_last_0;
	wire _mesh_5_0_io_out_valid_0;
	wire [31:0] _mesh_4_31_io_out_a_0;
	wire [31:0] _mesh_4_31_io_out_c_0;
	wire [31:0] _mesh_4_31_io_out_b_0;
	wire _mesh_4_31_io_out_control_0_dataflow;
	wire _mesh_4_31_io_out_control_0_propagate;
	wire [4:0] _mesh_4_31_io_out_control_0_shift;
	wire [2:0] _mesh_4_31_io_out_id_0;
	wire _mesh_4_31_io_out_last_0;
	wire _mesh_4_31_io_out_valid_0;
	wire [31:0] _mesh_4_30_io_out_a_0;
	wire [31:0] _mesh_4_30_io_out_c_0;
	wire [31:0] _mesh_4_30_io_out_b_0;
	wire _mesh_4_30_io_out_control_0_dataflow;
	wire _mesh_4_30_io_out_control_0_propagate;
	wire [4:0] _mesh_4_30_io_out_control_0_shift;
	wire [2:0] _mesh_4_30_io_out_id_0;
	wire _mesh_4_30_io_out_last_0;
	wire _mesh_4_30_io_out_valid_0;
	wire [31:0] _mesh_4_29_io_out_a_0;
	wire [31:0] _mesh_4_29_io_out_c_0;
	wire [31:0] _mesh_4_29_io_out_b_0;
	wire _mesh_4_29_io_out_control_0_dataflow;
	wire _mesh_4_29_io_out_control_0_propagate;
	wire [4:0] _mesh_4_29_io_out_control_0_shift;
	wire [2:0] _mesh_4_29_io_out_id_0;
	wire _mesh_4_29_io_out_last_0;
	wire _mesh_4_29_io_out_valid_0;
	wire [31:0] _mesh_4_28_io_out_a_0;
	wire [31:0] _mesh_4_28_io_out_c_0;
	wire [31:0] _mesh_4_28_io_out_b_0;
	wire _mesh_4_28_io_out_control_0_dataflow;
	wire _mesh_4_28_io_out_control_0_propagate;
	wire [4:0] _mesh_4_28_io_out_control_0_shift;
	wire [2:0] _mesh_4_28_io_out_id_0;
	wire _mesh_4_28_io_out_last_0;
	wire _mesh_4_28_io_out_valid_0;
	wire [31:0] _mesh_4_27_io_out_a_0;
	wire [31:0] _mesh_4_27_io_out_c_0;
	wire [31:0] _mesh_4_27_io_out_b_0;
	wire _mesh_4_27_io_out_control_0_dataflow;
	wire _mesh_4_27_io_out_control_0_propagate;
	wire [4:0] _mesh_4_27_io_out_control_0_shift;
	wire [2:0] _mesh_4_27_io_out_id_0;
	wire _mesh_4_27_io_out_last_0;
	wire _mesh_4_27_io_out_valid_0;
	wire [31:0] _mesh_4_26_io_out_a_0;
	wire [31:0] _mesh_4_26_io_out_c_0;
	wire [31:0] _mesh_4_26_io_out_b_0;
	wire _mesh_4_26_io_out_control_0_dataflow;
	wire _mesh_4_26_io_out_control_0_propagate;
	wire [4:0] _mesh_4_26_io_out_control_0_shift;
	wire [2:0] _mesh_4_26_io_out_id_0;
	wire _mesh_4_26_io_out_last_0;
	wire _mesh_4_26_io_out_valid_0;
	wire [31:0] _mesh_4_25_io_out_a_0;
	wire [31:0] _mesh_4_25_io_out_c_0;
	wire [31:0] _mesh_4_25_io_out_b_0;
	wire _mesh_4_25_io_out_control_0_dataflow;
	wire _mesh_4_25_io_out_control_0_propagate;
	wire [4:0] _mesh_4_25_io_out_control_0_shift;
	wire [2:0] _mesh_4_25_io_out_id_0;
	wire _mesh_4_25_io_out_last_0;
	wire _mesh_4_25_io_out_valid_0;
	wire [31:0] _mesh_4_24_io_out_a_0;
	wire [31:0] _mesh_4_24_io_out_c_0;
	wire [31:0] _mesh_4_24_io_out_b_0;
	wire _mesh_4_24_io_out_control_0_dataflow;
	wire _mesh_4_24_io_out_control_0_propagate;
	wire [4:0] _mesh_4_24_io_out_control_0_shift;
	wire [2:0] _mesh_4_24_io_out_id_0;
	wire _mesh_4_24_io_out_last_0;
	wire _mesh_4_24_io_out_valid_0;
	wire [31:0] _mesh_4_23_io_out_a_0;
	wire [31:0] _mesh_4_23_io_out_c_0;
	wire [31:0] _mesh_4_23_io_out_b_0;
	wire _mesh_4_23_io_out_control_0_dataflow;
	wire _mesh_4_23_io_out_control_0_propagate;
	wire [4:0] _mesh_4_23_io_out_control_0_shift;
	wire [2:0] _mesh_4_23_io_out_id_0;
	wire _mesh_4_23_io_out_last_0;
	wire _mesh_4_23_io_out_valid_0;
	wire [31:0] _mesh_4_22_io_out_a_0;
	wire [31:0] _mesh_4_22_io_out_c_0;
	wire [31:0] _mesh_4_22_io_out_b_0;
	wire _mesh_4_22_io_out_control_0_dataflow;
	wire _mesh_4_22_io_out_control_0_propagate;
	wire [4:0] _mesh_4_22_io_out_control_0_shift;
	wire [2:0] _mesh_4_22_io_out_id_0;
	wire _mesh_4_22_io_out_last_0;
	wire _mesh_4_22_io_out_valid_0;
	wire [31:0] _mesh_4_21_io_out_a_0;
	wire [31:0] _mesh_4_21_io_out_c_0;
	wire [31:0] _mesh_4_21_io_out_b_0;
	wire _mesh_4_21_io_out_control_0_dataflow;
	wire _mesh_4_21_io_out_control_0_propagate;
	wire [4:0] _mesh_4_21_io_out_control_0_shift;
	wire [2:0] _mesh_4_21_io_out_id_0;
	wire _mesh_4_21_io_out_last_0;
	wire _mesh_4_21_io_out_valid_0;
	wire [31:0] _mesh_4_20_io_out_a_0;
	wire [31:0] _mesh_4_20_io_out_c_0;
	wire [31:0] _mesh_4_20_io_out_b_0;
	wire _mesh_4_20_io_out_control_0_dataflow;
	wire _mesh_4_20_io_out_control_0_propagate;
	wire [4:0] _mesh_4_20_io_out_control_0_shift;
	wire [2:0] _mesh_4_20_io_out_id_0;
	wire _mesh_4_20_io_out_last_0;
	wire _mesh_4_20_io_out_valid_0;
	wire [31:0] _mesh_4_19_io_out_a_0;
	wire [31:0] _mesh_4_19_io_out_c_0;
	wire [31:0] _mesh_4_19_io_out_b_0;
	wire _mesh_4_19_io_out_control_0_dataflow;
	wire _mesh_4_19_io_out_control_0_propagate;
	wire [4:0] _mesh_4_19_io_out_control_0_shift;
	wire [2:0] _mesh_4_19_io_out_id_0;
	wire _mesh_4_19_io_out_last_0;
	wire _mesh_4_19_io_out_valid_0;
	wire [31:0] _mesh_4_18_io_out_a_0;
	wire [31:0] _mesh_4_18_io_out_c_0;
	wire [31:0] _mesh_4_18_io_out_b_0;
	wire _mesh_4_18_io_out_control_0_dataflow;
	wire _mesh_4_18_io_out_control_0_propagate;
	wire [4:0] _mesh_4_18_io_out_control_0_shift;
	wire [2:0] _mesh_4_18_io_out_id_0;
	wire _mesh_4_18_io_out_last_0;
	wire _mesh_4_18_io_out_valid_0;
	wire [31:0] _mesh_4_17_io_out_a_0;
	wire [31:0] _mesh_4_17_io_out_c_0;
	wire [31:0] _mesh_4_17_io_out_b_0;
	wire _mesh_4_17_io_out_control_0_dataflow;
	wire _mesh_4_17_io_out_control_0_propagate;
	wire [4:0] _mesh_4_17_io_out_control_0_shift;
	wire [2:0] _mesh_4_17_io_out_id_0;
	wire _mesh_4_17_io_out_last_0;
	wire _mesh_4_17_io_out_valid_0;
	wire [31:0] _mesh_4_16_io_out_a_0;
	wire [31:0] _mesh_4_16_io_out_c_0;
	wire [31:0] _mesh_4_16_io_out_b_0;
	wire _mesh_4_16_io_out_control_0_dataflow;
	wire _mesh_4_16_io_out_control_0_propagate;
	wire [4:0] _mesh_4_16_io_out_control_0_shift;
	wire [2:0] _mesh_4_16_io_out_id_0;
	wire _mesh_4_16_io_out_last_0;
	wire _mesh_4_16_io_out_valid_0;
	wire [31:0] _mesh_4_15_io_out_a_0;
	wire [31:0] _mesh_4_15_io_out_c_0;
	wire [31:0] _mesh_4_15_io_out_b_0;
	wire _mesh_4_15_io_out_control_0_dataflow;
	wire _mesh_4_15_io_out_control_0_propagate;
	wire [4:0] _mesh_4_15_io_out_control_0_shift;
	wire [2:0] _mesh_4_15_io_out_id_0;
	wire _mesh_4_15_io_out_last_0;
	wire _mesh_4_15_io_out_valid_0;
	wire [31:0] _mesh_4_14_io_out_a_0;
	wire [31:0] _mesh_4_14_io_out_c_0;
	wire [31:0] _mesh_4_14_io_out_b_0;
	wire _mesh_4_14_io_out_control_0_dataflow;
	wire _mesh_4_14_io_out_control_0_propagate;
	wire [4:0] _mesh_4_14_io_out_control_0_shift;
	wire [2:0] _mesh_4_14_io_out_id_0;
	wire _mesh_4_14_io_out_last_0;
	wire _mesh_4_14_io_out_valid_0;
	wire [31:0] _mesh_4_13_io_out_a_0;
	wire [31:0] _mesh_4_13_io_out_c_0;
	wire [31:0] _mesh_4_13_io_out_b_0;
	wire _mesh_4_13_io_out_control_0_dataflow;
	wire _mesh_4_13_io_out_control_0_propagate;
	wire [4:0] _mesh_4_13_io_out_control_0_shift;
	wire [2:0] _mesh_4_13_io_out_id_0;
	wire _mesh_4_13_io_out_last_0;
	wire _mesh_4_13_io_out_valid_0;
	wire [31:0] _mesh_4_12_io_out_a_0;
	wire [31:0] _mesh_4_12_io_out_c_0;
	wire [31:0] _mesh_4_12_io_out_b_0;
	wire _mesh_4_12_io_out_control_0_dataflow;
	wire _mesh_4_12_io_out_control_0_propagate;
	wire [4:0] _mesh_4_12_io_out_control_0_shift;
	wire [2:0] _mesh_4_12_io_out_id_0;
	wire _mesh_4_12_io_out_last_0;
	wire _mesh_4_12_io_out_valid_0;
	wire [31:0] _mesh_4_11_io_out_a_0;
	wire [31:0] _mesh_4_11_io_out_c_0;
	wire [31:0] _mesh_4_11_io_out_b_0;
	wire _mesh_4_11_io_out_control_0_dataflow;
	wire _mesh_4_11_io_out_control_0_propagate;
	wire [4:0] _mesh_4_11_io_out_control_0_shift;
	wire [2:0] _mesh_4_11_io_out_id_0;
	wire _mesh_4_11_io_out_last_0;
	wire _mesh_4_11_io_out_valid_0;
	wire [31:0] _mesh_4_10_io_out_a_0;
	wire [31:0] _mesh_4_10_io_out_c_0;
	wire [31:0] _mesh_4_10_io_out_b_0;
	wire _mesh_4_10_io_out_control_0_dataflow;
	wire _mesh_4_10_io_out_control_0_propagate;
	wire [4:0] _mesh_4_10_io_out_control_0_shift;
	wire [2:0] _mesh_4_10_io_out_id_0;
	wire _mesh_4_10_io_out_last_0;
	wire _mesh_4_10_io_out_valid_0;
	wire [31:0] _mesh_4_9_io_out_a_0;
	wire [31:0] _mesh_4_9_io_out_c_0;
	wire [31:0] _mesh_4_9_io_out_b_0;
	wire _mesh_4_9_io_out_control_0_dataflow;
	wire _mesh_4_9_io_out_control_0_propagate;
	wire [4:0] _mesh_4_9_io_out_control_0_shift;
	wire [2:0] _mesh_4_9_io_out_id_0;
	wire _mesh_4_9_io_out_last_0;
	wire _mesh_4_9_io_out_valid_0;
	wire [31:0] _mesh_4_8_io_out_a_0;
	wire [31:0] _mesh_4_8_io_out_c_0;
	wire [31:0] _mesh_4_8_io_out_b_0;
	wire _mesh_4_8_io_out_control_0_dataflow;
	wire _mesh_4_8_io_out_control_0_propagate;
	wire [4:0] _mesh_4_8_io_out_control_0_shift;
	wire [2:0] _mesh_4_8_io_out_id_0;
	wire _mesh_4_8_io_out_last_0;
	wire _mesh_4_8_io_out_valid_0;
	wire [31:0] _mesh_4_7_io_out_a_0;
	wire [31:0] _mesh_4_7_io_out_c_0;
	wire [31:0] _mesh_4_7_io_out_b_0;
	wire _mesh_4_7_io_out_control_0_dataflow;
	wire _mesh_4_7_io_out_control_0_propagate;
	wire [4:0] _mesh_4_7_io_out_control_0_shift;
	wire [2:0] _mesh_4_7_io_out_id_0;
	wire _mesh_4_7_io_out_last_0;
	wire _mesh_4_7_io_out_valid_0;
	wire [31:0] _mesh_4_6_io_out_a_0;
	wire [31:0] _mesh_4_6_io_out_c_0;
	wire [31:0] _mesh_4_6_io_out_b_0;
	wire _mesh_4_6_io_out_control_0_dataflow;
	wire _mesh_4_6_io_out_control_0_propagate;
	wire [4:0] _mesh_4_6_io_out_control_0_shift;
	wire [2:0] _mesh_4_6_io_out_id_0;
	wire _mesh_4_6_io_out_last_0;
	wire _mesh_4_6_io_out_valid_0;
	wire [31:0] _mesh_4_5_io_out_a_0;
	wire [31:0] _mesh_4_5_io_out_c_0;
	wire [31:0] _mesh_4_5_io_out_b_0;
	wire _mesh_4_5_io_out_control_0_dataflow;
	wire _mesh_4_5_io_out_control_0_propagate;
	wire [4:0] _mesh_4_5_io_out_control_0_shift;
	wire [2:0] _mesh_4_5_io_out_id_0;
	wire _mesh_4_5_io_out_last_0;
	wire _mesh_4_5_io_out_valid_0;
	wire [31:0] _mesh_4_4_io_out_a_0;
	wire [31:0] _mesh_4_4_io_out_c_0;
	wire [31:0] _mesh_4_4_io_out_b_0;
	wire _mesh_4_4_io_out_control_0_dataflow;
	wire _mesh_4_4_io_out_control_0_propagate;
	wire [4:0] _mesh_4_4_io_out_control_0_shift;
	wire [2:0] _mesh_4_4_io_out_id_0;
	wire _mesh_4_4_io_out_last_0;
	wire _mesh_4_4_io_out_valid_0;
	wire [31:0] _mesh_4_3_io_out_a_0;
	wire [31:0] _mesh_4_3_io_out_c_0;
	wire [31:0] _mesh_4_3_io_out_b_0;
	wire _mesh_4_3_io_out_control_0_dataflow;
	wire _mesh_4_3_io_out_control_0_propagate;
	wire [4:0] _mesh_4_3_io_out_control_0_shift;
	wire [2:0] _mesh_4_3_io_out_id_0;
	wire _mesh_4_3_io_out_last_0;
	wire _mesh_4_3_io_out_valid_0;
	wire [31:0] _mesh_4_2_io_out_a_0;
	wire [31:0] _mesh_4_2_io_out_c_0;
	wire [31:0] _mesh_4_2_io_out_b_0;
	wire _mesh_4_2_io_out_control_0_dataflow;
	wire _mesh_4_2_io_out_control_0_propagate;
	wire [4:0] _mesh_4_2_io_out_control_0_shift;
	wire [2:0] _mesh_4_2_io_out_id_0;
	wire _mesh_4_2_io_out_last_0;
	wire _mesh_4_2_io_out_valid_0;
	wire [31:0] _mesh_4_1_io_out_a_0;
	wire [31:0] _mesh_4_1_io_out_c_0;
	wire [31:0] _mesh_4_1_io_out_b_0;
	wire _mesh_4_1_io_out_control_0_dataflow;
	wire _mesh_4_1_io_out_control_0_propagate;
	wire [4:0] _mesh_4_1_io_out_control_0_shift;
	wire [2:0] _mesh_4_1_io_out_id_0;
	wire _mesh_4_1_io_out_last_0;
	wire _mesh_4_1_io_out_valid_0;
	wire [31:0] _mesh_4_0_io_out_a_0;
	wire [31:0] _mesh_4_0_io_out_c_0;
	wire [31:0] _mesh_4_0_io_out_b_0;
	wire _mesh_4_0_io_out_control_0_dataflow;
	wire _mesh_4_0_io_out_control_0_propagate;
	wire [4:0] _mesh_4_0_io_out_control_0_shift;
	wire [2:0] _mesh_4_0_io_out_id_0;
	wire _mesh_4_0_io_out_last_0;
	wire _mesh_4_0_io_out_valid_0;
	wire [31:0] _mesh_3_31_io_out_a_0;
	wire [31:0] _mesh_3_31_io_out_c_0;
	wire [31:0] _mesh_3_31_io_out_b_0;
	wire _mesh_3_31_io_out_control_0_dataflow;
	wire _mesh_3_31_io_out_control_0_propagate;
	wire [4:0] _mesh_3_31_io_out_control_0_shift;
	wire [2:0] _mesh_3_31_io_out_id_0;
	wire _mesh_3_31_io_out_last_0;
	wire _mesh_3_31_io_out_valid_0;
	wire [31:0] _mesh_3_30_io_out_a_0;
	wire [31:0] _mesh_3_30_io_out_c_0;
	wire [31:0] _mesh_3_30_io_out_b_0;
	wire _mesh_3_30_io_out_control_0_dataflow;
	wire _mesh_3_30_io_out_control_0_propagate;
	wire [4:0] _mesh_3_30_io_out_control_0_shift;
	wire [2:0] _mesh_3_30_io_out_id_0;
	wire _mesh_3_30_io_out_last_0;
	wire _mesh_3_30_io_out_valid_0;
	wire [31:0] _mesh_3_29_io_out_a_0;
	wire [31:0] _mesh_3_29_io_out_c_0;
	wire [31:0] _mesh_3_29_io_out_b_0;
	wire _mesh_3_29_io_out_control_0_dataflow;
	wire _mesh_3_29_io_out_control_0_propagate;
	wire [4:0] _mesh_3_29_io_out_control_0_shift;
	wire [2:0] _mesh_3_29_io_out_id_0;
	wire _mesh_3_29_io_out_last_0;
	wire _mesh_3_29_io_out_valid_0;
	wire [31:0] _mesh_3_28_io_out_a_0;
	wire [31:0] _mesh_3_28_io_out_c_0;
	wire [31:0] _mesh_3_28_io_out_b_0;
	wire _mesh_3_28_io_out_control_0_dataflow;
	wire _mesh_3_28_io_out_control_0_propagate;
	wire [4:0] _mesh_3_28_io_out_control_0_shift;
	wire [2:0] _mesh_3_28_io_out_id_0;
	wire _mesh_3_28_io_out_last_0;
	wire _mesh_3_28_io_out_valid_0;
	wire [31:0] _mesh_3_27_io_out_a_0;
	wire [31:0] _mesh_3_27_io_out_c_0;
	wire [31:0] _mesh_3_27_io_out_b_0;
	wire _mesh_3_27_io_out_control_0_dataflow;
	wire _mesh_3_27_io_out_control_0_propagate;
	wire [4:0] _mesh_3_27_io_out_control_0_shift;
	wire [2:0] _mesh_3_27_io_out_id_0;
	wire _mesh_3_27_io_out_last_0;
	wire _mesh_3_27_io_out_valid_0;
	wire [31:0] _mesh_3_26_io_out_a_0;
	wire [31:0] _mesh_3_26_io_out_c_0;
	wire [31:0] _mesh_3_26_io_out_b_0;
	wire _mesh_3_26_io_out_control_0_dataflow;
	wire _mesh_3_26_io_out_control_0_propagate;
	wire [4:0] _mesh_3_26_io_out_control_0_shift;
	wire [2:0] _mesh_3_26_io_out_id_0;
	wire _mesh_3_26_io_out_last_0;
	wire _mesh_3_26_io_out_valid_0;
	wire [31:0] _mesh_3_25_io_out_a_0;
	wire [31:0] _mesh_3_25_io_out_c_0;
	wire [31:0] _mesh_3_25_io_out_b_0;
	wire _mesh_3_25_io_out_control_0_dataflow;
	wire _mesh_3_25_io_out_control_0_propagate;
	wire [4:0] _mesh_3_25_io_out_control_0_shift;
	wire [2:0] _mesh_3_25_io_out_id_0;
	wire _mesh_3_25_io_out_last_0;
	wire _mesh_3_25_io_out_valid_0;
	wire [31:0] _mesh_3_24_io_out_a_0;
	wire [31:0] _mesh_3_24_io_out_c_0;
	wire [31:0] _mesh_3_24_io_out_b_0;
	wire _mesh_3_24_io_out_control_0_dataflow;
	wire _mesh_3_24_io_out_control_0_propagate;
	wire [4:0] _mesh_3_24_io_out_control_0_shift;
	wire [2:0] _mesh_3_24_io_out_id_0;
	wire _mesh_3_24_io_out_last_0;
	wire _mesh_3_24_io_out_valid_0;
	wire [31:0] _mesh_3_23_io_out_a_0;
	wire [31:0] _mesh_3_23_io_out_c_0;
	wire [31:0] _mesh_3_23_io_out_b_0;
	wire _mesh_3_23_io_out_control_0_dataflow;
	wire _mesh_3_23_io_out_control_0_propagate;
	wire [4:0] _mesh_3_23_io_out_control_0_shift;
	wire [2:0] _mesh_3_23_io_out_id_0;
	wire _mesh_3_23_io_out_last_0;
	wire _mesh_3_23_io_out_valid_0;
	wire [31:0] _mesh_3_22_io_out_a_0;
	wire [31:0] _mesh_3_22_io_out_c_0;
	wire [31:0] _mesh_3_22_io_out_b_0;
	wire _mesh_3_22_io_out_control_0_dataflow;
	wire _mesh_3_22_io_out_control_0_propagate;
	wire [4:0] _mesh_3_22_io_out_control_0_shift;
	wire [2:0] _mesh_3_22_io_out_id_0;
	wire _mesh_3_22_io_out_last_0;
	wire _mesh_3_22_io_out_valid_0;
	wire [31:0] _mesh_3_21_io_out_a_0;
	wire [31:0] _mesh_3_21_io_out_c_0;
	wire [31:0] _mesh_3_21_io_out_b_0;
	wire _mesh_3_21_io_out_control_0_dataflow;
	wire _mesh_3_21_io_out_control_0_propagate;
	wire [4:0] _mesh_3_21_io_out_control_0_shift;
	wire [2:0] _mesh_3_21_io_out_id_0;
	wire _mesh_3_21_io_out_last_0;
	wire _mesh_3_21_io_out_valid_0;
	wire [31:0] _mesh_3_20_io_out_a_0;
	wire [31:0] _mesh_3_20_io_out_c_0;
	wire [31:0] _mesh_3_20_io_out_b_0;
	wire _mesh_3_20_io_out_control_0_dataflow;
	wire _mesh_3_20_io_out_control_0_propagate;
	wire [4:0] _mesh_3_20_io_out_control_0_shift;
	wire [2:0] _mesh_3_20_io_out_id_0;
	wire _mesh_3_20_io_out_last_0;
	wire _mesh_3_20_io_out_valid_0;
	wire [31:0] _mesh_3_19_io_out_a_0;
	wire [31:0] _mesh_3_19_io_out_c_0;
	wire [31:0] _mesh_3_19_io_out_b_0;
	wire _mesh_3_19_io_out_control_0_dataflow;
	wire _mesh_3_19_io_out_control_0_propagate;
	wire [4:0] _mesh_3_19_io_out_control_0_shift;
	wire [2:0] _mesh_3_19_io_out_id_0;
	wire _mesh_3_19_io_out_last_0;
	wire _mesh_3_19_io_out_valid_0;
	wire [31:0] _mesh_3_18_io_out_a_0;
	wire [31:0] _mesh_3_18_io_out_c_0;
	wire [31:0] _mesh_3_18_io_out_b_0;
	wire _mesh_3_18_io_out_control_0_dataflow;
	wire _mesh_3_18_io_out_control_0_propagate;
	wire [4:0] _mesh_3_18_io_out_control_0_shift;
	wire [2:0] _mesh_3_18_io_out_id_0;
	wire _mesh_3_18_io_out_last_0;
	wire _mesh_3_18_io_out_valid_0;
	wire [31:0] _mesh_3_17_io_out_a_0;
	wire [31:0] _mesh_3_17_io_out_c_0;
	wire [31:0] _mesh_3_17_io_out_b_0;
	wire _mesh_3_17_io_out_control_0_dataflow;
	wire _mesh_3_17_io_out_control_0_propagate;
	wire [4:0] _mesh_3_17_io_out_control_0_shift;
	wire [2:0] _mesh_3_17_io_out_id_0;
	wire _mesh_3_17_io_out_last_0;
	wire _mesh_3_17_io_out_valid_0;
	wire [31:0] _mesh_3_16_io_out_a_0;
	wire [31:0] _mesh_3_16_io_out_c_0;
	wire [31:0] _mesh_3_16_io_out_b_0;
	wire _mesh_3_16_io_out_control_0_dataflow;
	wire _mesh_3_16_io_out_control_0_propagate;
	wire [4:0] _mesh_3_16_io_out_control_0_shift;
	wire [2:0] _mesh_3_16_io_out_id_0;
	wire _mesh_3_16_io_out_last_0;
	wire _mesh_3_16_io_out_valid_0;
	wire [31:0] _mesh_3_15_io_out_a_0;
	wire [31:0] _mesh_3_15_io_out_c_0;
	wire [31:0] _mesh_3_15_io_out_b_0;
	wire _mesh_3_15_io_out_control_0_dataflow;
	wire _mesh_3_15_io_out_control_0_propagate;
	wire [4:0] _mesh_3_15_io_out_control_0_shift;
	wire [2:0] _mesh_3_15_io_out_id_0;
	wire _mesh_3_15_io_out_last_0;
	wire _mesh_3_15_io_out_valid_0;
	wire [31:0] _mesh_3_14_io_out_a_0;
	wire [31:0] _mesh_3_14_io_out_c_0;
	wire [31:0] _mesh_3_14_io_out_b_0;
	wire _mesh_3_14_io_out_control_0_dataflow;
	wire _mesh_3_14_io_out_control_0_propagate;
	wire [4:0] _mesh_3_14_io_out_control_0_shift;
	wire [2:0] _mesh_3_14_io_out_id_0;
	wire _mesh_3_14_io_out_last_0;
	wire _mesh_3_14_io_out_valid_0;
	wire [31:0] _mesh_3_13_io_out_a_0;
	wire [31:0] _mesh_3_13_io_out_c_0;
	wire [31:0] _mesh_3_13_io_out_b_0;
	wire _mesh_3_13_io_out_control_0_dataflow;
	wire _mesh_3_13_io_out_control_0_propagate;
	wire [4:0] _mesh_3_13_io_out_control_0_shift;
	wire [2:0] _mesh_3_13_io_out_id_0;
	wire _mesh_3_13_io_out_last_0;
	wire _mesh_3_13_io_out_valid_0;
	wire [31:0] _mesh_3_12_io_out_a_0;
	wire [31:0] _mesh_3_12_io_out_c_0;
	wire [31:0] _mesh_3_12_io_out_b_0;
	wire _mesh_3_12_io_out_control_0_dataflow;
	wire _mesh_3_12_io_out_control_0_propagate;
	wire [4:0] _mesh_3_12_io_out_control_0_shift;
	wire [2:0] _mesh_3_12_io_out_id_0;
	wire _mesh_3_12_io_out_last_0;
	wire _mesh_3_12_io_out_valid_0;
	wire [31:0] _mesh_3_11_io_out_a_0;
	wire [31:0] _mesh_3_11_io_out_c_0;
	wire [31:0] _mesh_3_11_io_out_b_0;
	wire _mesh_3_11_io_out_control_0_dataflow;
	wire _mesh_3_11_io_out_control_0_propagate;
	wire [4:0] _mesh_3_11_io_out_control_0_shift;
	wire [2:0] _mesh_3_11_io_out_id_0;
	wire _mesh_3_11_io_out_last_0;
	wire _mesh_3_11_io_out_valid_0;
	wire [31:0] _mesh_3_10_io_out_a_0;
	wire [31:0] _mesh_3_10_io_out_c_0;
	wire [31:0] _mesh_3_10_io_out_b_0;
	wire _mesh_3_10_io_out_control_0_dataflow;
	wire _mesh_3_10_io_out_control_0_propagate;
	wire [4:0] _mesh_3_10_io_out_control_0_shift;
	wire [2:0] _mesh_3_10_io_out_id_0;
	wire _mesh_3_10_io_out_last_0;
	wire _mesh_3_10_io_out_valid_0;
	wire [31:0] _mesh_3_9_io_out_a_0;
	wire [31:0] _mesh_3_9_io_out_c_0;
	wire [31:0] _mesh_3_9_io_out_b_0;
	wire _mesh_3_9_io_out_control_0_dataflow;
	wire _mesh_3_9_io_out_control_0_propagate;
	wire [4:0] _mesh_3_9_io_out_control_0_shift;
	wire [2:0] _mesh_3_9_io_out_id_0;
	wire _mesh_3_9_io_out_last_0;
	wire _mesh_3_9_io_out_valid_0;
	wire [31:0] _mesh_3_8_io_out_a_0;
	wire [31:0] _mesh_3_8_io_out_c_0;
	wire [31:0] _mesh_3_8_io_out_b_0;
	wire _mesh_3_8_io_out_control_0_dataflow;
	wire _mesh_3_8_io_out_control_0_propagate;
	wire [4:0] _mesh_3_8_io_out_control_0_shift;
	wire [2:0] _mesh_3_8_io_out_id_0;
	wire _mesh_3_8_io_out_last_0;
	wire _mesh_3_8_io_out_valid_0;
	wire [31:0] _mesh_3_7_io_out_a_0;
	wire [31:0] _mesh_3_7_io_out_c_0;
	wire [31:0] _mesh_3_7_io_out_b_0;
	wire _mesh_3_7_io_out_control_0_dataflow;
	wire _mesh_3_7_io_out_control_0_propagate;
	wire [4:0] _mesh_3_7_io_out_control_0_shift;
	wire [2:0] _mesh_3_7_io_out_id_0;
	wire _mesh_3_7_io_out_last_0;
	wire _mesh_3_7_io_out_valid_0;
	wire [31:0] _mesh_3_6_io_out_a_0;
	wire [31:0] _mesh_3_6_io_out_c_0;
	wire [31:0] _mesh_3_6_io_out_b_0;
	wire _mesh_3_6_io_out_control_0_dataflow;
	wire _mesh_3_6_io_out_control_0_propagate;
	wire [4:0] _mesh_3_6_io_out_control_0_shift;
	wire [2:0] _mesh_3_6_io_out_id_0;
	wire _mesh_3_6_io_out_last_0;
	wire _mesh_3_6_io_out_valid_0;
	wire [31:0] _mesh_3_5_io_out_a_0;
	wire [31:0] _mesh_3_5_io_out_c_0;
	wire [31:0] _mesh_3_5_io_out_b_0;
	wire _mesh_3_5_io_out_control_0_dataflow;
	wire _mesh_3_5_io_out_control_0_propagate;
	wire [4:0] _mesh_3_5_io_out_control_0_shift;
	wire [2:0] _mesh_3_5_io_out_id_0;
	wire _mesh_3_5_io_out_last_0;
	wire _mesh_3_5_io_out_valid_0;
	wire [31:0] _mesh_3_4_io_out_a_0;
	wire [31:0] _mesh_3_4_io_out_c_0;
	wire [31:0] _mesh_3_4_io_out_b_0;
	wire _mesh_3_4_io_out_control_0_dataflow;
	wire _mesh_3_4_io_out_control_0_propagate;
	wire [4:0] _mesh_3_4_io_out_control_0_shift;
	wire [2:0] _mesh_3_4_io_out_id_0;
	wire _mesh_3_4_io_out_last_0;
	wire _mesh_3_4_io_out_valid_0;
	wire [31:0] _mesh_3_3_io_out_a_0;
	wire [31:0] _mesh_3_3_io_out_c_0;
	wire [31:0] _mesh_3_3_io_out_b_0;
	wire _mesh_3_3_io_out_control_0_dataflow;
	wire _mesh_3_3_io_out_control_0_propagate;
	wire [4:0] _mesh_3_3_io_out_control_0_shift;
	wire [2:0] _mesh_3_3_io_out_id_0;
	wire _mesh_3_3_io_out_last_0;
	wire _mesh_3_3_io_out_valid_0;
	wire [31:0] _mesh_3_2_io_out_a_0;
	wire [31:0] _mesh_3_2_io_out_c_0;
	wire [31:0] _mesh_3_2_io_out_b_0;
	wire _mesh_3_2_io_out_control_0_dataflow;
	wire _mesh_3_2_io_out_control_0_propagate;
	wire [4:0] _mesh_3_2_io_out_control_0_shift;
	wire [2:0] _mesh_3_2_io_out_id_0;
	wire _mesh_3_2_io_out_last_0;
	wire _mesh_3_2_io_out_valid_0;
	wire [31:0] _mesh_3_1_io_out_a_0;
	wire [31:0] _mesh_3_1_io_out_c_0;
	wire [31:0] _mesh_3_1_io_out_b_0;
	wire _mesh_3_1_io_out_control_0_dataflow;
	wire _mesh_3_1_io_out_control_0_propagate;
	wire [4:0] _mesh_3_1_io_out_control_0_shift;
	wire [2:0] _mesh_3_1_io_out_id_0;
	wire _mesh_3_1_io_out_last_0;
	wire _mesh_3_1_io_out_valid_0;
	wire [31:0] _mesh_3_0_io_out_a_0;
	wire [31:0] _mesh_3_0_io_out_c_0;
	wire [31:0] _mesh_3_0_io_out_b_0;
	wire _mesh_3_0_io_out_control_0_dataflow;
	wire _mesh_3_0_io_out_control_0_propagate;
	wire [4:0] _mesh_3_0_io_out_control_0_shift;
	wire [2:0] _mesh_3_0_io_out_id_0;
	wire _mesh_3_0_io_out_last_0;
	wire _mesh_3_0_io_out_valid_0;
	wire [31:0] _mesh_2_31_io_out_a_0;
	wire [31:0] _mesh_2_31_io_out_c_0;
	wire [31:0] _mesh_2_31_io_out_b_0;
	wire _mesh_2_31_io_out_control_0_dataflow;
	wire _mesh_2_31_io_out_control_0_propagate;
	wire [4:0] _mesh_2_31_io_out_control_0_shift;
	wire [2:0] _mesh_2_31_io_out_id_0;
	wire _mesh_2_31_io_out_last_0;
	wire _mesh_2_31_io_out_valid_0;
	wire [31:0] _mesh_2_30_io_out_a_0;
	wire [31:0] _mesh_2_30_io_out_c_0;
	wire [31:0] _mesh_2_30_io_out_b_0;
	wire _mesh_2_30_io_out_control_0_dataflow;
	wire _mesh_2_30_io_out_control_0_propagate;
	wire [4:0] _mesh_2_30_io_out_control_0_shift;
	wire [2:0] _mesh_2_30_io_out_id_0;
	wire _mesh_2_30_io_out_last_0;
	wire _mesh_2_30_io_out_valid_0;
	wire [31:0] _mesh_2_29_io_out_a_0;
	wire [31:0] _mesh_2_29_io_out_c_0;
	wire [31:0] _mesh_2_29_io_out_b_0;
	wire _mesh_2_29_io_out_control_0_dataflow;
	wire _mesh_2_29_io_out_control_0_propagate;
	wire [4:0] _mesh_2_29_io_out_control_0_shift;
	wire [2:0] _mesh_2_29_io_out_id_0;
	wire _mesh_2_29_io_out_last_0;
	wire _mesh_2_29_io_out_valid_0;
	wire [31:0] _mesh_2_28_io_out_a_0;
	wire [31:0] _mesh_2_28_io_out_c_0;
	wire [31:0] _mesh_2_28_io_out_b_0;
	wire _mesh_2_28_io_out_control_0_dataflow;
	wire _mesh_2_28_io_out_control_0_propagate;
	wire [4:0] _mesh_2_28_io_out_control_0_shift;
	wire [2:0] _mesh_2_28_io_out_id_0;
	wire _mesh_2_28_io_out_last_0;
	wire _mesh_2_28_io_out_valid_0;
	wire [31:0] _mesh_2_27_io_out_a_0;
	wire [31:0] _mesh_2_27_io_out_c_0;
	wire [31:0] _mesh_2_27_io_out_b_0;
	wire _mesh_2_27_io_out_control_0_dataflow;
	wire _mesh_2_27_io_out_control_0_propagate;
	wire [4:0] _mesh_2_27_io_out_control_0_shift;
	wire [2:0] _mesh_2_27_io_out_id_0;
	wire _mesh_2_27_io_out_last_0;
	wire _mesh_2_27_io_out_valid_0;
	wire [31:0] _mesh_2_26_io_out_a_0;
	wire [31:0] _mesh_2_26_io_out_c_0;
	wire [31:0] _mesh_2_26_io_out_b_0;
	wire _mesh_2_26_io_out_control_0_dataflow;
	wire _mesh_2_26_io_out_control_0_propagate;
	wire [4:0] _mesh_2_26_io_out_control_0_shift;
	wire [2:0] _mesh_2_26_io_out_id_0;
	wire _mesh_2_26_io_out_last_0;
	wire _mesh_2_26_io_out_valid_0;
	wire [31:0] _mesh_2_25_io_out_a_0;
	wire [31:0] _mesh_2_25_io_out_c_0;
	wire [31:0] _mesh_2_25_io_out_b_0;
	wire _mesh_2_25_io_out_control_0_dataflow;
	wire _mesh_2_25_io_out_control_0_propagate;
	wire [4:0] _mesh_2_25_io_out_control_0_shift;
	wire [2:0] _mesh_2_25_io_out_id_0;
	wire _mesh_2_25_io_out_last_0;
	wire _mesh_2_25_io_out_valid_0;
	wire [31:0] _mesh_2_24_io_out_a_0;
	wire [31:0] _mesh_2_24_io_out_c_0;
	wire [31:0] _mesh_2_24_io_out_b_0;
	wire _mesh_2_24_io_out_control_0_dataflow;
	wire _mesh_2_24_io_out_control_0_propagate;
	wire [4:0] _mesh_2_24_io_out_control_0_shift;
	wire [2:0] _mesh_2_24_io_out_id_0;
	wire _mesh_2_24_io_out_last_0;
	wire _mesh_2_24_io_out_valid_0;
	wire [31:0] _mesh_2_23_io_out_a_0;
	wire [31:0] _mesh_2_23_io_out_c_0;
	wire [31:0] _mesh_2_23_io_out_b_0;
	wire _mesh_2_23_io_out_control_0_dataflow;
	wire _mesh_2_23_io_out_control_0_propagate;
	wire [4:0] _mesh_2_23_io_out_control_0_shift;
	wire [2:0] _mesh_2_23_io_out_id_0;
	wire _mesh_2_23_io_out_last_0;
	wire _mesh_2_23_io_out_valid_0;
	wire [31:0] _mesh_2_22_io_out_a_0;
	wire [31:0] _mesh_2_22_io_out_c_0;
	wire [31:0] _mesh_2_22_io_out_b_0;
	wire _mesh_2_22_io_out_control_0_dataflow;
	wire _mesh_2_22_io_out_control_0_propagate;
	wire [4:0] _mesh_2_22_io_out_control_0_shift;
	wire [2:0] _mesh_2_22_io_out_id_0;
	wire _mesh_2_22_io_out_last_0;
	wire _mesh_2_22_io_out_valid_0;
	wire [31:0] _mesh_2_21_io_out_a_0;
	wire [31:0] _mesh_2_21_io_out_c_0;
	wire [31:0] _mesh_2_21_io_out_b_0;
	wire _mesh_2_21_io_out_control_0_dataflow;
	wire _mesh_2_21_io_out_control_0_propagate;
	wire [4:0] _mesh_2_21_io_out_control_0_shift;
	wire [2:0] _mesh_2_21_io_out_id_0;
	wire _mesh_2_21_io_out_last_0;
	wire _mesh_2_21_io_out_valid_0;
	wire [31:0] _mesh_2_20_io_out_a_0;
	wire [31:0] _mesh_2_20_io_out_c_0;
	wire [31:0] _mesh_2_20_io_out_b_0;
	wire _mesh_2_20_io_out_control_0_dataflow;
	wire _mesh_2_20_io_out_control_0_propagate;
	wire [4:0] _mesh_2_20_io_out_control_0_shift;
	wire [2:0] _mesh_2_20_io_out_id_0;
	wire _mesh_2_20_io_out_last_0;
	wire _mesh_2_20_io_out_valid_0;
	wire [31:0] _mesh_2_19_io_out_a_0;
	wire [31:0] _mesh_2_19_io_out_c_0;
	wire [31:0] _mesh_2_19_io_out_b_0;
	wire _mesh_2_19_io_out_control_0_dataflow;
	wire _mesh_2_19_io_out_control_0_propagate;
	wire [4:0] _mesh_2_19_io_out_control_0_shift;
	wire [2:0] _mesh_2_19_io_out_id_0;
	wire _mesh_2_19_io_out_last_0;
	wire _mesh_2_19_io_out_valid_0;
	wire [31:0] _mesh_2_18_io_out_a_0;
	wire [31:0] _mesh_2_18_io_out_c_0;
	wire [31:0] _mesh_2_18_io_out_b_0;
	wire _mesh_2_18_io_out_control_0_dataflow;
	wire _mesh_2_18_io_out_control_0_propagate;
	wire [4:0] _mesh_2_18_io_out_control_0_shift;
	wire [2:0] _mesh_2_18_io_out_id_0;
	wire _mesh_2_18_io_out_last_0;
	wire _mesh_2_18_io_out_valid_0;
	wire [31:0] _mesh_2_17_io_out_a_0;
	wire [31:0] _mesh_2_17_io_out_c_0;
	wire [31:0] _mesh_2_17_io_out_b_0;
	wire _mesh_2_17_io_out_control_0_dataflow;
	wire _mesh_2_17_io_out_control_0_propagate;
	wire [4:0] _mesh_2_17_io_out_control_0_shift;
	wire [2:0] _mesh_2_17_io_out_id_0;
	wire _mesh_2_17_io_out_last_0;
	wire _mesh_2_17_io_out_valid_0;
	wire [31:0] _mesh_2_16_io_out_a_0;
	wire [31:0] _mesh_2_16_io_out_c_0;
	wire [31:0] _mesh_2_16_io_out_b_0;
	wire _mesh_2_16_io_out_control_0_dataflow;
	wire _mesh_2_16_io_out_control_0_propagate;
	wire [4:0] _mesh_2_16_io_out_control_0_shift;
	wire [2:0] _mesh_2_16_io_out_id_0;
	wire _mesh_2_16_io_out_last_0;
	wire _mesh_2_16_io_out_valid_0;
	wire [31:0] _mesh_2_15_io_out_a_0;
	wire [31:0] _mesh_2_15_io_out_c_0;
	wire [31:0] _mesh_2_15_io_out_b_0;
	wire _mesh_2_15_io_out_control_0_dataflow;
	wire _mesh_2_15_io_out_control_0_propagate;
	wire [4:0] _mesh_2_15_io_out_control_0_shift;
	wire [2:0] _mesh_2_15_io_out_id_0;
	wire _mesh_2_15_io_out_last_0;
	wire _mesh_2_15_io_out_valid_0;
	wire [31:0] _mesh_2_14_io_out_a_0;
	wire [31:0] _mesh_2_14_io_out_c_0;
	wire [31:0] _mesh_2_14_io_out_b_0;
	wire _mesh_2_14_io_out_control_0_dataflow;
	wire _mesh_2_14_io_out_control_0_propagate;
	wire [4:0] _mesh_2_14_io_out_control_0_shift;
	wire [2:0] _mesh_2_14_io_out_id_0;
	wire _mesh_2_14_io_out_last_0;
	wire _mesh_2_14_io_out_valid_0;
	wire [31:0] _mesh_2_13_io_out_a_0;
	wire [31:0] _mesh_2_13_io_out_c_0;
	wire [31:0] _mesh_2_13_io_out_b_0;
	wire _mesh_2_13_io_out_control_0_dataflow;
	wire _mesh_2_13_io_out_control_0_propagate;
	wire [4:0] _mesh_2_13_io_out_control_0_shift;
	wire [2:0] _mesh_2_13_io_out_id_0;
	wire _mesh_2_13_io_out_last_0;
	wire _mesh_2_13_io_out_valid_0;
	wire [31:0] _mesh_2_12_io_out_a_0;
	wire [31:0] _mesh_2_12_io_out_c_0;
	wire [31:0] _mesh_2_12_io_out_b_0;
	wire _mesh_2_12_io_out_control_0_dataflow;
	wire _mesh_2_12_io_out_control_0_propagate;
	wire [4:0] _mesh_2_12_io_out_control_0_shift;
	wire [2:0] _mesh_2_12_io_out_id_0;
	wire _mesh_2_12_io_out_last_0;
	wire _mesh_2_12_io_out_valid_0;
	wire [31:0] _mesh_2_11_io_out_a_0;
	wire [31:0] _mesh_2_11_io_out_c_0;
	wire [31:0] _mesh_2_11_io_out_b_0;
	wire _mesh_2_11_io_out_control_0_dataflow;
	wire _mesh_2_11_io_out_control_0_propagate;
	wire [4:0] _mesh_2_11_io_out_control_0_shift;
	wire [2:0] _mesh_2_11_io_out_id_0;
	wire _mesh_2_11_io_out_last_0;
	wire _mesh_2_11_io_out_valid_0;
	wire [31:0] _mesh_2_10_io_out_a_0;
	wire [31:0] _mesh_2_10_io_out_c_0;
	wire [31:0] _mesh_2_10_io_out_b_0;
	wire _mesh_2_10_io_out_control_0_dataflow;
	wire _mesh_2_10_io_out_control_0_propagate;
	wire [4:0] _mesh_2_10_io_out_control_0_shift;
	wire [2:0] _mesh_2_10_io_out_id_0;
	wire _mesh_2_10_io_out_last_0;
	wire _mesh_2_10_io_out_valid_0;
	wire [31:0] _mesh_2_9_io_out_a_0;
	wire [31:0] _mesh_2_9_io_out_c_0;
	wire [31:0] _mesh_2_9_io_out_b_0;
	wire _mesh_2_9_io_out_control_0_dataflow;
	wire _mesh_2_9_io_out_control_0_propagate;
	wire [4:0] _mesh_2_9_io_out_control_0_shift;
	wire [2:0] _mesh_2_9_io_out_id_0;
	wire _mesh_2_9_io_out_last_0;
	wire _mesh_2_9_io_out_valid_0;
	wire [31:0] _mesh_2_8_io_out_a_0;
	wire [31:0] _mesh_2_8_io_out_c_0;
	wire [31:0] _mesh_2_8_io_out_b_0;
	wire _mesh_2_8_io_out_control_0_dataflow;
	wire _mesh_2_8_io_out_control_0_propagate;
	wire [4:0] _mesh_2_8_io_out_control_0_shift;
	wire [2:0] _mesh_2_8_io_out_id_0;
	wire _mesh_2_8_io_out_last_0;
	wire _mesh_2_8_io_out_valid_0;
	wire [31:0] _mesh_2_7_io_out_a_0;
	wire [31:0] _mesh_2_7_io_out_c_0;
	wire [31:0] _mesh_2_7_io_out_b_0;
	wire _mesh_2_7_io_out_control_0_dataflow;
	wire _mesh_2_7_io_out_control_0_propagate;
	wire [4:0] _mesh_2_7_io_out_control_0_shift;
	wire [2:0] _mesh_2_7_io_out_id_0;
	wire _mesh_2_7_io_out_last_0;
	wire _mesh_2_7_io_out_valid_0;
	wire [31:0] _mesh_2_6_io_out_a_0;
	wire [31:0] _mesh_2_6_io_out_c_0;
	wire [31:0] _mesh_2_6_io_out_b_0;
	wire _mesh_2_6_io_out_control_0_dataflow;
	wire _mesh_2_6_io_out_control_0_propagate;
	wire [4:0] _mesh_2_6_io_out_control_0_shift;
	wire [2:0] _mesh_2_6_io_out_id_0;
	wire _mesh_2_6_io_out_last_0;
	wire _mesh_2_6_io_out_valid_0;
	wire [31:0] _mesh_2_5_io_out_a_0;
	wire [31:0] _mesh_2_5_io_out_c_0;
	wire [31:0] _mesh_2_5_io_out_b_0;
	wire _mesh_2_5_io_out_control_0_dataflow;
	wire _mesh_2_5_io_out_control_0_propagate;
	wire [4:0] _mesh_2_5_io_out_control_0_shift;
	wire [2:0] _mesh_2_5_io_out_id_0;
	wire _mesh_2_5_io_out_last_0;
	wire _mesh_2_5_io_out_valid_0;
	wire [31:0] _mesh_2_4_io_out_a_0;
	wire [31:0] _mesh_2_4_io_out_c_0;
	wire [31:0] _mesh_2_4_io_out_b_0;
	wire _mesh_2_4_io_out_control_0_dataflow;
	wire _mesh_2_4_io_out_control_0_propagate;
	wire [4:0] _mesh_2_4_io_out_control_0_shift;
	wire [2:0] _mesh_2_4_io_out_id_0;
	wire _mesh_2_4_io_out_last_0;
	wire _mesh_2_4_io_out_valid_0;
	wire [31:0] _mesh_2_3_io_out_a_0;
	wire [31:0] _mesh_2_3_io_out_c_0;
	wire [31:0] _mesh_2_3_io_out_b_0;
	wire _mesh_2_3_io_out_control_0_dataflow;
	wire _mesh_2_3_io_out_control_0_propagate;
	wire [4:0] _mesh_2_3_io_out_control_0_shift;
	wire [2:0] _mesh_2_3_io_out_id_0;
	wire _mesh_2_3_io_out_last_0;
	wire _mesh_2_3_io_out_valid_0;
	wire [31:0] _mesh_2_2_io_out_a_0;
	wire [31:0] _mesh_2_2_io_out_c_0;
	wire [31:0] _mesh_2_2_io_out_b_0;
	wire _mesh_2_2_io_out_control_0_dataflow;
	wire _mesh_2_2_io_out_control_0_propagate;
	wire [4:0] _mesh_2_2_io_out_control_0_shift;
	wire [2:0] _mesh_2_2_io_out_id_0;
	wire _mesh_2_2_io_out_last_0;
	wire _mesh_2_2_io_out_valid_0;
	wire [31:0] _mesh_2_1_io_out_a_0;
	wire [31:0] _mesh_2_1_io_out_c_0;
	wire [31:0] _mesh_2_1_io_out_b_0;
	wire _mesh_2_1_io_out_control_0_dataflow;
	wire _mesh_2_1_io_out_control_0_propagate;
	wire [4:0] _mesh_2_1_io_out_control_0_shift;
	wire [2:0] _mesh_2_1_io_out_id_0;
	wire _mesh_2_1_io_out_last_0;
	wire _mesh_2_1_io_out_valid_0;
	wire [31:0] _mesh_2_0_io_out_a_0;
	wire [31:0] _mesh_2_0_io_out_c_0;
	wire [31:0] _mesh_2_0_io_out_b_0;
	wire _mesh_2_0_io_out_control_0_dataflow;
	wire _mesh_2_0_io_out_control_0_propagate;
	wire [4:0] _mesh_2_0_io_out_control_0_shift;
	wire [2:0] _mesh_2_0_io_out_id_0;
	wire _mesh_2_0_io_out_last_0;
	wire _mesh_2_0_io_out_valid_0;
	wire [31:0] _mesh_1_31_io_out_a_0;
	wire [31:0] _mesh_1_31_io_out_c_0;
	wire [31:0] _mesh_1_31_io_out_b_0;
	wire _mesh_1_31_io_out_control_0_dataflow;
	wire _mesh_1_31_io_out_control_0_propagate;
	wire [4:0] _mesh_1_31_io_out_control_0_shift;
	wire [2:0] _mesh_1_31_io_out_id_0;
	wire _mesh_1_31_io_out_last_0;
	wire _mesh_1_31_io_out_valid_0;
	wire [31:0] _mesh_1_30_io_out_a_0;
	wire [31:0] _mesh_1_30_io_out_c_0;
	wire [31:0] _mesh_1_30_io_out_b_0;
	wire _mesh_1_30_io_out_control_0_dataflow;
	wire _mesh_1_30_io_out_control_0_propagate;
	wire [4:0] _mesh_1_30_io_out_control_0_shift;
	wire [2:0] _mesh_1_30_io_out_id_0;
	wire _mesh_1_30_io_out_last_0;
	wire _mesh_1_30_io_out_valid_0;
	wire [31:0] _mesh_1_29_io_out_a_0;
	wire [31:0] _mesh_1_29_io_out_c_0;
	wire [31:0] _mesh_1_29_io_out_b_0;
	wire _mesh_1_29_io_out_control_0_dataflow;
	wire _mesh_1_29_io_out_control_0_propagate;
	wire [4:0] _mesh_1_29_io_out_control_0_shift;
	wire [2:0] _mesh_1_29_io_out_id_0;
	wire _mesh_1_29_io_out_last_0;
	wire _mesh_1_29_io_out_valid_0;
	wire [31:0] _mesh_1_28_io_out_a_0;
	wire [31:0] _mesh_1_28_io_out_c_0;
	wire [31:0] _mesh_1_28_io_out_b_0;
	wire _mesh_1_28_io_out_control_0_dataflow;
	wire _mesh_1_28_io_out_control_0_propagate;
	wire [4:0] _mesh_1_28_io_out_control_0_shift;
	wire [2:0] _mesh_1_28_io_out_id_0;
	wire _mesh_1_28_io_out_last_0;
	wire _mesh_1_28_io_out_valid_0;
	wire [31:0] _mesh_1_27_io_out_a_0;
	wire [31:0] _mesh_1_27_io_out_c_0;
	wire [31:0] _mesh_1_27_io_out_b_0;
	wire _mesh_1_27_io_out_control_0_dataflow;
	wire _mesh_1_27_io_out_control_0_propagate;
	wire [4:0] _mesh_1_27_io_out_control_0_shift;
	wire [2:0] _mesh_1_27_io_out_id_0;
	wire _mesh_1_27_io_out_last_0;
	wire _mesh_1_27_io_out_valid_0;
	wire [31:0] _mesh_1_26_io_out_a_0;
	wire [31:0] _mesh_1_26_io_out_c_0;
	wire [31:0] _mesh_1_26_io_out_b_0;
	wire _mesh_1_26_io_out_control_0_dataflow;
	wire _mesh_1_26_io_out_control_0_propagate;
	wire [4:0] _mesh_1_26_io_out_control_0_shift;
	wire [2:0] _mesh_1_26_io_out_id_0;
	wire _mesh_1_26_io_out_last_0;
	wire _mesh_1_26_io_out_valid_0;
	wire [31:0] _mesh_1_25_io_out_a_0;
	wire [31:0] _mesh_1_25_io_out_c_0;
	wire [31:0] _mesh_1_25_io_out_b_0;
	wire _mesh_1_25_io_out_control_0_dataflow;
	wire _mesh_1_25_io_out_control_0_propagate;
	wire [4:0] _mesh_1_25_io_out_control_0_shift;
	wire [2:0] _mesh_1_25_io_out_id_0;
	wire _mesh_1_25_io_out_last_0;
	wire _mesh_1_25_io_out_valid_0;
	wire [31:0] _mesh_1_24_io_out_a_0;
	wire [31:0] _mesh_1_24_io_out_c_0;
	wire [31:0] _mesh_1_24_io_out_b_0;
	wire _mesh_1_24_io_out_control_0_dataflow;
	wire _mesh_1_24_io_out_control_0_propagate;
	wire [4:0] _mesh_1_24_io_out_control_0_shift;
	wire [2:0] _mesh_1_24_io_out_id_0;
	wire _mesh_1_24_io_out_last_0;
	wire _mesh_1_24_io_out_valid_0;
	wire [31:0] _mesh_1_23_io_out_a_0;
	wire [31:0] _mesh_1_23_io_out_c_0;
	wire [31:0] _mesh_1_23_io_out_b_0;
	wire _mesh_1_23_io_out_control_0_dataflow;
	wire _mesh_1_23_io_out_control_0_propagate;
	wire [4:0] _mesh_1_23_io_out_control_0_shift;
	wire [2:0] _mesh_1_23_io_out_id_0;
	wire _mesh_1_23_io_out_last_0;
	wire _mesh_1_23_io_out_valid_0;
	wire [31:0] _mesh_1_22_io_out_a_0;
	wire [31:0] _mesh_1_22_io_out_c_0;
	wire [31:0] _mesh_1_22_io_out_b_0;
	wire _mesh_1_22_io_out_control_0_dataflow;
	wire _mesh_1_22_io_out_control_0_propagate;
	wire [4:0] _mesh_1_22_io_out_control_0_shift;
	wire [2:0] _mesh_1_22_io_out_id_0;
	wire _mesh_1_22_io_out_last_0;
	wire _mesh_1_22_io_out_valid_0;
	wire [31:0] _mesh_1_21_io_out_a_0;
	wire [31:0] _mesh_1_21_io_out_c_0;
	wire [31:0] _mesh_1_21_io_out_b_0;
	wire _mesh_1_21_io_out_control_0_dataflow;
	wire _mesh_1_21_io_out_control_0_propagate;
	wire [4:0] _mesh_1_21_io_out_control_0_shift;
	wire [2:0] _mesh_1_21_io_out_id_0;
	wire _mesh_1_21_io_out_last_0;
	wire _mesh_1_21_io_out_valid_0;
	wire [31:0] _mesh_1_20_io_out_a_0;
	wire [31:0] _mesh_1_20_io_out_c_0;
	wire [31:0] _mesh_1_20_io_out_b_0;
	wire _mesh_1_20_io_out_control_0_dataflow;
	wire _mesh_1_20_io_out_control_0_propagate;
	wire [4:0] _mesh_1_20_io_out_control_0_shift;
	wire [2:0] _mesh_1_20_io_out_id_0;
	wire _mesh_1_20_io_out_last_0;
	wire _mesh_1_20_io_out_valid_0;
	wire [31:0] _mesh_1_19_io_out_a_0;
	wire [31:0] _mesh_1_19_io_out_c_0;
	wire [31:0] _mesh_1_19_io_out_b_0;
	wire _mesh_1_19_io_out_control_0_dataflow;
	wire _mesh_1_19_io_out_control_0_propagate;
	wire [4:0] _mesh_1_19_io_out_control_0_shift;
	wire [2:0] _mesh_1_19_io_out_id_0;
	wire _mesh_1_19_io_out_last_0;
	wire _mesh_1_19_io_out_valid_0;
	wire [31:0] _mesh_1_18_io_out_a_0;
	wire [31:0] _mesh_1_18_io_out_c_0;
	wire [31:0] _mesh_1_18_io_out_b_0;
	wire _mesh_1_18_io_out_control_0_dataflow;
	wire _mesh_1_18_io_out_control_0_propagate;
	wire [4:0] _mesh_1_18_io_out_control_0_shift;
	wire [2:0] _mesh_1_18_io_out_id_0;
	wire _mesh_1_18_io_out_last_0;
	wire _mesh_1_18_io_out_valid_0;
	wire [31:0] _mesh_1_17_io_out_a_0;
	wire [31:0] _mesh_1_17_io_out_c_0;
	wire [31:0] _mesh_1_17_io_out_b_0;
	wire _mesh_1_17_io_out_control_0_dataflow;
	wire _mesh_1_17_io_out_control_0_propagate;
	wire [4:0] _mesh_1_17_io_out_control_0_shift;
	wire [2:0] _mesh_1_17_io_out_id_0;
	wire _mesh_1_17_io_out_last_0;
	wire _mesh_1_17_io_out_valid_0;
	wire [31:0] _mesh_1_16_io_out_a_0;
	wire [31:0] _mesh_1_16_io_out_c_0;
	wire [31:0] _mesh_1_16_io_out_b_0;
	wire _mesh_1_16_io_out_control_0_dataflow;
	wire _mesh_1_16_io_out_control_0_propagate;
	wire [4:0] _mesh_1_16_io_out_control_0_shift;
	wire [2:0] _mesh_1_16_io_out_id_0;
	wire _mesh_1_16_io_out_last_0;
	wire _mesh_1_16_io_out_valid_0;
	wire [31:0] _mesh_1_15_io_out_a_0;
	wire [31:0] _mesh_1_15_io_out_c_0;
	wire [31:0] _mesh_1_15_io_out_b_0;
	wire _mesh_1_15_io_out_control_0_dataflow;
	wire _mesh_1_15_io_out_control_0_propagate;
	wire [4:0] _mesh_1_15_io_out_control_0_shift;
	wire [2:0] _mesh_1_15_io_out_id_0;
	wire _mesh_1_15_io_out_last_0;
	wire _mesh_1_15_io_out_valid_0;
	wire [31:0] _mesh_1_14_io_out_a_0;
	wire [31:0] _mesh_1_14_io_out_c_0;
	wire [31:0] _mesh_1_14_io_out_b_0;
	wire _mesh_1_14_io_out_control_0_dataflow;
	wire _mesh_1_14_io_out_control_0_propagate;
	wire [4:0] _mesh_1_14_io_out_control_0_shift;
	wire [2:0] _mesh_1_14_io_out_id_0;
	wire _mesh_1_14_io_out_last_0;
	wire _mesh_1_14_io_out_valid_0;
	wire [31:0] _mesh_1_13_io_out_a_0;
	wire [31:0] _mesh_1_13_io_out_c_0;
	wire [31:0] _mesh_1_13_io_out_b_0;
	wire _mesh_1_13_io_out_control_0_dataflow;
	wire _mesh_1_13_io_out_control_0_propagate;
	wire [4:0] _mesh_1_13_io_out_control_0_shift;
	wire [2:0] _mesh_1_13_io_out_id_0;
	wire _mesh_1_13_io_out_last_0;
	wire _mesh_1_13_io_out_valid_0;
	wire [31:0] _mesh_1_12_io_out_a_0;
	wire [31:0] _mesh_1_12_io_out_c_0;
	wire [31:0] _mesh_1_12_io_out_b_0;
	wire _mesh_1_12_io_out_control_0_dataflow;
	wire _mesh_1_12_io_out_control_0_propagate;
	wire [4:0] _mesh_1_12_io_out_control_0_shift;
	wire [2:0] _mesh_1_12_io_out_id_0;
	wire _mesh_1_12_io_out_last_0;
	wire _mesh_1_12_io_out_valid_0;
	wire [31:0] _mesh_1_11_io_out_a_0;
	wire [31:0] _mesh_1_11_io_out_c_0;
	wire [31:0] _mesh_1_11_io_out_b_0;
	wire _mesh_1_11_io_out_control_0_dataflow;
	wire _mesh_1_11_io_out_control_0_propagate;
	wire [4:0] _mesh_1_11_io_out_control_0_shift;
	wire [2:0] _mesh_1_11_io_out_id_0;
	wire _mesh_1_11_io_out_last_0;
	wire _mesh_1_11_io_out_valid_0;
	wire [31:0] _mesh_1_10_io_out_a_0;
	wire [31:0] _mesh_1_10_io_out_c_0;
	wire [31:0] _mesh_1_10_io_out_b_0;
	wire _mesh_1_10_io_out_control_0_dataflow;
	wire _mesh_1_10_io_out_control_0_propagate;
	wire [4:0] _mesh_1_10_io_out_control_0_shift;
	wire [2:0] _mesh_1_10_io_out_id_0;
	wire _mesh_1_10_io_out_last_0;
	wire _mesh_1_10_io_out_valid_0;
	wire [31:0] _mesh_1_9_io_out_a_0;
	wire [31:0] _mesh_1_9_io_out_c_0;
	wire [31:0] _mesh_1_9_io_out_b_0;
	wire _mesh_1_9_io_out_control_0_dataflow;
	wire _mesh_1_9_io_out_control_0_propagate;
	wire [4:0] _mesh_1_9_io_out_control_0_shift;
	wire [2:0] _mesh_1_9_io_out_id_0;
	wire _mesh_1_9_io_out_last_0;
	wire _mesh_1_9_io_out_valid_0;
	wire [31:0] _mesh_1_8_io_out_a_0;
	wire [31:0] _mesh_1_8_io_out_c_0;
	wire [31:0] _mesh_1_8_io_out_b_0;
	wire _mesh_1_8_io_out_control_0_dataflow;
	wire _mesh_1_8_io_out_control_0_propagate;
	wire [4:0] _mesh_1_8_io_out_control_0_shift;
	wire [2:0] _mesh_1_8_io_out_id_0;
	wire _mesh_1_8_io_out_last_0;
	wire _mesh_1_8_io_out_valid_0;
	wire [31:0] _mesh_1_7_io_out_a_0;
	wire [31:0] _mesh_1_7_io_out_c_0;
	wire [31:0] _mesh_1_7_io_out_b_0;
	wire _mesh_1_7_io_out_control_0_dataflow;
	wire _mesh_1_7_io_out_control_0_propagate;
	wire [4:0] _mesh_1_7_io_out_control_0_shift;
	wire [2:0] _mesh_1_7_io_out_id_0;
	wire _mesh_1_7_io_out_last_0;
	wire _mesh_1_7_io_out_valid_0;
	wire [31:0] _mesh_1_6_io_out_a_0;
	wire [31:0] _mesh_1_6_io_out_c_0;
	wire [31:0] _mesh_1_6_io_out_b_0;
	wire _mesh_1_6_io_out_control_0_dataflow;
	wire _mesh_1_6_io_out_control_0_propagate;
	wire [4:0] _mesh_1_6_io_out_control_0_shift;
	wire [2:0] _mesh_1_6_io_out_id_0;
	wire _mesh_1_6_io_out_last_0;
	wire _mesh_1_6_io_out_valid_0;
	wire [31:0] _mesh_1_5_io_out_a_0;
	wire [31:0] _mesh_1_5_io_out_c_0;
	wire [31:0] _mesh_1_5_io_out_b_0;
	wire _mesh_1_5_io_out_control_0_dataflow;
	wire _mesh_1_5_io_out_control_0_propagate;
	wire [4:0] _mesh_1_5_io_out_control_0_shift;
	wire [2:0] _mesh_1_5_io_out_id_0;
	wire _mesh_1_5_io_out_last_0;
	wire _mesh_1_5_io_out_valid_0;
	wire [31:0] _mesh_1_4_io_out_a_0;
	wire [31:0] _mesh_1_4_io_out_c_0;
	wire [31:0] _mesh_1_4_io_out_b_0;
	wire _mesh_1_4_io_out_control_0_dataflow;
	wire _mesh_1_4_io_out_control_0_propagate;
	wire [4:0] _mesh_1_4_io_out_control_0_shift;
	wire [2:0] _mesh_1_4_io_out_id_0;
	wire _mesh_1_4_io_out_last_0;
	wire _mesh_1_4_io_out_valid_0;
	wire [31:0] _mesh_1_3_io_out_a_0;
	wire [31:0] _mesh_1_3_io_out_c_0;
	wire [31:0] _mesh_1_3_io_out_b_0;
	wire _mesh_1_3_io_out_control_0_dataflow;
	wire _mesh_1_3_io_out_control_0_propagate;
	wire [4:0] _mesh_1_3_io_out_control_0_shift;
	wire [2:0] _mesh_1_3_io_out_id_0;
	wire _mesh_1_3_io_out_last_0;
	wire _mesh_1_3_io_out_valid_0;
	wire [31:0] _mesh_1_2_io_out_a_0;
	wire [31:0] _mesh_1_2_io_out_c_0;
	wire [31:0] _mesh_1_2_io_out_b_0;
	wire _mesh_1_2_io_out_control_0_dataflow;
	wire _mesh_1_2_io_out_control_0_propagate;
	wire [4:0] _mesh_1_2_io_out_control_0_shift;
	wire [2:0] _mesh_1_2_io_out_id_0;
	wire _mesh_1_2_io_out_last_0;
	wire _mesh_1_2_io_out_valid_0;
	wire [31:0] _mesh_1_1_io_out_a_0;
	wire [31:0] _mesh_1_1_io_out_c_0;
	wire [31:0] _mesh_1_1_io_out_b_0;
	wire _mesh_1_1_io_out_control_0_dataflow;
	wire _mesh_1_1_io_out_control_0_propagate;
	wire [4:0] _mesh_1_1_io_out_control_0_shift;
	wire [2:0] _mesh_1_1_io_out_id_0;
	wire _mesh_1_1_io_out_last_0;
	wire _mesh_1_1_io_out_valid_0;
	wire [31:0] _mesh_1_0_io_out_a_0;
	wire [31:0] _mesh_1_0_io_out_c_0;
	wire [31:0] _mesh_1_0_io_out_b_0;
	wire _mesh_1_0_io_out_control_0_dataflow;
	wire _mesh_1_0_io_out_control_0_propagate;
	wire [4:0] _mesh_1_0_io_out_control_0_shift;
	wire [2:0] _mesh_1_0_io_out_id_0;
	wire _mesh_1_0_io_out_last_0;
	wire _mesh_1_0_io_out_valid_0;
	wire [31:0] _mesh_0_31_io_out_a_0;
	wire [31:0] _mesh_0_31_io_out_c_0;
	wire [31:0] _mesh_0_31_io_out_b_0;
	wire _mesh_0_31_io_out_control_0_dataflow;
	wire _mesh_0_31_io_out_control_0_propagate;
	wire [4:0] _mesh_0_31_io_out_control_0_shift;
	wire [2:0] _mesh_0_31_io_out_id_0;
	wire _mesh_0_31_io_out_last_0;
	wire _mesh_0_31_io_out_valid_0;
	wire [31:0] _mesh_0_30_io_out_a_0;
	wire [31:0] _mesh_0_30_io_out_c_0;
	wire [31:0] _mesh_0_30_io_out_b_0;
	wire _mesh_0_30_io_out_control_0_dataflow;
	wire _mesh_0_30_io_out_control_0_propagate;
	wire [4:0] _mesh_0_30_io_out_control_0_shift;
	wire [2:0] _mesh_0_30_io_out_id_0;
	wire _mesh_0_30_io_out_last_0;
	wire _mesh_0_30_io_out_valid_0;
	wire [31:0] _mesh_0_29_io_out_a_0;
	wire [31:0] _mesh_0_29_io_out_c_0;
	wire [31:0] _mesh_0_29_io_out_b_0;
	wire _mesh_0_29_io_out_control_0_dataflow;
	wire _mesh_0_29_io_out_control_0_propagate;
	wire [4:0] _mesh_0_29_io_out_control_0_shift;
	wire [2:0] _mesh_0_29_io_out_id_0;
	wire _mesh_0_29_io_out_last_0;
	wire _mesh_0_29_io_out_valid_0;
	wire [31:0] _mesh_0_28_io_out_a_0;
	wire [31:0] _mesh_0_28_io_out_c_0;
	wire [31:0] _mesh_0_28_io_out_b_0;
	wire _mesh_0_28_io_out_control_0_dataflow;
	wire _mesh_0_28_io_out_control_0_propagate;
	wire [4:0] _mesh_0_28_io_out_control_0_shift;
	wire [2:0] _mesh_0_28_io_out_id_0;
	wire _mesh_0_28_io_out_last_0;
	wire _mesh_0_28_io_out_valid_0;
	wire [31:0] _mesh_0_27_io_out_a_0;
	wire [31:0] _mesh_0_27_io_out_c_0;
	wire [31:0] _mesh_0_27_io_out_b_0;
	wire _mesh_0_27_io_out_control_0_dataflow;
	wire _mesh_0_27_io_out_control_0_propagate;
	wire [4:0] _mesh_0_27_io_out_control_0_shift;
	wire [2:0] _mesh_0_27_io_out_id_0;
	wire _mesh_0_27_io_out_last_0;
	wire _mesh_0_27_io_out_valid_0;
	wire [31:0] _mesh_0_26_io_out_a_0;
	wire [31:0] _mesh_0_26_io_out_c_0;
	wire [31:0] _mesh_0_26_io_out_b_0;
	wire _mesh_0_26_io_out_control_0_dataflow;
	wire _mesh_0_26_io_out_control_0_propagate;
	wire [4:0] _mesh_0_26_io_out_control_0_shift;
	wire [2:0] _mesh_0_26_io_out_id_0;
	wire _mesh_0_26_io_out_last_0;
	wire _mesh_0_26_io_out_valid_0;
	wire [31:0] _mesh_0_25_io_out_a_0;
	wire [31:0] _mesh_0_25_io_out_c_0;
	wire [31:0] _mesh_0_25_io_out_b_0;
	wire _mesh_0_25_io_out_control_0_dataflow;
	wire _mesh_0_25_io_out_control_0_propagate;
	wire [4:0] _mesh_0_25_io_out_control_0_shift;
	wire [2:0] _mesh_0_25_io_out_id_0;
	wire _mesh_0_25_io_out_last_0;
	wire _mesh_0_25_io_out_valid_0;
	wire [31:0] _mesh_0_24_io_out_a_0;
	wire [31:0] _mesh_0_24_io_out_c_0;
	wire [31:0] _mesh_0_24_io_out_b_0;
	wire _mesh_0_24_io_out_control_0_dataflow;
	wire _mesh_0_24_io_out_control_0_propagate;
	wire [4:0] _mesh_0_24_io_out_control_0_shift;
	wire [2:0] _mesh_0_24_io_out_id_0;
	wire _mesh_0_24_io_out_last_0;
	wire _mesh_0_24_io_out_valid_0;
	wire [31:0] _mesh_0_23_io_out_a_0;
	wire [31:0] _mesh_0_23_io_out_c_0;
	wire [31:0] _mesh_0_23_io_out_b_0;
	wire _mesh_0_23_io_out_control_0_dataflow;
	wire _mesh_0_23_io_out_control_0_propagate;
	wire [4:0] _mesh_0_23_io_out_control_0_shift;
	wire [2:0] _mesh_0_23_io_out_id_0;
	wire _mesh_0_23_io_out_last_0;
	wire _mesh_0_23_io_out_valid_0;
	wire [31:0] _mesh_0_22_io_out_a_0;
	wire [31:0] _mesh_0_22_io_out_c_0;
	wire [31:0] _mesh_0_22_io_out_b_0;
	wire _mesh_0_22_io_out_control_0_dataflow;
	wire _mesh_0_22_io_out_control_0_propagate;
	wire [4:0] _mesh_0_22_io_out_control_0_shift;
	wire [2:0] _mesh_0_22_io_out_id_0;
	wire _mesh_0_22_io_out_last_0;
	wire _mesh_0_22_io_out_valid_0;
	wire [31:0] _mesh_0_21_io_out_a_0;
	wire [31:0] _mesh_0_21_io_out_c_0;
	wire [31:0] _mesh_0_21_io_out_b_0;
	wire _mesh_0_21_io_out_control_0_dataflow;
	wire _mesh_0_21_io_out_control_0_propagate;
	wire [4:0] _mesh_0_21_io_out_control_0_shift;
	wire [2:0] _mesh_0_21_io_out_id_0;
	wire _mesh_0_21_io_out_last_0;
	wire _mesh_0_21_io_out_valid_0;
	wire [31:0] _mesh_0_20_io_out_a_0;
	wire [31:0] _mesh_0_20_io_out_c_0;
	wire [31:0] _mesh_0_20_io_out_b_0;
	wire _mesh_0_20_io_out_control_0_dataflow;
	wire _mesh_0_20_io_out_control_0_propagate;
	wire [4:0] _mesh_0_20_io_out_control_0_shift;
	wire [2:0] _mesh_0_20_io_out_id_0;
	wire _mesh_0_20_io_out_last_0;
	wire _mesh_0_20_io_out_valid_0;
	wire [31:0] _mesh_0_19_io_out_a_0;
	wire [31:0] _mesh_0_19_io_out_c_0;
	wire [31:0] _mesh_0_19_io_out_b_0;
	wire _mesh_0_19_io_out_control_0_dataflow;
	wire _mesh_0_19_io_out_control_0_propagate;
	wire [4:0] _mesh_0_19_io_out_control_0_shift;
	wire [2:0] _mesh_0_19_io_out_id_0;
	wire _mesh_0_19_io_out_last_0;
	wire _mesh_0_19_io_out_valid_0;
	wire [31:0] _mesh_0_18_io_out_a_0;
	wire [31:0] _mesh_0_18_io_out_c_0;
	wire [31:0] _mesh_0_18_io_out_b_0;
	wire _mesh_0_18_io_out_control_0_dataflow;
	wire _mesh_0_18_io_out_control_0_propagate;
	wire [4:0] _mesh_0_18_io_out_control_0_shift;
	wire [2:0] _mesh_0_18_io_out_id_0;
	wire _mesh_0_18_io_out_last_0;
	wire _mesh_0_18_io_out_valid_0;
	wire [31:0] _mesh_0_17_io_out_a_0;
	wire [31:0] _mesh_0_17_io_out_c_0;
	wire [31:0] _mesh_0_17_io_out_b_0;
	wire _mesh_0_17_io_out_control_0_dataflow;
	wire _mesh_0_17_io_out_control_0_propagate;
	wire [4:0] _mesh_0_17_io_out_control_0_shift;
	wire [2:0] _mesh_0_17_io_out_id_0;
	wire _mesh_0_17_io_out_last_0;
	wire _mesh_0_17_io_out_valid_0;
	wire [31:0] _mesh_0_16_io_out_a_0;
	wire [31:0] _mesh_0_16_io_out_c_0;
	wire [31:0] _mesh_0_16_io_out_b_0;
	wire _mesh_0_16_io_out_control_0_dataflow;
	wire _mesh_0_16_io_out_control_0_propagate;
	wire [4:0] _mesh_0_16_io_out_control_0_shift;
	wire [2:0] _mesh_0_16_io_out_id_0;
	wire _mesh_0_16_io_out_last_0;
	wire _mesh_0_16_io_out_valid_0;
	wire [31:0] _mesh_0_15_io_out_a_0;
	wire [31:0] _mesh_0_15_io_out_c_0;
	wire [31:0] _mesh_0_15_io_out_b_0;
	wire _mesh_0_15_io_out_control_0_dataflow;
	wire _mesh_0_15_io_out_control_0_propagate;
	wire [4:0] _mesh_0_15_io_out_control_0_shift;
	wire [2:0] _mesh_0_15_io_out_id_0;
	wire _mesh_0_15_io_out_last_0;
	wire _mesh_0_15_io_out_valid_0;
	wire [31:0] _mesh_0_14_io_out_a_0;
	wire [31:0] _mesh_0_14_io_out_c_0;
	wire [31:0] _mesh_0_14_io_out_b_0;
	wire _mesh_0_14_io_out_control_0_dataflow;
	wire _mesh_0_14_io_out_control_0_propagate;
	wire [4:0] _mesh_0_14_io_out_control_0_shift;
	wire [2:0] _mesh_0_14_io_out_id_0;
	wire _mesh_0_14_io_out_last_0;
	wire _mesh_0_14_io_out_valid_0;
	wire [31:0] _mesh_0_13_io_out_a_0;
	wire [31:0] _mesh_0_13_io_out_c_0;
	wire [31:0] _mesh_0_13_io_out_b_0;
	wire _mesh_0_13_io_out_control_0_dataflow;
	wire _mesh_0_13_io_out_control_0_propagate;
	wire [4:0] _mesh_0_13_io_out_control_0_shift;
	wire [2:0] _mesh_0_13_io_out_id_0;
	wire _mesh_0_13_io_out_last_0;
	wire _mesh_0_13_io_out_valid_0;
	wire [31:0] _mesh_0_12_io_out_a_0;
	wire [31:0] _mesh_0_12_io_out_c_0;
	wire [31:0] _mesh_0_12_io_out_b_0;
	wire _mesh_0_12_io_out_control_0_dataflow;
	wire _mesh_0_12_io_out_control_0_propagate;
	wire [4:0] _mesh_0_12_io_out_control_0_shift;
	wire [2:0] _mesh_0_12_io_out_id_0;
	wire _mesh_0_12_io_out_last_0;
	wire _mesh_0_12_io_out_valid_0;
	wire [31:0] _mesh_0_11_io_out_a_0;
	wire [31:0] _mesh_0_11_io_out_c_0;
	wire [31:0] _mesh_0_11_io_out_b_0;
	wire _mesh_0_11_io_out_control_0_dataflow;
	wire _mesh_0_11_io_out_control_0_propagate;
	wire [4:0] _mesh_0_11_io_out_control_0_shift;
	wire [2:0] _mesh_0_11_io_out_id_0;
	wire _mesh_0_11_io_out_last_0;
	wire _mesh_0_11_io_out_valid_0;
	wire [31:0] _mesh_0_10_io_out_a_0;
	wire [31:0] _mesh_0_10_io_out_c_0;
	wire [31:0] _mesh_0_10_io_out_b_0;
	wire _mesh_0_10_io_out_control_0_dataflow;
	wire _mesh_0_10_io_out_control_0_propagate;
	wire [4:0] _mesh_0_10_io_out_control_0_shift;
	wire [2:0] _mesh_0_10_io_out_id_0;
	wire _mesh_0_10_io_out_last_0;
	wire _mesh_0_10_io_out_valid_0;
	wire [31:0] _mesh_0_9_io_out_a_0;
	wire [31:0] _mesh_0_9_io_out_c_0;
	wire [31:0] _mesh_0_9_io_out_b_0;
	wire _mesh_0_9_io_out_control_0_dataflow;
	wire _mesh_0_9_io_out_control_0_propagate;
	wire [4:0] _mesh_0_9_io_out_control_0_shift;
	wire [2:0] _mesh_0_9_io_out_id_0;
	wire _mesh_0_9_io_out_last_0;
	wire _mesh_0_9_io_out_valid_0;
	wire [31:0] _mesh_0_8_io_out_a_0;
	wire [31:0] _mesh_0_8_io_out_c_0;
	wire [31:0] _mesh_0_8_io_out_b_0;
	wire _mesh_0_8_io_out_control_0_dataflow;
	wire _mesh_0_8_io_out_control_0_propagate;
	wire [4:0] _mesh_0_8_io_out_control_0_shift;
	wire [2:0] _mesh_0_8_io_out_id_0;
	wire _mesh_0_8_io_out_last_0;
	wire _mesh_0_8_io_out_valid_0;
	wire [31:0] _mesh_0_7_io_out_a_0;
	wire [31:0] _mesh_0_7_io_out_c_0;
	wire [31:0] _mesh_0_7_io_out_b_0;
	wire _mesh_0_7_io_out_control_0_dataflow;
	wire _mesh_0_7_io_out_control_0_propagate;
	wire [4:0] _mesh_0_7_io_out_control_0_shift;
	wire [2:0] _mesh_0_7_io_out_id_0;
	wire _mesh_0_7_io_out_last_0;
	wire _mesh_0_7_io_out_valid_0;
	wire [31:0] _mesh_0_6_io_out_a_0;
	wire [31:0] _mesh_0_6_io_out_c_0;
	wire [31:0] _mesh_0_6_io_out_b_0;
	wire _mesh_0_6_io_out_control_0_dataflow;
	wire _mesh_0_6_io_out_control_0_propagate;
	wire [4:0] _mesh_0_6_io_out_control_0_shift;
	wire [2:0] _mesh_0_6_io_out_id_0;
	wire _mesh_0_6_io_out_last_0;
	wire _mesh_0_6_io_out_valid_0;
	wire [31:0] _mesh_0_5_io_out_a_0;
	wire [31:0] _mesh_0_5_io_out_c_0;
	wire [31:0] _mesh_0_5_io_out_b_0;
	wire _mesh_0_5_io_out_control_0_dataflow;
	wire _mesh_0_5_io_out_control_0_propagate;
	wire [4:0] _mesh_0_5_io_out_control_0_shift;
	wire [2:0] _mesh_0_5_io_out_id_0;
	wire _mesh_0_5_io_out_last_0;
	wire _mesh_0_5_io_out_valid_0;
	wire [31:0] _mesh_0_4_io_out_a_0;
	wire [31:0] _mesh_0_4_io_out_c_0;
	wire [31:0] _mesh_0_4_io_out_b_0;
	wire _mesh_0_4_io_out_control_0_dataflow;
	wire _mesh_0_4_io_out_control_0_propagate;
	wire [4:0] _mesh_0_4_io_out_control_0_shift;
	wire [2:0] _mesh_0_4_io_out_id_0;
	wire _mesh_0_4_io_out_last_0;
	wire _mesh_0_4_io_out_valid_0;
	wire [31:0] _mesh_0_3_io_out_a_0;
	wire [31:0] _mesh_0_3_io_out_c_0;
	wire [31:0] _mesh_0_3_io_out_b_0;
	wire _mesh_0_3_io_out_control_0_dataflow;
	wire _mesh_0_3_io_out_control_0_propagate;
	wire [4:0] _mesh_0_3_io_out_control_0_shift;
	wire [2:0] _mesh_0_3_io_out_id_0;
	wire _mesh_0_3_io_out_last_0;
	wire _mesh_0_3_io_out_valid_0;
	wire [31:0] _mesh_0_2_io_out_a_0;
	wire [31:0] _mesh_0_2_io_out_c_0;
	wire [31:0] _mesh_0_2_io_out_b_0;
	wire _mesh_0_2_io_out_control_0_dataflow;
	wire _mesh_0_2_io_out_control_0_propagate;
	wire [4:0] _mesh_0_2_io_out_control_0_shift;
	wire [2:0] _mesh_0_2_io_out_id_0;
	wire _mesh_0_2_io_out_last_0;
	wire _mesh_0_2_io_out_valid_0;
	wire [31:0] _mesh_0_1_io_out_a_0;
	wire [31:0] _mesh_0_1_io_out_c_0;
	wire [31:0] _mesh_0_1_io_out_b_0;
	wire _mesh_0_1_io_out_control_0_dataflow;
	wire _mesh_0_1_io_out_control_0_propagate;
	wire [4:0] _mesh_0_1_io_out_control_0_shift;
	wire [2:0] _mesh_0_1_io_out_id_0;
	wire _mesh_0_1_io_out_last_0;
	wire _mesh_0_1_io_out_valid_0;
	wire [31:0] _mesh_0_0_io_out_a_0;
	wire [31:0] _mesh_0_0_io_out_c_0;
	wire [31:0] _mesh_0_0_io_out_b_0;
	wire _mesh_0_0_io_out_control_0_dataflow;
	wire _mesh_0_0_io_out_control_0_propagate;
	wire [4:0] _mesh_0_0_io_out_control_0_shift;
	wire [2:0] _mesh_0_0_io_out_id_0;
	wire _mesh_0_0_io_out_last_0;
	wire _mesh_0_0_io_out_valid_0;
	reg [31:0] r_0;
	reg [31:0] r_1_0;
	reg [31:0] r_2_0;
	reg [31:0] r_3_0;
	reg [31:0] r_4_0;
	reg [31:0] r_5_0;
	reg [31:0] r_6_0;
	reg [31:0] r_7_0;
	reg [31:0] r_8_0;
	reg [31:0] r_9_0;
	reg [31:0] r_10_0;
	reg [31:0] r_11_0;
	reg [31:0] r_12_0;
	reg [31:0] r_13_0;
	reg [31:0] r_14_0;
	reg [31:0] r_15_0;
	reg [31:0] r_16_0;
	reg [31:0] r_17_0;
	reg [31:0] r_18_0;
	reg [31:0] r_19_0;
	reg [31:0] r_20_0;
	reg [31:0] r_21_0;
	reg [31:0] r_22_0;
	reg [31:0] r_23_0;
	reg [31:0] r_24_0;
	reg [31:0] r_25_0;
	reg [31:0] r_26_0;
	reg [31:0] r_27_0;
	reg [31:0] r_28_0;
	reg [31:0] r_29_0;
	reg [31:0] r_30_0;
	reg [31:0] r_31_0;
	reg [31:0] r_32_0;
	reg [31:0] r_33_0;
	reg [31:0] r_34_0;
	reg [31:0] r_35_0;
	reg [31:0] r_36_0;
	reg [31:0] r_37_0;
	reg [31:0] r_38_0;
	reg [31:0] r_39_0;
	reg [31:0] r_40_0;
	reg [31:0] r_41_0;
	reg [31:0] r_42_0;
	reg [31:0] r_43_0;
	reg [31:0] r_44_0;
	reg [31:0] r_45_0;
	reg [31:0] r_46_0;
	reg [31:0] r_47_0;
	reg [31:0] r_48_0;
	reg [31:0] r_49_0;
	reg [31:0] r_50_0;
	reg [31:0] r_51_0;
	reg [31:0] r_52_0;
	reg [31:0] r_53_0;
	reg [31:0] r_54_0;
	reg [31:0] r_55_0;
	reg [31:0] r_56_0;
	reg [31:0] r_57_0;
	reg [31:0] r_58_0;
	reg [31:0] r_59_0;
	reg [31:0] r_60_0;
	reg [31:0] r_61_0;
	reg [31:0] r_62_0;
	reg [31:0] r_63_0;
	reg [31:0] r_64_0;
	reg [31:0] r_65_0;
	reg [31:0] r_66_0;
	reg [31:0] r_67_0;
	reg [31:0] r_68_0;
	reg [31:0] r_69_0;
	reg [31:0] r_70_0;
	reg [31:0] r_71_0;
	reg [31:0] r_72_0;
	reg [31:0] r_73_0;
	reg [31:0] r_74_0;
	reg [31:0] r_75_0;
	reg [31:0] r_76_0;
	reg [31:0] r_77_0;
	reg [31:0] r_78_0;
	reg [31:0] r_79_0;
	reg [31:0] r_80_0;
	reg [31:0] r_81_0;
	reg [31:0] r_82_0;
	reg [31:0] r_83_0;
	reg [31:0] r_84_0;
	reg [31:0] r_85_0;
	reg [31:0] r_86_0;
	reg [31:0] r_87_0;
	reg [31:0] r_88_0;
	reg [31:0] r_89_0;
	reg [31:0] r_90_0;
	reg [31:0] r_91_0;
	reg [31:0] r_92_0;
	reg [31:0] r_93_0;
	reg [31:0] r_94_0;
	reg [31:0] r_95_0;
	reg [31:0] r_96_0;
	reg [31:0] r_97_0;
	reg [31:0] r_98_0;
	reg [31:0] r_99_0;
	reg [31:0] r_100_0;
	reg [31:0] r_101_0;
	reg [31:0] r_102_0;
	reg [31:0] r_103_0;
	reg [31:0] r_104_0;
	reg [31:0] r_105_0;
	reg [31:0] r_106_0;
	reg [31:0] r_107_0;
	reg [31:0] r_108_0;
	reg [31:0] r_109_0;
	reg [31:0] r_110_0;
	reg [31:0] r_111_0;
	reg [31:0] r_112_0;
	reg [31:0] r_113_0;
	reg [31:0] r_114_0;
	reg [31:0] r_115_0;
	reg [31:0] r_116_0;
	reg [31:0] r_117_0;
	reg [31:0] r_118_0;
	reg [31:0] r_119_0;
	reg [31:0] r_120_0;
	reg [31:0] r_121_0;
	reg [31:0] r_122_0;
	reg [31:0] r_123_0;
	reg [31:0] r_124_0;
	reg [31:0] r_125_0;
	reg [31:0] r_126_0;
	reg [31:0] r_127_0;
	reg [31:0] r_128_0;
	reg [31:0] r_129_0;
	reg [31:0] r_130_0;
	reg [31:0] r_131_0;
	reg [31:0] r_132_0;
	reg [31:0] r_133_0;
	reg [31:0] r_134_0;
	reg [31:0] r_135_0;
	reg [31:0] r_136_0;
	reg [31:0] r_137_0;
	reg [31:0] r_138_0;
	reg [31:0] r_139_0;
	reg [31:0] r_140_0;
	reg [31:0] r_141_0;
	reg [31:0] r_142_0;
	reg [31:0] r_143_0;
	reg [31:0] r_144_0;
	reg [31:0] r_145_0;
	reg [31:0] r_146_0;
	reg [31:0] r_147_0;
	reg [31:0] r_148_0;
	reg [31:0] r_149_0;
	reg [31:0] r_150_0;
	reg [31:0] r_151_0;
	reg [31:0] r_152_0;
	reg [31:0] r_153_0;
	reg [31:0] r_154_0;
	reg [31:0] r_155_0;
	reg [31:0] r_156_0;
	reg [31:0] r_157_0;
	reg [31:0] r_158_0;
	reg [31:0] r_159_0;
	reg [31:0] r_160_0;
	reg [31:0] r_161_0;
	reg [31:0] r_162_0;
	reg [31:0] r_163_0;
	reg [31:0] r_164_0;
	reg [31:0] r_165_0;
	reg [31:0] r_166_0;
	reg [31:0] r_167_0;
	reg [31:0] r_168_0;
	reg [31:0] r_169_0;
	reg [31:0] r_170_0;
	reg [31:0] r_171_0;
	reg [31:0] r_172_0;
	reg [31:0] r_173_0;
	reg [31:0] r_174_0;
	reg [31:0] r_175_0;
	reg [31:0] r_176_0;
	reg [31:0] r_177_0;
	reg [31:0] r_178_0;
	reg [31:0] r_179_0;
	reg [31:0] r_180_0;
	reg [31:0] r_181_0;
	reg [31:0] r_182_0;
	reg [31:0] r_183_0;
	reg [31:0] r_184_0;
	reg [31:0] r_185_0;
	reg [31:0] r_186_0;
	reg [31:0] r_187_0;
	reg [31:0] r_188_0;
	reg [31:0] r_189_0;
	reg [31:0] r_190_0;
	reg [31:0] r_191_0;
	reg [31:0] r_192_0;
	reg [31:0] r_193_0;
	reg [31:0] r_194_0;
	reg [31:0] r_195_0;
	reg [31:0] r_196_0;
	reg [31:0] r_197_0;
	reg [31:0] r_198_0;
	reg [31:0] r_199_0;
	reg [31:0] r_200_0;
	reg [31:0] r_201_0;
	reg [31:0] r_202_0;
	reg [31:0] r_203_0;
	reg [31:0] r_204_0;
	reg [31:0] r_205_0;
	reg [31:0] r_206_0;
	reg [31:0] r_207_0;
	reg [31:0] r_208_0;
	reg [31:0] r_209_0;
	reg [31:0] r_210_0;
	reg [31:0] r_211_0;
	reg [31:0] r_212_0;
	reg [31:0] r_213_0;
	reg [31:0] r_214_0;
	reg [31:0] r_215_0;
	reg [31:0] r_216_0;
	reg [31:0] r_217_0;
	reg [31:0] r_218_0;
	reg [31:0] r_219_0;
	reg [31:0] r_220_0;
	reg [31:0] r_221_0;
	reg [31:0] r_222_0;
	reg [31:0] r_223_0;
	reg [31:0] r_224_0;
	reg [31:0] r_225_0;
	reg [31:0] r_226_0;
	reg [31:0] r_227_0;
	reg [31:0] r_228_0;
	reg [31:0] r_229_0;
	reg [31:0] r_230_0;
	reg [31:0] r_231_0;
	reg [31:0] r_232_0;
	reg [31:0] r_233_0;
	reg [31:0] r_234_0;
	reg [31:0] r_235_0;
	reg [31:0] r_236_0;
	reg [31:0] r_237_0;
	reg [31:0] r_238_0;
	reg [31:0] r_239_0;
	reg [31:0] r_240_0;
	reg [31:0] r_241_0;
	reg [31:0] r_242_0;
	reg [31:0] r_243_0;
	reg [31:0] r_244_0;
	reg [31:0] r_245_0;
	reg [31:0] r_246_0;
	reg [31:0] r_247_0;
	reg [31:0] r_248_0;
	reg [31:0] r_249_0;
	reg [31:0] r_250_0;
	reg [31:0] r_251_0;
	reg [31:0] r_252_0;
	reg [31:0] r_253_0;
	reg [31:0] r_254_0;
	reg [31:0] r_255_0;
	reg [31:0] r_256_0;
	reg [31:0] r_257_0;
	reg [31:0] r_258_0;
	reg [31:0] r_259_0;
	reg [31:0] r_260_0;
	reg [31:0] r_261_0;
	reg [31:0] r_262_0;
	reg [31:0] r_263_0;
	reg [31:0] r_264_0;
	reg [31:0] r_265_0;
	reg [31:0] r_266_0;
	reg [31:0] r_267_0;
	reg [31:0] r_268_0;
	reg [31:0] r_269_0;
	reg [31:0] r_270_0;
	reg [31:0] r_271_0;
	reg [31:0] r_272_0;
	reg [31:0] r_273_0;
	reg [31:0] r_274_0;
	reg [31:0] r_275_0;
	reg [31:0] r_276_0;
	reg [31:0] r_277_0;
	reg [31:0] r_278_0;
	reg [31:0] r_279_0;
	reg [31:0] r_280_0;
	reg [31:0] r_281_0;
	reg [31:0] r_282_0;
	reg [31:0] r_283_0;
	reg [31:0] r_284_0;
	reg [31:0] r_285_0;
	reg [31:0] r_286_0;
	reg [31:0] r_287_0;
	reg [31:0] r_288_0;
	reg [31:0] r_289_0;
	reg [31:0] r_290_0;
	reg [31:0] r_291_0;
	reg [31:0] r_292_0;
	reg [31:0] r_293_0;
	reg [31:0] r_294_0;
	reg [31:0] r_295_0;
	reg [31:0] r_296_0;
	reg [31:0] r_297_0;
	reg [31:0] r_298_0;
	reg [31:0] r_299_0;
	reg [31:0] r_300_0;
	reg [31:0] r_301_0;
	reg [31:0] r_302_0;
	reg [31:0] r_303_0;
	reg [31:0] r_304_0;
	reg [31:0] r_305_0;
	reg [31:0] r_306_0;
	reg [31:0] r_307_0;
	reg [31:0] r_308_0;
	reg [31:0] r_309_0;
	reg [31:0] r_310_0;
	reg [31:0] r_311_0;
	reg [31:0] r_312_0;
	reg [31:0] r_313_0;
	reg [31:0] r_314_0;
	reg [31:0] r_315_0;
	reg [31:0] r_316_0;
	reg [31:0] r_317_0;
	reg [31:0] r_318_0;
	reg [31:0] r_319_0;
	reg [31:0] r_320_0;
	reg [31:0] r_321_0;
	reg [31:0] r_322_0;
	reg [31:0] r_323_0;
	reg [31:0] r_324_0;
	reg [31:0] r_325_0;
	reg [31:0] r_326_0;
	reg [31:0] r_327_0;
	reg [31:0] r_328_0;
	reg [31:0] r_329_0;
	reg [31:0] r_330_0;
	reg [31:0] r_331_0;
	reg [31:0] r_332_0;
	reg [31:0] r_333_0;
	reg [31:0] r_334_0;
	reg [31:0] r_335_0;
	reg [31:0] r_336_0;
	reg [31:0] r_337_0;
	reg [31:0] r_338_0;
	reg [31:0] r_339_0;
	reg [31:0] r_340_0;
	reg [31:0] r_341_0;
	reg [31:0] r_342_0;
	reg [31:0] r_343_0;
	reg [31:0] r_344_0;
	reg [31:0] r_345_0;
	reg [31:0] r_346_0;
	reg [31:0] r_347_0;
	reg [31:0] r_348_0;
	reg [31:0] r_349_0;
	reg [31:0] r_350_0;
	reg [31:0] r_351_0;
	reg [31:0] r_352_0;
	reg [31:0] r_353_0;
	reg [31:0] r_354_0;
	reg [31:0] r_355_0;
	reg [31:0] r_356_0;
	reg [31:0] r_357_0;
	reg [31:0] r_358_0;
	reg [31:0] r_359_0;
	reg [31:0] r_360_0;
	reg [31:0] r_361_0;
	reg [31:0] r_362_0;
	reg [31:0] r_363_0;
	reg [31:0] r_364_0;
	reg [31:0] r_365_0;
	reg [31:0] r_366_0;
	reg [31:0] r_367_0;
	reg [31:0] r_368_0;
	reg [31:0] r_369_0;
	reg [31:0] r_370_0;
	reg [31:0] r_371_0;
	reg [31:0] r_372_0;
	reg [31:0] r_373_0;
	reg [31:0] r_374_0;
	reg [31:0] r_375_0;
	reg [31:0] r_376_0;
	reg [31:0] r_377_0;
	reg [31:0] r_378_0;
	reg [31:0] r_379_0;
	reg [31:0] r_380_0;
	reg [31:0] r_381_0;
	reg [31:0] r_382_0;
	reg [31:0] r_383_0;
	reg [31:0] r_384_0;
	reg [31:0] r_385_0;
	reg [31:0] r_386_0;
	reg [31:0] r_387_0;
	reg [31:0] r_388_0;
	reg [31:0] r_389_0;
	reg [31:0] r_390_0;
	reg [31:0] r_391_0;
	reg [31:0] r_392_0;
	reg [31:0] r_393_0;
	reg [31:0] r_394_0;
	reg [31:0] r_395_0;
	reg [31:0] r_396_0;
	reg [31:0] r_397_0;
	reg [31:0] r_398_0;
	reg [31:0] r_399_0;
	reg [31:0] r_400_0;
	reg [31:0] r_401_0;
	reg [31:0] r_402_0;
	reg [31:0] r_403_0;
	reg [31:0] r_404_0;
	reg [31:0] r_405_0;
	reg [31:0] r_406_0;
	reg [31:0] r_407_0;
	reg [31:0] r_408_0;
	reg [31:0] r_409_0;
	reg [31:0] r_410_0;
	reg [31:0] r_411_0;
	reg [31:0] r_412_0;
	reg [31:0] r_413_0;
	reg [31:0] r_414_0;
	reg [31:0] r_415_0;
	reg [31:0] r_416_0;
	reg [31:0] r_417_0;
	reg [31:0] r_418_0;
	reg [31:0] r_419_0;
	reg [31:0] r_420_0;
	reg [31:0] r_421_0;
	reg [31:0] r_422_0;
	reg [31:0] r_423_0;
	reg [31:0] r_424_0;
	reg [31:0] r_425_0;
	reg [31:0] r_426_0;
	reg [31:0] r_427_0;
	reg [31:0] r_428_0;
	reg [31:0] r_429_0;
	reg [31:0] r_430_0;
	reg [31:0] r_431_0;
	reg [31:0] r_432_0;
	reg [31:0] r_433_0;
	reg [31:0] r_434_0;
	reg [31:0] r_435_0;
	reg [31:0] r_436_0;
	reg [31:0] r_437_0;
	reg [31:0] r_438_0;
	reg [31:0] r_439_0;
	reg [31:0] r_440_0;
	reg [31:0] r_441_0;
	reg [31:0] r_442_0;
	reg [31:0] r_443_0;
	reg [31:0] r_444_0;
	reg [31:0] r_445_0;
	reg [31:0] r_446_0;
	reg [31:0] r_447_0;
	reg [31:0] r_448_0;
	reg [31:0] r_449_0;
	reg [31:0] r_450_0;
	reg [31:0] r_451_0;
	reg [31:0] r_452_0;
	reg [31:0] r_453_0;
	reg [31:0] r_454_0;
	reg [31:0] r_455_0;
	reg [31:0] r_456_0;
	reg [31:0] r_457_0;
	reg [31:0] r_458_0;
	reg [31:0] r_459_0;
	reg [31:0] r_460_0;
	reg [31:0] r_461_0;
	reg [31:0] r_462_0;
	reg [31:0] r_463_0;
	reg [31:0] r_464_0;
	reg [31:0] r_465_0;
	reg [31:0] r_466_0;
	reg [31:0] r_467_0;
	reg [31:0] r_468_0;
	reg [31:0] r_469_0;
	reg [31:0] r_470_0;
	reg [31:0] r_471_0;
	reg [31:0] r_472_0;
	reg [31:0] r_473_0;
	reg [31:0] r_474_0;
	reg [31:0] r_475_0;
	reg [31:0] r_476_0;
	reg [31:0] r_477_0;
	reg [31:0] r_478_0;
	reg [31:0] r_479_0;
	reg [31:0] r_480_0;
	reg [31:0] r_481_0;
	reg [31:0] r_482_0;
	reg [31:0] r_483_0;
	reg [31:0] r_484_0;
	reg [31:0] r_485_0;
	reg [31:0] r_486_0;
	reg [31:0] r_487_0;
	reg [31:0] r_488_0;
	reg [31:0] r_489_0;
	reg [31:0] r_490_0;
	reg [31:0] r_491_0;
	reg [31:0] r_492_0;
	reg [31:0] r_493_0;
	reg [31:0] r_494_0;
	reg [31:0] r_495_0;
	reg [31:0] r_496_0;
	reg [31:0] r_497_0;
	reg [31:0] r_498_0;
	reg [31:0] r_499_0;
	reg [31:0] r_500_0;
	reg [31:0] r_501_0;
	reg [31:0] r_502_0;
	reg [31:0] r_503_0;
	reg [31:0] r_504_0;
	reg [31:0] r_505_0;
	reg [31:0] r_506_0;
	reg [31:0] r_507_0;
	reg [31:0] r_508_0;
	reg [31:0] r_509_0;
	reg [31:0] r_510_0;
	reg [31:0] r_511_0;
	reg [31:0] r_512_0;
	reg [31:0] r_513_0;
	reg [31:0] r_514_0;
	reg [31:0] r_515_0;
	reg [31:0] r_516_0;
	reg [31:0] r_517_0;
	reg [31:0] r_518_0;
	reg [31:0] r_519_0;
	reg [31:0] r_520_0;
	reg [31:0] r_521_0;
	reg [31:0] r_522_0;
	reg [31:0] r_523_0;
	reg [31:0] r_524_0;
	reg [31:0] r_525_0;
	reg [31:0] r_526_0;
	reg [31:0] r_527_0;
	reg [31:0] r_528_0;
	reg [31:0] r_529_0;
	reg [31:0] r_530_0;
	reg [31:0] r_531_0;
	reg [31:0] r_532_0;
	reg [31:0] r_533_0;
	reg [31:0] r_534_0;
	reg [31:0] r_535_0;
	reg [31:0] r_536_0;
	reg [31:0] r_537_0;
	reg [31:0] r_538_0;
	reg [31:0] r_539_0;
	reg [31:0] r_540_0;
	reg [31:0] r_541_0;
	reg [31:0] r_542_0;
	reg [31:0] r_543_0;
	reg [31:0] r_544_0;
	reg [31:0] r_545_0;
	reg [31:0] r_546_0;
	reg [31:0] r_547_0;
	reg [31:0] r_548_0;
	reg [31:0] r_549_0;
	reg [31:0] r_550_0;
	reg [31:0] r_551_0;
	reg [31:0] r_552_0;
	reg [31:0] r_553_0;
	reg [31:0] r_554_0;
	reg [31:0] r_555_0;
	reg [31:0] r_556_0;
	reg [31:0] r_557_0;
	reg [31:0] r_558_0;
	reg [31:0] r_559_0;
	reg [31:0] r_560_0;
	reg [31:0] r_561_0;
	reg [31:0] r_562_0;
	reg [31:0] r_563_0;
	reg [31:0] r_564_0;
	reg [31:0] r_565_0;
	reg [31:0] r_566_0;
	reg [31:0] r_567_0;
	reg [31:0] r_568_0;
	reg [31:0] r_569_0;
	reg [31:0] r_570_0;
	reg [31:0] r_571_0;
	reg [31:0] r_572_0;
	reg [31:0] r_573_0;
	reg [31:0] r_574_0;
	reg [31:0] r_575_0;
	reg [31:0] r_576_0;
	reg [31:0] r_577_0;
	reg [31:0] r_578_0;
	reg [31:0] r_579_0;
	reg [31:0] r_580_0;
	reg [31:0] r_581_0;
	reg [31:0] r_582_0;
	reg [31:0] r_583_0;
	reg [31:0] r_584_0;
	reg [31:0] r_585_0;
	reg [31:0] r_586_0;
	reg [31:0] r_587_0;
	reg [31:0] r_588_0;
	reg [31:0] r_589_0;
	reg [31:0] r_590_0;
	reg [31:0] r_591_0;
	reg [31:0] r_592_0;
	reg [31:0] r_593_0;
	reg [31:0] r_594_0;
	reg [31:0] r_595_0;
	reg [31:0] r_596_0;
	reg [31:0] r_597_0;
	reg [31:0] r_598_0;
	reg [31:0] r_599_0;
	reg [31:0] r_600_0;
	reg [31:0] r_601_0;
	reg [31:0] r_602_0;
	reg [31:0] r_603_0;
	reg [31:0] r_604_0;
	reg [31:0] r_605_0;
	reg [31:0] r_606_0;
	reg [31:0] r_607_0;
	reg [31:0] r_608_0;
	reg [31:0] r_609_0;
	reg [31:0] r_610_0;
	reg [31:0] r_611_0;
	reg [31:0] r_612_0;
	reg [31:0] r_613_0;
	reg [31:0] r_614_0;
	reg [31:0] r_615_0;
	reg [31:0] r_616_0;
	reg [31:0] r_617_0;
	reg [31:0] r_618_0;
	reg [31:0] r_619_0;
	reg [31:0] r_620_0;
	reg [31:0] r_621_0;
	reg [31:0] r_622_0;
	reg [31:0] r_623_0;
	reg [31:0] r_624_0;
	reg [31:0] r_625_0;
	reg [31:0] r_626_0;
	reg [31:0] r_627_0;
	reg [31:0] r_628_0;
	reg [31:0] r_629_0;
	reg [31:0] r_630_0;
	reg [31:0] r_631_0;
	reg [31:0] r_632_0;
	reg [31:0] r_633_0;
	reg [31:0] r_634_0;
	reg [31:0] r_635_0;
	reg [31:0] r_636_0;
	reg [31:0] r_637_0;
	reg [31:0] r_638_0;
	reg [31:0] r_639_0;
	reg [31:0] r_640_0;
	reg [31:0] r_641_0;
	reg [31:0] r_642_0;
	reg [31:0] r_643_0;
	reg [31:0] r_644_0;
	reg [31:0] r_645_0;
	reg [31:0] r_646_0;
	reg [31:0] r_647_0;
	reg [31:0] r_648_0;
	reg [31:0] r_649_0;
	reg [31:0] r_650_0;
	reg [31:0] r_651_0;
	reg [31:0] r_652_0;
	reg [31:0] r_653_0;
	reg [31:0] r_654_0;
	reg [31:0] r_655_0;
	reg [31:0] r_656_0;
	reg [31:0] r_657_0;
	reg [31:0] r_658_0;
	reg [31:0] r_659_0;
	reg [31:0] r_660_0;
	reg [31:0] r_661_0;
	reg [31:0] r_662_0;
	reg [31:0] r_663_0;
	reg [31:0] r_664_0;
	reg [31:0] r_665_0;
	reg [31:0] r_666_0;
	reg [31:0] r_667_0;
	reg [31:0] r_668_0;
	reg [31:0] r_669_0;
	reg [31:0] r_670_0;
	reg [31:0] r_671_0;
	reg [31:0] r_672_0;
	reg [31:0] r_673_0;
	reg [31:0] r_674_0;
	reg [31:0] r_675_0;
	reg [31:0] r_676_0;
	reg [31:0] r_677_0;
	reg [31:0] r_678_0;
	reg [31:0] r_679_0;
	reg [31:0] r_680_0;
	reg [31:0] r_681_0;
	reg [31:0] r_682_0;
	reg [31:0] r_683_0;
	reg [31:0] r_684_0;
	reg [31:0] r_685_0;
	reg [31:0] r_686_0;
	reg [31:0] r_687_0;
	reg [31:0] r_688_0;
	reg [31:0] r_689_0;
	reg [31:0] r_690_0;
	reg [31:0] r_691_0;
	reg [31:0] r_692_0;
	reg [31:0] r_693_0;
	reg [31:0] r_694_0;
	reg [31:0] r_695_0;
	reg [31:0] r_696_0;
	reg [31:0] r_697_0;
	reg [31:0] r_698_0;
	reg [31:0] r_699_0;
	reg [31:0] r_700_0;
	reg [31:0] r_701_0;
	reg [31:0] r_702_0;
	reg [31:0] r_703_0;
	reg [31:0] r_704_0;
	reg [31:0] r_705_0;
	reg [31:0] r_706_0;
	reg [31:0] r_707_0;
	reg [31:0] r_708_0;
	reg [31:0] r_709_0;
	reg [31:0] r_710_0;
	reg [31:0] r_711_0;
	reg [31:0] r_712_0;
	reg [31:0] r_713_0;
	reg [31:0] r_714_0;
	reg [31:0] r_715_0;
	reg [31:0] r_716_0;
	reg [31:0] r_717_0;
	reg [31:0] r_718_0;
	reg [31:0] r_719_0;
	reg [31:0] r_720_0;
	reg [31:0] r_721_0;
	reg [31:0] r_722_0;
	reg [31:0] r_723_0;
	reg [31:0] r_724_0;
	reg [31:0] r_725_0;
	reg [31:0] r_726_0;
	reg [31:0] r_727_0;
	reg [31:0] r_728_0;
	reg [31:0] r_729_0;
	reg [31:0] r_730_0;
	reg [31:0] r_731_0;
	reg [31:0] r_732_0;
	reg [31:0] r_733_0;
	reg [31:0] r_734_0;
	reg [31:0] r_735_0;
	reg [31:0] r_736_0;
	reg [31:0] r_737_0;
	reg [31:0] r_738_0;
	reg [31:0] r_739_0;
	reg [31:0] r_740_0;
	reg [31:0] r_741_0;
	reg [31:0] r_742_0;
	reg [31:0] r_743_0;
	reg [31:0] r_744_0;
	reg [31:0] r_745_0;
	reg [31:0] r_746_0;
	reg [31:0] r_747_0;
	reg [31:0] r_748_0;
	reg [31:0] r_749_0;
	reg [31:0] r_750_0;
	reg [31:0] r_751_0;
	reg [31:0] r_752_0;
	reg [31:0] r_753_0;
	reg [31:0] r_754_0;
	reg [31:0] r_755_0;
	reg [31:0] r_756_0;
	reg [31:0] r_757_0;
	reg [31:0] r_758_0;
	reg [31:0] r_759_0;
	reg [31:0] r_760_0;
	reg [31:0] r_761_0;
	reg [31:0] r_762_0;
	reg [31:0] r_763_0;
	reg [31:0] r_764_0;
	reg [31:0] r_765_0;
	reg [31:0] r_766_0;
	reg [31:0] r_767_0;
	reg [31:0] r_768_0;
	reg [31:0] r_769_0;
	reg [31:0] r_770_0;
	reg [31:0] r_771_0;
	reg [31:0] r_772_0;
	reg [31:0] r_773_0;
	reg [31:0] r_774_0;
	reg [31:0] r_775_0;
	reg [31:0] r_776_0;
	reg [31:0] r_777_0;
	reg [31:0] r_778_0;
	reg [31:0] r_779_0;
	reg [31:0] r_780_0;
	reg [31:0] r_781_0;
	reg [31:0] r_782_0;
	reg [31:0] r_783_0;
	reg [31:0] r_784_0;
	reg [31:0] r_785_0;
	reg [31:0] r_786_0;
	reg [31:0] r_787_0;
	reg [31:0] r_788_0;
	reg [31:0] r_789_0;
	reg [31:0] r_790_0;
	reg [31:0] r_791_0;
	reg [31:0] r_792_0;
	reg [31:0] r_793_0;
	reg [31:0] r_794_0;
	reg [31:0] r_795_0;
	reg [31:0] r_796_0;
	reg [31:0] r_797_0;
	reg [31:0] r_798_0;
	reg [31:0] r_799_0;
	reg [31:0] r_800_0;
	reg [31:0] r_801_0;
	reg [31:0] r_802_0;
	reg [31:0] r_803_0;
	reg [31:0] r_804_0;
	reg [31:0] r_805_0;
	reg [31:0] r_806_0;
	reg [31:0] r_807_0;
	reg [31:0] r_808_0;
	reg [31:0] r_809_0;
	reg [31:0] r_810_0;
	reg [31:0] r_811_0;
	reg [31:0] r_812_0;
	reg [31:0] r_813_0;
	reg [31:0] r_814_0;
	reg [31:0] r_815_0;
	reg [31:0] r_816_0;
	reg [31:0] r_817_0;
	reg [31:0] r_818_0;
	reg [31:0] r_819_0;
	reg [31:0] r_820_0;
	reg [31:0] r_821_0;
	reg [31:0] r_822_0;
	reg [31:0] r_823_0;
	reg [31:0] r_824_0;
	reg [31:0] r_825_0;
	reg [31:0] r_826_0;
	reg [31:0] r_827_0;
	reg [31:0] r_828_0;
	reg [31:0] r_829_0;
	reg [31:0] r_830_0;
	reg [31:0] r_831_0;
	reg [31:0] r_832_0;
	reg [31:0] r_833_0;
	reg [31:0] r_834_0;
	reg [31:0] r_835_0;
	reg [31:0] r_836_0;
	reg [31:0] r_837_0;
	reg [31:0] r_838_0;
	reg [31:0] r_839_0;
	reg [31:0] r_840_0;
	reg [31:0] r_841_0;
	reg [31:0] r_842_0;
	reg [31:0] r_843_0;
	reg [31:0] r_844_0;
	reg [31:0] r_845_0;
	reg [31:0] r_846_0;
	reg [31:0] r_847_0;
	reg [31:0] r_848_0;
	reg [31:0] r_849_0;
	reg [31:0] r_850_0;
	reg [31:0] r_851_0;
	reg [31:0] r_852_0;
	reg [31:0] r_853_0;
	reg [31:0] r_854_0;
	reg [31:0] r_855_0;
	reg [31:0] r_856_0;
	reg [31:0] r_857_0;
	reg [31:0] r_858_0;
	reg [31:0] r_859_0;
	reg [31:0] r_860_0;
	reg [31:0] r_861_0;
	reg [31:0] r_862_0;
	reg [31:0] r_863_0;
	reg [31:0] r_864_0;
	reg [31:0] r_865_0;
	reg [31:0] r_866_0;
	reg [31:0] r_867_0;
	reg [31:0] r_868_0;
	reg [31:0] r_869_0;
	reg [31:0] r_870_0;
	reg [31:0] r_871_0;
	reg [31:0] r_872_0;
	reg [31:0] r_873_0;
	reg [31:0] r_874_0;
	reg [31:0] r_875_0;
	reg [31:0] r_876_0;
	reg [31:0] r_877_0;
	reg [31:0] r_878_0;
	reg [31:0] r_879_0;
	reg [31:0] r_880_0;
	reg [31:0] r_881_0;
	reg [31:0] r_882_0;
	reg [31:0] r_883_0;
	reg [31:0] r_884_0;
	reg [31:0] r_885_0;
	reg [31:0] r_886_0;
	reg [31:0] r_887_0;
	reg [31:0] r_888_0;
	reg [31:0] r_889_0;
	reg [31:0] r_890_0;
	reg [31:0] r_891_0;
	reg [31:0] r_892_0;
	reg [31:0] r_893_0;
	reg [31:0] r_894_0;
	reg [31:0] r_895_0;
	reg [31:0] r_896_0;
	reg [31:0] r_897_0;
	reg [31:0] r_898_0;
	reg [31:0] r_899_0;
	reg [31:0] r_900_0;
	reg [31:0] r_901_0;
	reg [31:0] r_902_0;
	reg [31:0] r_903_0;
	reg [31:0] r_904_0;
	reg [31:0] r_905_0;
	reg [31:0] r_906_0;
	reg [31:0] r_907_0;
	reg [31:0] r_908_0;
	reg [31:0] r_909_0;
	reg [31:0] r_910_0;
	reg [31:0] r_911_0;
	reg [31:0] r_912_0;
	reg [31:0] r_913_0;
	reg [31:0] r_914_0;
	reg [31:0] r_915_0;
	reg [31:0] r_916_0;
	reg [31:0] r_917_0;
	reg [31:0] r_918_0;
	reg [31:0] r_919_0;
	reg [31:0] r_920_0;
	reg [31:0] r_921_0;
	reg [31:0] r_922_0;
	reg [31:0] r_923_0;
	reg [31:0] r_924_0;
	reg [31:0] r_925_0;
	reg [31:0] r_926_0;
	reg [31:0] r_927_0;
	reg [31:0] r_928_0;
	reg [31:0] r_929_0;
	reg [31:0] r_930_0;
	reg [31:0] r_931_0;
	reg [31:0] r_932_0;
	reg [31:0] r_933_0;
	reg [31:0] r_934_0;
	reg [31:0] r_935_0;
	reg [31:0] r_936_0;
	reg [31:0] r_937_0;
	reg [31:0] r_938_0;
	reg [31:0] r_939_0;
	reg [31:0] r_940_0;
	reg [31:0] r_941_0;
	reg [31:0] r_942_0;
	reg [31:0] r_943_0;
	reg [31:0] r_944_0;
	reg [31:0] r_945_0;
	reg [31:0] r_946_0;
	reg [31:0] r_947_0;
	reg [31:0] r_948_0;
	reg [31:0] r_949_0;
	reg [31:0] r_950_0;
	reg [31:0] r_951_0;
	reg [31:0] r_952_0;
	reg [31:0] r_953_0;
	reg [31:0] r_954_0;
	reg [31:0] r_955_0;
	reg [31:0] r_956_0;
	reg [31:0] r_957_0;
	reg [31:0] r_958_0;
	reg [31:0] r_959_0;
	reg [31:0] r_960_0;
	reg [31:0] r_961_0;
	reg [31:0] r_962_0;
	reg [31:0] r_963_0;
	reg [31:0] r_964_0;
	reg [31:0] r_965_0;
	reg [31:0] r_966_0;
	reg [31:0] r_967_0;
	reg [31:0] r_968_0;
	reg [31:0] r_969_0;
	reg [31:0] r_970_0;
	reg [31:0] r_971_0;
	reg [31:0] r_972_0;
	reg [31:0] r_973_0;
	reg [31:0] r_974_0;
	reg [31:0] r_975_0;
	reg [31:0] r_976_0;
	reg [31:0] r_977_0;
	reg [31:0] r_978_0;
	reg [31:0] r_979_0;
	reg [31:0] r_980_0;
	reg [31:0] r_981_0;
	reg [31:0] r_982_0;
	reg [31:0] r_983_0;
	reg [31:0] r_984_0;
	reg [31:0] r_985_0;
	reg [31:0] r_986_0;
	reg [31:0] r_987_0;
	reg [31:0] r_988_0;
	reg [31:0] r_989_0;
	reg [31:0] r_990_0;
	reg [31:0] r_991_0;
	reg [31:0] r_992_0;
	reg [31:0] r_993_0;
	reg [31:0] r_994_0;
	reg [31:0] r_995_0;
	reg [31:0] r_996_0;
	reg [31:0] r_997_0;
	reg [31:0] r_998_0;
	reg [31:0] r_999_0;
	reg [31:0] r_1000_0;
	reg [31:0] r_1001_0;
	reg [31:0] r_1002_0;
	reg [31:0] r_1003_0;
	reg [31:0] r_1004_0;
	reg [31:0] r_1005_0;
	reg [31:0] r_1006_0;
	reg [31:0] r_1007_0;
	reg [31:0] r_1008_0;
	reg [31:0] r_1009_0;
	reg [31:0] r_1010_0;
	reg [31:0] r_1011_0;
	reg [31:0] r_1012_0;
	reg [31:0] r_1013_0;
	reg [31:0] r_1014_0;
	reg [31:0] r_1015_0;
	reg [31:0] r_1016_0;
	reg [31:0] r_1017_0;
	reg [31:0] r_1018_0;
	reg [31:0] r_1019_0;
	reg [31:0] r_1020_0;
	reg [31:0] r_1021_0;
	reg [31:0] r_1022_0;
	reg [31:0] r_1023_0;
	reg [31:0] b_0;
	reg [31:0] b_1_0;
	reg [31:0] b_2_0;
	reg [31:0] b_3_0;
	reg [31:0] b_4_0;
	reg [31:0] b_5_0;
	reg [31:0] b_6_0;
	reg [31:0] b_7_0;
	reg [31:0] b_8_0;
	reg [31:0] b_9_0;
	reg [31:0] b_10_0;
	reg [31:0] b_11_0;
	reg [31:0] b_12_0;
	reg [31:0] b_13_0;
	reg [31:0] b_14_0;
	reg [31:0] b_15_0;
	reg [31:0] b_16_0;
	reg [31:0] b_17_0;
	reg [31:0] b_18_0;
	reg [31:0] b_19_0;
	reg [31:0] b_20_0;
	reg [31:0] b_21_0;
	reg [31:0] b_22_0;
	reg [31:0] b_23_0;
	reg [31:0] b_24_0;
	reg [31:0] b_25_0;
	reg [31:0] b_26_0;
	reg [31:0] b_27_0;
	reg [31:0] b_28_0;
	reg [31:0] b_29_0;
	reg [31:0] b_30_0;
	reg [31:0] b_31_0;
	reg [31:0] b_32_0;
	reg [31:0] b_33_0;
	reg [31:0] b_34_0;
	reg [31:0] b_35_0;
	reg [31:0] b_36_0;
	reg [31:0] b_37_0;
	reg [31:0] b_38_0;
	reg [31:0] b_39_0;
	reg [31:0] b_40_0;
	reg [31:0] b_41_0;
	reg [31:0] b_42_0;
	reg [31:0] b_43_0;
	reg [31:0] b_44_0;
	reg [31:0] b_45_0;
	reg [31:0] b_46_0;
	reg [31:0] b_47_0;
	reg [31:0] b_48_0;
	reg [31:0] b_49_0;
	reg [31:0] b_50_0;
	reg [31:0] b_51_0;
	reg [31:0] b_52_0;
	reg [31:0] b_53_0;
	reg [31:0] b_54_0;
	reg [31:0] b_55_0;
	reg [31:0] b_56_0;
	reg [31:0] b_57_0;
	reg [31:0] b_58_0;
	reg [31:0] b_59_0;
	reg [31:0] b_60_0;
	reg [31:0] b_61_0;
	reg [31:0] b_62_0;
	reg [31:0] b_63_0;
	reg [31:0] b_64_0;
	reg [31:0] b_65_0;
	reg [31:0] b_66_0;
	reg [31:0] b_67_0;
	reg [31:0] b_68_0;
	reg [31:0] b_69_0;
	reg [31:0] b_70_0;
	reg [31:0] b_71_0;
	reg [31:0] b_72_0;
	reg [31:0] b_73_0;
	reg [31:0] b_74_0;
	reg [31:0] b_75_0;
	reg [31:0] b_76_0;
	reg [31:0] b_77_0;
	reg [31:0] b_78_0;
	reg [31:0] b_79_0;
	reg [31:0] b_80_0;
	reg [31:0] b_81_0;
	reg [31:0] b_82_0;
	reg [31:0] b_83_0;
	reg [31:0] b_84_0;
	reg [31:0] b_85_0;
	reg [31:0] b_86_0;
	reg [31:0] b_87_0;
	reg [31:0] b_88_0;
	reg [31:0] b_89_0;
	reg [31:0] b_90_0;
	reg [31:0] b_91_0;
	reg [31:0] b_92_0;
	reg [31:0] b_93_0;
	reg [31:0] b_94_0;
	reg [31:0] b_95_0;
	reg [31:0] b_96_0;
	reg [31:0] b_97_0;
	reg [31:0] b_98_0;
	reg [31:0] b_99_0;
	reg [31:0] b_100_0;
	reg [31:0] b_101_0;
	reg [31:0] b_102_0;
	reg [31:0] b_103_0;
	reg [31:0] b_104_0;
	reg [31:0] b_105_0;
	reg [31:0] b_106_0;
	reg [31:0] b_107_0;
	reg [31:0] b_108_0;
	reg [31:0] b_109_0;
	reg [31:0] b_110_0;
	reg [31:0] b_111_0;
	reg [31:0] b_112_0;
	reg [31:0] b_113_0;
	reg [31:0] b_114_0;
	reg [31:0] b_115_0;
	reg [31:0] b_116_0;
	reg [31:0] b_117_0;
	reg [31:0] b_118_0;
	reg [31:0] b_119_0;
	reg [31:0] b_120_0;
	reg [31:0] b_121_0;
	reg [31:0] b_122_0;
	reg [31:0] b_123_0;
	reg [31:0] b_124_0;
	reg [31:0] b_125_0;
	reg [31:0] b_126_0;
	reg [31:0] b_127_0;
	reg [31:0] b_128_0;
	reg [31:0] b_129_0;
	reg [31:0] b_130_0;
	reg [31:0] b_131_0;
	reg [31:0] b_132_0;
	reg [31:0] b_133_0;
	reg [31:0] b_134_0;
	reg [31:0] b_135_0;
	reg [31:0] b_136_0;
	reg [31:0] b_137_0;
	reg [31:0] b_138_0;
	reg [31:0] b_139_0;
	reg [31:0] b_140_0;
	reg [31:0] b_141_0;
	reg [31:0] b_142_0;
	reg [31:0] b_143_0;
	reg [31:0] b_144_0;
	reg [31:0] b_145_0;
	reg [31:0] b_146_0;
	reg [31:0] b_147_0;
	reg [31:0] b_148_0;
	reg [31:0] b_149_0;
	reg [31:0] b_150_0;
	reg [31:0] b_151_0;
	reg [31:0] b_152_0;
	reg [31:0] b_153_0;
	reg [31:0] b_154_0;
	reg [31:0] b_155_0;
	reg [31:0] b_156_0;
	reg [31:0] b_157_0;
	reg [31:0] b_158_0;
	reg [31:0] b_159_0;
	reg [31:0] b_160_0;
	reg [31:0] b_161_0;
	reg [31:0] b_162_0;
	reg [31:0] b_163_0;
	reg [31:0] b_164_0;
	reg [31:0] b_165_0;
	reg [31:0] b_166_0;
	reg [31:0] b_167_0;
	reg [31:0] b_168_0;
	reg [31:0] b_169_0;
	reg [31:0] b_170_0;
	reg [31:0] b_171_0;
	reg [31:0] b_172_0;
	reg [31:0] b_173_0;
	reg [31:0] b_174_0;
	reg [31:0] b_175_0;
	reg [31:0] b_176_0;
	reg [31:0] b_177_0;
	reg [31:0] b_178_0;
	reg [31:0] b_179_0;
	reg [31:0] b_180_0;
	reg [31:0] b_181_0;
	reg [31:0] b_182_0;
	reg [31:0] b_183_0;
	reg [31:0] b_184_0;
	reg [31:0] b_185_0;
	reg [31:0] b_186_0;
	reg [31:0] b_187_0;
	reg [31:0] b_188_0;
	reg [31:0] b_189_0;
	reg [31:0] b_190_0;
	reg [31:0] b_191_0;
	reg [31:0] b_192_0;
	reg [31:0] b_193_0;
	reg [31:0] b_194_0;
	reg [31:0] b_195_0;
	reg [31:0] b_196_0;
	reg [31:0] b_197_0;
	reg [31:0] b_198_0;
	reg [31:0] b_199_0;
	reg [31:0] b_200_0;
	reg [31:0] b_201_0;
	reg [31:0] b_202_0;
	reg [31:0] b_203_0;
	reg [31:0] b_204_0;
	reg [31:0] b_205_0;
	reg [31:0] b_206_0;
	reg [31:0] b_207_0;
	reg [31:0] b_208_0;
	reg [31:0] b_209_0;
	reg [31:0] b_210_0;
	reg [31:0] b_211_0;
	reg [31:0] b_212_0;
	reg [31:0] b_213_0;
	reg [31:0] b_214_0;
	reg [31:0] b_215_0;
	reg [31:0] b_216_0;
	reg [31:0] b_217_0;
	reg [31:0] b_218_0;
	reg [31:0] b_219_0;
	reg [31:0] b_220_0;
	reg [31:0] b_221_0;
	reg [31:0] b_222_0;
	reg [31:0] b_223_0;
	reg [31:0] b_224_0;
	reg [31:0] b_225_0;
	reg [31:0] b_226_0;
	reg [31:0] b_227_0;
	reg [31:0] b_228_0;
	reg [31:0] b_229_0;
	reg [31:0] b_230_0;
	reg [31:0] b_231_0;
	reg [31:0] b_232_0;
	reg [31:0] b_233_0;
	reg [31:0] b_234_0;
	reg [31:0] b_235_0;
	reg [31:0] b_236_0;
	reg [31:0] b_237_0;
	reg [31:0] b_238_0;
	reg [31:0] b_239_0;
	reg [31:0] b_240_0;
	reg [31:0] b_241_0;
	reg [31:0] b_242_0;
	reg [31:0] b_243_0;
	reg [31:0] b_244_0;
	reg [31:0] b_245_0;
	reg [31:0] b_246_0;
	reg [31:0] b_247_0;
	reg [31:0] b_248_0;
	reg [31:0] b_249_0;
	reg [31:0] b_250_0;
	reg [31:0] b_251_0;
	reg [31:0] b_252_0;
	reg [31:0] b_253_0;
	reg [31:0] b_254_0;
	reg [31:0] b_255_0;
	reg [31:0] b_256_0;
	reg [31:0] b_257_0;
	reg [31:0] b_258_0;
	reg [31:0] b_259_0;
	reg [31:0] b_260_0;
	reg [31:0] b_261_0;
	reg [31:0] b_262_0;
	reg [31:0] b_263_0;
	reg [31:0] b_264_0;
	reg [31:0] b_265_0;
	reg [31:0] b_266_0;
	reg [31:0] b_267_0;
	reg [31:0] b_268_0;
	reg [31:0] b_269_0;
	reg [31:0] b_270_0;
	reg [31:0] b_271_0;
	reg [31:0] b_272_0;
	reg [31:0] b_273_0;
	reg [31:0] b_274_0;
	reg [31:0] b_275_0;
	reg [31:0] b_276_0;
	reg [31:0] b_277_0;
	reg [31:0] b_278_0;
	reg [31:0] b_279_0;
	reg [31:0] b_280_0;
	reg [31:0] b_281_0;
	reg [31:0] b_282_0;
	reg [31:0] b_283_0;
	reg [31:0] b_284_0;
	reg [31:0] b_285_0;
	reg [31:0] b_286_0;
	reg [31:0] b_287_0;
	reg [31:0] b_288_0;
	reg [31:0] b_289_0;
	reg [31:0] b_290_0;
	reg [31:0] b_291_0;
	reg [31:0] b_292_0;
	reg [31:0] b_293_0;
	reg [31:0] b_294_0;
	reg [31:0] b_295_0;
	reg [31:0] b_296_0;
	reg [31:0] b_297_0;
	reg [31:0] b_298_0;
	reg [31:0] b_299_0;
	reg [31:0] b_300_0;
	reg [31:0] b_301_0;
	reg [31:0] b_302_0;
	reg [31:0] b_303_0;
	reg [31:0] b_304_0;
	reg [31:0] b_305_0;
	reg [31:0] b_306_0;
	reg [31:0] b_307_0;
	reg [31:0] b_308_0;
	reg [31:0] b_309_0;
	reg [31:0] b_310_0;
	reg [31:0] b_311_0;
	reg [31:0] b_312_0;
	reg [31:0] b_313_0;
	reg [31:0] b_314_0;
	reg [31:0] b_315_0;
	reg [31:0] b_316_0;
	reg [31:0] b_317_0;
	reg [31:0] b_318_0;
	reg [31:0] b_319_0;
	reg [31:0] b_320_0;
	reg [31:0] b_321_0;
	reg [31:0] b_322_0;
	reg [31:0] b_323_0;
	reg [31:0] b_324_0;
	reg [31:0] b_325_0;
	reg [31:0] b_326_0;
	reg [31:0] b_327_0;
	reg [31:0] b_328_0;
	reg [31:0] b_329_0;
	reg [31:0] b_330_0;
	reg [31:0] b_331_0;
	reg [31:0] b_332_0;
	reg [31:0] b_333_0;
	reg [31:0] b_334_0;
	reg [31:0] b_335_0;
	reg [31:0] b_336_0;
	reg [31:0] b_337_0;
	reg [31:0] b_338_0;
	reg [31:0] b_339_0;
	reg [31:0] b_340_0;
	reg [31:0] b_341_0;
	reg [31:0] b_342_0;
	reg [31:0] b_343_0;
	reg [31:0] b_344_0;
	reg [31:0] b_345_0;
	reg [31:0] b_346_0;
	reg [31:0] b_347_0;
	reg [31:0] b_348_0;
	reg [31:0] b_349_0;
	reg [31:0] b_350_0;
	reg [31:0] b_351_0;
	reg [31:0] b_352_0;
	reg [31:0] b_353_0;
	reg [31:0] b_354_0;
	reg [31:0] b_355_0;
	reg [31:0] b_356_0;
	reg [31:0] b_357_0;
	reg [31:0] b_358_0;
	reg [31:0] b_359_0;
	reg [31:0] b_360_0;
	reg [31:0] b_361_0;
	reg [31:0] b_362_0;
	reg [31:0] b_363_0;
	reg [31:0] b_364_0;
	reg [31:0] b_365_0;
	reg [31:0] b_366_0;
	reg [31:0] b_367_0;
	reg [31:0] b_368_0;
	reg [31:0] b_369_0;
	reg [31:0] b_370_0;
	reg [31:0] b_371_0;
	reg [31:0] b_372_0;
	reg [31:0] b_373_0;
	reg [31:0] b_374_0;
	reg [31:0] b_375_0;
	reg [31:0] b_376_0;
	reg [31:0] b_377_0;
	reg [31:0] b_378_0;
	reg [31:0] b_379_0;
	reg [31:0] b_380_0;
	reg [31:0] b_381_0;
	reg [31:0] b_382_0;
	reg [31:0] b_383_0;
	reg [31:0] b_384_0;
	reg [31:0] b_385_0;
	reg [31:0] b_386_0;
	reg [31:0] b_387_0;
	reg [31:0] b_388_0;
	reg [31:0] b_389_0;
	reg [31:0] b_390_0;
	reg [31:0] b_391_0;
	reg [31:0] b_392_0;
	reg [31:0] b_393_0;
	reg [31:0] b_394_0;
	reg [31:0] b_395_0;
	reg [31:0] b_396_0;
	reg [31:0] b_397_0;
	reg [31:0] b_398_0;
	reg [31:0] b_399_0;
	reg [31:0] b_400_0;
	reg [31:0] b_401_0;
	reg [31:0] b_402_0;
	reg [31:0] b_403_0;
	reg [31:0] b_404_0;
	reg [31:0] b_405_0;
	reg [31:0] b_406_0;
	reg [31:0] b_407_0;
	reg [31:0] b_408_0;
	reg [31:0] b_409_0;
	reg [31:0] b_410_0;
	reg [31:0] b_411_0;
	reg [31:0] b_412_0;
	reg [31:0] b_413_0;
	reg [31:0] b_414_0;
	reg [31:0] b_415_0;
	reg [31:0] b_416_0;
	reg [31:0] b_417_0;
	reg [31:0] b_418_0;
	reg [31:0] b_419_0;
	reg [31:0] b_420_0;
	reg [31:0] b_421_0;
	reg [31:0] b_422_0;
	reg [31:0] b_423_0;
	reg [31:0] b_424_0;
	reg [31:0] b_425_0;
	reg [31:0] b_426_0;
	reg [31:0] b_427_0;
	reg [31:0] b_428_0;
	reg [31:0] b_429_0;
	reg [31:0] b_430_0;
	reg [31:0] b_431_0;
	reg [31:0] b_432_0;
	reg [31:0] b_433_0;
	reg [31:0] b_434_0;
	reg [31:0] b_435_0;
	reg [31:0] b_436_0;
	reg [31:0] b_437_0;
	reg [31:0] b_438_0;
	reg [31:0] b_439_0;
	reg [31:0] b_440_0;
	reg [31:0] b_441_0;
	reg [31:0] b_442_0;
	reg [31:0] b_443_0;
	reg [31:0] b_444_0;
	reg [31:0] b_445_0;
	reg [31:0] b_446_0;
	reg [31:0] b_447_0;
	reg [31:0] b_448_0;
	reg [31:0] b_449_0;
	reg [31:0] b_450_0;
	reg [31:0] b_451_0;
	reg [31:0] b_452_0;
	reg [31:0] b_453_0;
	reg [31:0] b_454_0;
	reg [31:0] b_455_0;
	reg [31:0] b_456_0;
	reg [31:0] b_457_0;
	reg [31:0] b_458_0;
	reg [31:0] b_459_0;
	reg [31:0] b_460_0;
	reg [31:0] b_461_0;
	reg [31:0] b_462_0;
	reg [31:0] b_463_0;
	reg [31:0] b_464_0;
	reg [31:0] b_465_0;
	reg [31:0] b_466_0;
	reg [31:0] b_467_0;
	reg [31:0] b_468_0;
	reg [31:0] b_469_0;
	reg [31:0] b_470_0;
	reg [31:0] b_471_0;
	reg [31:0] b_472_0;
	reg [31:0] b_473_0;
	reg [31:0] b_474_0;
	reg [31:0] b_475_0;
	reg [31:0] b_476_0;
	reg [31:0] b_477_0;
	reg [31:0] b_478_0;
	reg [31:0] b_479_0;
	reg [31:0] b_480_0;
	reg [31:0] b_481_0;
	reg [31:0] b_482_0;
	reg [31:0] b_483_0;
	reg [31:0] b_484_0;
	reg [31:0] b_485_0;
	reg [31:0] b_486_0;
	reg [31:0] b_487_0;
	reg [31:0] b_488_0;
	reg [31:0] b_489_0;
	reg [31:0] b_490_0;
	reg [31:0] b_491_0;
	reg [31:0] b_492_0;
	reg [31:0] b_493_0;
	reg [31:0] b_494_0;
	reg [31:0] b_495_0;
	reg [31:0] b_496_0;
	reg [31:0] b_497_0;
	reg [31:0] b_498_0;
	reg [31:0] b_499_0;
	reg [31:0] b_500_0;
	reg [31:0] b_501_0;
	reg [31:0] b_502_0;
	reg [31:0] b_503_0;
	reg [31:0] b_504_0;
	reg [31:0] b_505_0;
	reg [31:0] b_506_0;
	reg [31:0] b_507_0;
	reg [31:0] b_508_0;
	reg [31:0] b_509_0;
	reg [31:0] b_510_0;
	reg [31:0] b_511_0;
	reg [31:0] b_512_0;
	reg [31:0] b_513_0;
	reg [31:0] b_514_0;
	reg [31:0] b_515_0;
	reg [31:0] b_516_0;
	reg [31:0] b_517_0;
	reg [31:0] b_518_0;
	reg [31:0] b_519_0;
	reg [31:0] b_520_0;
	reg [31:0] b_521_0;
	reg [31:0] b_522_0;
	reg [31:0] b_523_0;
	reg [31:0] b_524_0;
	reg [31:0] b_525_0;
	reg [31:0] b_526_0;
	reg [31:0] b_527_0;
	reg [31:0] b_528_0;
	reg [31:0] b_529_0;
	reg [31:0] b_530_0;
	reg [31:0] b_531_0;
	reg [31:0] b_532_0;
	reg [31:0] b_533_0;
	reg [31:0] b_534_0;
	reg [31:0] b_535_0;
	reg [31:0] b_536_0;
	reg [31:0] b_537_0;
	reg [31:0] b_538_0;
	reg [31:0] b_539_0;
	reg [31:0] b_540_0;
	reg [31:0] b_541_0;
	reg [31:0] b_542_0;
	reg [31:0] b_543_0;
	reg [31:0] b_544_0;
	reg [31:0] b_545_0;
	reg [31:0] b_546_0;
	reg [31:0] b_547_0;
	reg [31:0] b_548_0;
	reg [31:0] b_549_0;
	reg [31:0] b_550_0;
	reg [31:0] b_551_0;
	reg [31:0] b_552_0;
	reg [31:0] b_553_0;
	reg [31:0] b_554_0;
	reg [31:0] b_555_0;
	reg [31:0] b_556_0;
	reg [31:0] b_557_0;
	reg [31:0] b_558_0;
	reg [31:0] b_559_0;
	reg [31:0] b_560_0;
	reg [31:0] b_561_0;
	reg [31:0] b_562_0;
	reg [31:0] b_563_0;
	reg [31:0] b_564_0;
	reg [31:0] b_565_0;
	reg [31:0] b_566_0;
	reg [31:0] b_567_0;
	reg [31:0] b_568_0;
	reg [31:0] b_569_0;
	reg [31:0] b_570_0;
	reg [31:0] b_571_0;
	reg [31:0] b_572_0;
	reg [31:0] b_573_0;
	reg [31:0] b_574_0;
	reg [31:0] b_575_0;
	reg [31:0] b_576_0;
	reg [31:0] b_577_0;
	reg [31:0] b_578_0;
	reg [31:0] b_579_0;
	reg [31:0] b_580_0;
	reg [31:0] b_581_0;
	reg [31:0] b_582_0;
	reg [31:0] b_583_0;
	reg [31:0] b_584_0;
	reg [31:0] b_585_0;
	reg [31:0] b_586_0;
	reg [31:0] b_587_0;
	reg [31:0] b_588_0;
	reg [31:0] b_589_0;
	reg [31:0] b_590_0;
	reg [31:0] b_591_0;
	reg [31:0] b_592_0;
	reg [31:0] b_593_0;
	reg [31:0] b_594_0;
	reg [31:0] b_595_0;
	reg [31:0] b_596_0;
	reg [31:0] b_597_0;
	reg [31:0] b_598_0;
	reg [31:0] b_599_0;
	reg [31:0] b_600_0;
	reg [31:0] b_601_0;
	reg [31:0] b_602_0;
	reg [31:0] b_603_0;
	reg [31:0] b_604_0;
	reg [31:0] b_605_0;
	reg [31:0] b_606_0;
	reg [31:0] b_607_0;
	reg [31:0] b_608_0;
	reg [31:0] b_609_0;
	reg [31:0] b_610_0;
	reg [31:0] b_611_0;
	reg [31:0] b_612_0;
	reg [31:0] b_613_0;
	reg [31:0] b_614_0;
	reg [31:0] b_615_0;
	reg [31:0] b_616_0;
	reg [31:0] b_617_0;
	reg [31:0] b_618_0;
	reg [31:0] b_619_0;
	reg [31:0] b_620_0;
	reg [31:0] b_621_0;
	reg [31:0] b_622_0;
	reg [31:0] b_623_0;
	reg [31:0] b_624_0;
	reg [31:0] b_625_0;
	reg [31:0] b_626_0;
	reg [31:0] b_627_0;
	reg [31:0] b_628_0;
	reg [31:0] b_629_0;
	reg [31:0] b_630_0;
	reg [31:0] b_631_0;
	reg [31:0] b_632_0;
	reg [31:0] b_633_0;
	reg [31:0] b_634_0;
	reg [31:0] b_635_0;
	reg [31:0] b_636_0;
	reg [31:0] b_637_0;
	reg [31:0] b_638_0;
	reg [31:0] b_639_0;
	reg [31:0] b_640_0;
	reg [31:0] b_641_0;
	reg [31:0] b_642_0;
	reg [31:0] b_643_0;
	reg [31:0] b_644_0;
	reg [31:0] b_645_0;
	reg [31:0] b_646_0;
	reg [31:0] b_647_0;
	reg [31:0] b_648_0;
	reg [31:0] b_649_0;
	reg [31:0] b_650_0;
	reg [31:0] b_651_0;
	reg [31:0] b_652_0;
	reg [31:0] b_653_0;
	reg [31:0] b_654_0;
	reg [31:0] b_655_0;
	reg [31:0] b_656_0;
	reg [31:0] b_657_0;
	reg [31:0] b_658_0;
	reg [31:0] b_659_0;
	reg [31:0] b_660_0;
	reg [31:0] b_661_0;
	reg [31:0] b_662_0;
	reg [31:0] b_663_0;
	reg [31:0] b_664_0;
	reg [31:0] b_665_0;
	reg [31:0] b_666_0;
	reg [31:0] b_667_0;
	reg [31:0] b_668_0;
	reg [31:0] b_669_0;
	reg [31:0] b_670_0;
	reg [31:0] b_671_0;
	reg [31:0] b_672_0;
	reg [31:0] b_673_0;
	reg [31:0] b_674_0;
	reg [31:0] b_675_0;
	reg [31:0] b_676_0;
	reg [31:0] b_677_0;
	reg [31:0] b_678_0;
	reg [31:0] b_679_0;
	reg [31:0] b_680_0;
	reg [31:0] b_681_0;
	reg [31:0] b_682_0;
	reg [31:0] b_683_0;
	reg [31:0] b_684_0;
	reg [31:0] b_685_0;
	reg [31:0] b_686_0;
	reg [31:0] b_687_0;
	reg [31:0] b_688_0;
	reg [31:0] b_689_0;
	reg [31:0] b_690_0;
	reg [31:0] b_691_0;
	reg [31:0] b_692_0;
	reg [31:0] b_693_0;
	reg [31:0] b_694_0;
	reg [31:0] b_695_0;
	reg [31:0] b_696_0;
	reg [31:0] b_697_0;
	reg [31:0] b_698_0;
	reg [31:0] b_699_0;
	reg [31:0] b_700_0;
	reg [31:0] b_701_0;
	reg [31:0] b_702_0;
	reg [31:0] b_703_0;
	reg [31:0] b_704_0;
	reg [31:0] b_705_0;
	reg [31:0] b_706_0;
	reg [31:0] b_707_0;
	reg [31:0] b_708_0;
	reg [31:0] b_709_0;
	reg [31:0] b_710_0;
	reg [31:0] b_711_0;
	reg [31:0] b_712_0;
	reg [31:0] b_713_0;
	reg [31:0] b_714_0;
	reg [31:0] b_715_0;
	reg [31:0] b_716_0;
	reg [31:0] b_717_0;
	reg [31:0] b_718_0;
	reg [31:0] b_719_0;
	reg [31:0] b_720_0;
	reg [31:0] b_721_0;
	reg [31:0] b_722_0;
	reg [31:0] b_723_0;
	reg [31:0] b_724_0;
	reg [31:0] b_725_0;
	reg [31:0] b_726_0;
	reg [31:0] b_727_0;
	reg [31:0] b_728_0;
	reg [31:0] b_729_0;
	reg [31:0] b_730_0;
	reg [31:0] b_731_0;
	reg [31:0] b_732_0;
	reg [31:0] b_733_0;
	reg [31:0] b_734_0;
	reg [31:0] b_735_0;
	reg [31:0] b_736_0;
	reg [31:0] b_737_0;
	reg [31:0] b_738_0;
	reg [31:0] b_739_0;
	reg [31:0] b_740_0;
	reg [31:0] b_741_0;
	reg [31:0] b_742_0;
	reg [31:0] b_743_0;
	reg [31:0] b_744_0;
	reg [31:0] b_745_0;
	reg [31:0] b_746_0;
	reg [31:0] b_747_0;
	reg [31:0] b_748_0;
	reg [31:0] b_749_0;
	reg [31:0] b_750_0;
	reg [31:0] b_751_0;
	reg [31:0] b_752_0;
	reg [31:0] b_753_0;
	reg [31:0] b_754_0;
	reg [31:0] b_755_0;
	reg [31:0] b_756_0;
	reg [31:0] b_757_0;
	reg [31:0] b_758_0;
	reg [31:0] b_759_0;
	reg [31:0] b_760_0;
	reg [31:0] b_761_0;
	reg [31:0] b_762_0;
	reg [31:0] b_763_0;
	reg [31:0] b_764_0;
	reg [31:0] b_765_0;
	reg [31:0] b_766_0;
	reg [31:0] b_767_0;
	reg [31:0] b_768_0;
	reg [31:0] b_769_0;
	reg [31:0] b_770_0;
	reg [31:0] b_771_0;
	reg [31:0] b_772_0;
	reg [31:0] b_773_0;
	reg [31:0] b_774_0;
	reg [31:0] b_775_0;
	reg [31:0] b_776_0;
	reg [31:0] b_777_0;
	reg [31:0] b_778_0;
	reg [31:0] b_779_0;
	reg [31:0] b_780_0;
	reg [31:0] b_781_0;
	reg [31:0] b_782_0;
	reg [31:0] b_783_0;
	reg [31:0] b_784_0;
	reg [31:0] b_785_0;
	reg [31:0] b_786_0;
	reg [31:0] b_787_0;
	reg [31:0] b_788_0;
	reg [31:0] b_789_0;
	reg [31:0] b_790_0;
	reg [31:0] b_791_0;
	reg [31:0] b_792_0;
	reg [31:0] b_793_0;
	reg [31:0] b_794_0;
	reg [31:0] b_795_0;
	reg [31:0] b_796_0;
	reg [31:0] b_797_0;
	reg [31:0] b_798_0;
	reg [31:0] b_799_0;
	reg [31:0] b_800_0;
	reg [31:0] b_801_0;
	reg [31:0] b_802_0;
	reg [31:0] b_803_0;
	reg [31:0] b_804_0;
	reg [31:0] b_805_0;
	reg [31:0] b_806_0;
	reg [31:0] b_807_0;
	reg [31:0] b_808_0;
	reg [31:0] b_809_0;
	reg [31:0] b_810_0;
	reg [31:0] b_811_0;
	reg [31:0] b_812_0;
	reg [31:0] b_813_0;
	reg [31:0] b_814_0;
	reg [31:0] b_815_0;
	reg [31:0] b_816_0;
	reg [31:0] b_817_0;
	reg [31:0] b_818_0;
	reg [31:0] b_819_0;
	reg [31:0] b_820_0;
	reg [31:0] b_821_0;
	reg [31:0] b_822_0;
	reg [31:0] b_823_0;
	reg [31:0] b_824_0;
	reg [31:0] b_825_0;
	reg [31:0] b_826_0;
	reg [31:0] b_827_0;
	reg [31:0] b_828_0;
	reg [31:0] b_829_0;
	reg [31:0] b_830_0;
	reg [31:0] b_831_0;
	reg [31:0] b_832_0;
	reg [31:0] b_833_0;
	reg [31:0] b_834_0;
	reg [31:0] b_835_0;
	reg [31:0] b_836_0;
	reg [31:0] b_837_0;
	reg [31:0] b_838_0;
	reg [31:0] b_839_0;
	reg [31:0] b_840_0;
	reg [31:0] b_841_0;
	reg [31:0] b_842_0;
	reg [31:0] b_843_0;
	reg [31:0] b_844_0;
	reg [31:0] b_845_0;
	reg [31:0] b_846_0;
	reg [31:0] b_847_0;
	reg [31:0] b_848_0;
	reg [31:0] b_849_0;
	reg [31:0] b_850_0;
	reg [31:0] b_851_0;
	reg [31:0] b_852_0;
	reg [31:0] b_853_0;
	reg [31:0] b_854_0;
	reg [31:0] b_855_0;
	reg [31:0] b_856_0;
	reg [31:0] b_857_0;
	reg [31:0] b_858_0;
	reg [31:0] b_859_0;
	reg [31:0] b_860_0;
	reg [31:0] b_861_0;
	reg [31:0] b_862_0;
	reg [31:0] b_863_0;
	reg [31:0] b_864_0;
	reg [31:0] b_865_0;
	reg [31:0] b_866_0;
	reg [31:0] b_867_0;
	reg [31:0] b_868_0;
	reg [31:0] b_869_0;
	reg [31:0] b_870_0;
	reg [31:0] b_871_0;
	reg [31:0] b_872_0;
	reg [31:0] b_873_0;
	reg [31:0] b_874_0;
	reg [31:0] b_875_0;
	reg [31:0] b_876_0;
	reg [31:0] b_877_0;
	reg [31:0] b_878_0;
	reg [31:0] b_879_0;
	reg [31:0] b_880_0;
	reg [31:0] b_881_0;
	reg [31:0] b_882_0;
	reg [31:0] b_883_0;
	reg [31:0] b_884_0;
	reg [31:0] b_885_0;
	reg [31:0] b_886_0;
	reg [31:0] b_887_0;
	reg [31:0] b_888_0;
	reg [31:0] b_889_0;
	reg [31:0] b_890_0;
	reg [31:0] b_891_0;
	reg [31:0] b_892_0;
	reg [31:0] b_893_0;
	reg [31:0] b_894_0;
	reg [31:0] b_895_0;
	reg [31:0] b_896_0;
	reg [31:0] b_897_0;
	reg [31:0] b_898_0;
	reg [31:0] b_899_0;
	reg [31:0] b_900_0;
	reg [31:0] b_901_0;
	reg [31:0] b_902_0;
	reg [31:0] b_903_0;
	reg [31:0] b_904_0;
	reg [31:0] b_905_0;
	reg [31:0] b_906_0;
	reg [31:0] b_907_0;
	reg [31:0] b_908_0;
	reg [31:0] b_909_0;
	reg [31:0] b_910_0;
	reg [31:0] b_911_0;
	reg [31:0] b_912_0;
	reg [31:0] b_913_0;
	reg [31:0] b_914_0;
	reg [31:0] b_915_0;
	reg [31:0] b_916_0;
	reg [31:0] b_917_0;
	reg [31:0] b_918_0;
	reg [31:0] b_919_0;
	reg [31:0] b_920_0;
	reg [31:0] b_921_0;
	reg [31:0] b_922_0;
	reg [31:0] b_923_0;
	reg [31:0] b_924_0;
	reg [31:0] b_925_0;
	reg [31:0] b_926_0;
	reg [31:0] b_927_0;
	reg [31:0] b_928_0;
	reg [31:0] b_929_0;
	reg [31:0] b_930_0;
	reg [31:0] b_931_0;
	reg [31:0] b_932_0;
	reg [31:0] b_933_0;
	reg [31:0] b_934_0;
	reg [31:0] b_935_0;
	reg [31:0] b_936_0;
	reg [31:0] b_937_0;
	reg [31:0] b_938_0;
	reg [31:0] b_939_0;
	reg [31:0] b_940_0;
	reg [31:0] b_941_0;
	reg [31:0] b_942_0;
	reg [31:0] b_943_0;
	reg [31:0] b_944_0;
	reg [31:0] b_945_0;
	reg [31:0] b_946_0;
	reg [31:0] b_947_0;
	reg [31:0] b_948_0;
	reg [31:0] b_949_0;
	reg [31:0] b_950_0;
	reg [31:0] b_951_0;
	reg [31:0] b_952_0;
	reg [31:0] b_953_0;
	reg [31:0] b_954_0;
	reg [31:0] b_955_0;
	reg [31:0] b_956_0;
	reg [31:0] b_957_0;
	reg [31:0] b_958_0;
	reg [31:0] b_959_0;
	reg [31:0] b_960_0;
	reg [31:0] b_961_0;
	reg [31:0] b_962_0;
	reg [31:0] b_963_0;
	reg [31:0] b_964_0;
	reg [31:0] b_965_0;
	reg [31:0] b_966_0;
	reg [31:0] b_967_0;
	reg [31:0] b_968_0;
	reg [31:0] b_969_0;
	reg [31:0] b_970_0;
	reg [31:0] b_971_0;
	reg [31:0] b_972_0;
	reg [31:0] b_973_0;
	reg [31:0] b_974_0;
	reg [31:0] b_975_0;
	reg [31:0] b_976_0;
	reg [31:0] b_977_0;
	reg [31:0] b_978_0;
	reg [31:0] b_979_0;
	reg [31:0] b_980_0;
	reg [31:0] b_981_0;
	reg [31:0] b_982_0;
	reg [31:0] b_983_0;
	reg [31:0] b_984_0;
	reg [31:0] b_985_0;
	reg [31:0] b_986_0;
	reg [31:0] b_987_0;
	reg [31:0] b_988_0;
	reg [31:0] b_989_0;
	reg [31:0] b_990_0;
	reg [31:0] b_991_0;
	reg [31:0] b_992_0;
	reg [31:0] b_993_0;
	reg [31:0] b_994_0;
	reg [31:0] b_995_0;
	reg [31:0] b_996_0;
	reg [31:0] b_997_0;
	reg [31:0] b_998_0;
	reg [31:0] b_999_0;
	reg [31:0] b_1000_0;
	reg [31:0] b_1001_0;
	reg [31:0] b_1002_0;
	reg [31:0] b_1003_0;
	reg [31:0] b_1004_0;
	reg [31:0] b_1005_0;
	reg [31:0] b_1006_0;
	reg [31:0] b_1007_0;
	reg [31:0] b_1008_0;
	reg [31:0] b_1009_0;
	reg [31:0] b_1010_0;
	reg [31:0] b_1011_0;
	reg [31:0] b_1012_0;
	reg [31:0] b_1013_0;
	reg [31:0] b_1014_0;
	reg [31:0] b_1015_0;
	reg [31:0] b_1016_0;
	reg [31:0] b_1017_0;
	reg [31:0] b_1018_0;
	reg [31:0] b_1019_0;
	reg [31:0] b_1020_0;
	reg [31:0] b_1021_0;
	reg [31:0] b_1022_0;
	reg [31:0] b_1023_0;
	reg [31:0] b_1024_0;
	reg [31:0] b_1025_0;
	reg [31:0] b_1026_0;
	reg [31:0] b_1027_0;
	reg [31:0] b_1028_0;
	reg [31:0] b_1029_0;
	reg [31:0] b_1030_0;
	reg [31:0] b_1031_0;
	reg [31:0] b_1032_0;
	reg [31:0] b_1033_0;
	reg [31:0] b_1034_0;
	reg [31:0] b_1035_0;
	reg [31:0] b_1036_0;
	reg [31:0] b_1037_0;
	reg [31:0] b_1038_0;
	reg [31:0] b_1039_0;
	reg [31:0] b_1040_0;
	reg [31:0] b_1041_0;
	reg [31:0] b_1042_0;
	reg [31:0] b_1043_0;
	reg [31:0] b_1044_0;
	reg [31:0] b_1045_0;
	reg [31:0] b_1046_0;
	reg [31:0] b_1047_0;
	reg [31:0] b_1048_0;
	reg [31:0] b_1049_0;
	reg [31:0] b_1050_0;
	reg [31:0] b_1051_0;
	reg [31:0] b_1052_0;
	reg [31:0] b_1053_0;
	reg [31:0] b_1054_0;
	reg [31:0] b_1055_0;
	reg [31:0] b_1056_0;
	reg [31:0] b_1057_0;
	reg [31:0] b_1058_0;
	reg [31:0] b_1059_0;
	reg [31:0] b_1060_0;
	reg [31:0] b_1061_0;
	reg [31:0] b_1062_0;
	reg [31:0] b_1063_0;
	reg [31:0] b_1064_0;
	reg [31:0] b_1065_0;
	reg [31:0] b_1066_0;
	reg [31:0] b_1067_0;
	reg [31:0] b_1068_0;
	reg [31:0] b_1069_0;
	reg [31:0] b_1070_0;
	reg [31:0] b_1071_0;
	reg [31:0] b_1072_0;
	reg [31:0] b_1073_0;
	reg [31:0] b_1074_0;
	reg [31:0] b_1075_0;
	reg [31:0] b_1076_0;
	reg [31:0] b_1077_0;
	reg [31:0] b_1078_0;
	reg [31:0] b_1079_0;
	reg [31:0] b_1080_0;
	reg [31:0] b_1081_0;
	reg [31:0] b_1082_0;
	reg [31:0] b_1083_0;
	reg [31:0] b_1084_0;
	reg [31:0] b_1085_0;
	reg [31:0] b_1086_0;
	reg [31:0] b_1087_0;
	reg [31:0] b_1088_0;
	reg [31:0] b_1089_0;
	reg [31:0] b_1090_0;
	reg [31:0] b_1091_0;
	reg [31:0] b_1092_0;
	reg [31:0] b_1093_0;
	reg [31:0] b_1094_0;
	reg [31:0] b_1095_0;
	reg [31:0] b_1096_0;
	reg [31:0] b_1097_0;
	reg [31:0] b_1098_0;
	reg [31:0] b_1099_0;
	reg [31:0] b_1100_0;
	reg [31:0] b_1101_0;
	reg [31:0] b_1102_0;
	reg [31:0] b_1103_0;
	reg [31:0] b_1104_0;
	reg [31:0] b_1105_0;
	reg [31:0] b_1106_0;
	reg [31:0] b_1107_0;
	reg [31:0] b_1108_0;
	reg [31:0] b_1109_0;
	reg [31:0] b_1110_0;
	reg [31:0] b_1111_0;
	reg [31:0] b_1112_0;
	reg [31:0] b_1113_0;
	reg [31:0] b_1114_0;
	reg [31:0] b_1115_0;
	reg [31:0] b_1116_0;
	reg [31:0] b_1117_0;
	reg [31:0] b_1118_0;
	reg [31:0] b_1119_0;
	reg [31:0] b_1120_0;
	reg [31:0] b_1121_0;
	reg [31:0] b_1122_0;
	reg [31:0] b_1123_0;
	reg [31:0] b_1124_0;
	reg [31:0] b_1125_0;
	reg [31:0] b_1126_0;
	reg [31:0] b_1127_0;
	reg [31:0] b_1128_0;
	reg [31:0] b_1129_0;
	reg [31:0] b_1130_0;
	reg [31:0] b_1131_0;
	reg [31:0] b_1132_0;
	reg [31:0] b_1133_0;
	reg [31:0] b_1134_0;
	reg [31:0] b_1135_0;
	reg [31:0] b_1136_0;
	reg [31:0] b_1137_0;
	reg [31:0] b_1138_0;
	reg [31:0] b_1139_0;
	reg [31:0] b_1140_0;
	reg [31:0] b_1141_0;
	reg [31:0] b_1142_0;
	reg [31:0] b_1143_0;
	reg [31:0] b_1144_0;
	reg [31:0] b_1145_0;
	reg [31:0] b_1146_0;
	reg [31:0] b_1147_0;
	reg [31:0] b_1148_0;
	reg [31:0] b_1149_0;
	reg [31:0] b_1150_0;
	reg [31:0] b_1151_0;
	reg [31:0] b_1152_0;
	reg [31:0] b_1153_0;
	reg [31:0] b_1154_0;
	reg [31:0] b_1155_0;
	reg [31:0] b_1156_0;
	reg [31:0] b_1157_0;
	reg [31:0] b_1158_0;
	reg [31:0] b_1159_0;
	reg [31:0] b_1160_0;
	reg [31:0] b_1161_0;
	reg [31:0] b_1162_0;
	reg [31:0] b_1163_0;
	reg [31:0] b_1164_0;
	reg [31:0] b_1165_0;
	reg [31:0] b_1166_0;
	reg [31:0] b_1167_0;
	reg [31:0] b_1168_0;
	reg [31:0] b_1169_0;
	reg [31:0] b_1170_0;
	reg [31:0] b_1171_0;
	reg [31:0] b_1172_0;
	reg [31:0] b_1173_0;
	reg [31:0] b_1174_0;
	reg [31:0] b_1175_0;
	reg [31:0] b_1176_0;
	reg [31:0] b_1177_0;
	reg [31:0] b_1178_0;
	reg [31:0] b_1179_0;
	reg [31:0] b_1180_0;
	reg [31:0] b_1181_0;
	reg [31:0] b_1182_0;
	reg [31:0] b_1183_0;
	reg [31:0] b_1184_0;
	reg [31:0] b_1185_0;
	reg [31:0] b_1186_0;
	reg [31:0] b_1187_0;
	reg [31:0] b_1188_0;
	reg [31:0] b_1189_0;
	reg [31:0] b_1190_0;
	reg [31:0] b_1191_0;
	reg [31:0] b_1192_0;
	reg [31:0] b_1193_0;
	reg [31:0] b_1194_0;
	reg [31:0] b_1195_0;
	reg [31:0] b_1196_0;
	reg [31:0] b_1197_0;
	reg [31:0] b_1198_0;
	reg [31:0] b_1199_0;
	reg [31:0] b_1200_0;
	reg [31:0] b_1201_0;
	reg [31:0] b_1202_0;
	reg [31:0] b_1203_0;
	reg [31:0] b_1204_0;
	reg [31:0] b_1205_0;
	reg [31:0] b_1206_0;
	reg [31:0] b_1207_0;
	reg [31:0] b_1208_0;
	reg [31:0] b_1209_0;
	reg [31:0] b_1210_0;
	reg [31:0] b_1211_0;
	reg [31:0] b_1212_0;
	reg [31:0] b_1213_0;
	reg [31:0] b_1214_0;
	reg [31:0] b_1215_0;
	reg [31:0] b_1216_0;
	reg [31:0] b_1217_0;
	reg [31:0] b_1218_0;
	reg [31:0] b_1219_0;
	reg [31:0] b_1220_0;
	reg [31:0] b_1221_0;
	reg [31:0] b_1222_0;
	reg [31:0] b_1223_0;
	reg [31:0] b_1224_0;
	reg [31:0] b_1225_0;
	reg [31:0] b_1226_0;
	reg [31:0] b_1227_0;
	reg [31:0] b_1228_0;
	reg [31:0] b_1229_0;
	reg [31:0] b_1230_0;
	reg [31:0] b_1231_0;
	reg [31:0] b_1232_0;
	reg [31:0] b_1233_0;
	reg [31:0] b_1234_0;
	reg [31:0] b_1235_0;
	reg [31:0] b_1236_0;
	reg [31:0] b_1237_0;
	reg [31:0] b_1238_0;
	reg [31:0] b_1239_0;
	reg [31:0] b_1240_0;
	reg [31:0] b_1241_0;
	reg [31:0] b_1242_0;
	reg [31:0] b_1243_0;
	reg [31:0] b_1244_0;
	reg [31:0] b_1245_0;
	reg [31:0] b_1246_0;
	reg [31:0] b_1247_0;
	reg [31:0] b_1248_0;
	reg [31:0] b_1249_0;
	reg [31:0] b_1250_0;
	reg [31:0] b_1251_0;
	reg [31:0] b_1252_0;
	reg [31:0] b_1253_0;
	reg [31:0] b_1254_0;
	reg [31:0] b_1255_0;
	reg [31:0] b_1256_0;
	reg [31:0] b_1257_0;
	reg [31:0] b_1258_0;
	reg [31:0] b_1259_0;
	reg [31:0] b_1260_0;
	reg [31:0] b_1261_0;
	reg [31:0] b_1262_0;
	reg [31:0] b_1263_0;
	reg [31:0] b_1264_0;
	reg [31:0] b_1265_0;
	reg [31:0] b_1266_0;
	reg [31:0] b_1267_0;
	reg [31:0] b_1268_0;
	reg [31:0] b_1269_0;
	reg [31:0] b_1270_0;
	reg [31:0] b_1271_0;
	reg [31:0] b_1272_0;
	reg [31:0] b_1273_0;
	reg [31:0] b_1274_0;
	reg [31:0] b_1275_0;
	reg [31:0] b_1276_0;
	reg [31:0] b_1277_0;
	reg [31:0] b_1278_0;
	reg [31:0] b_1279_0;
	reg [31:0] b_1280_0;
	reg [31:0] b_1281_0;
	reg [31:0] b_1282_0;
	reg [31:0] b_1283_0;
	reg [31:0] b_1284_0;
	reg [31:0] b_1285_0;
	reg [31:0] b_1286_0;
	reg [31:0] b_1287_0;
	reg [31:0] b_1288_0;
	reg [31:0] b_1289_0;
	reg [31:0] b_1290_0;
	reg [31:0] b_1291_0;
	reg [31:0] b_1292_0;
	reg [31:0] b_1293_0;
	reg [31:0] b_1294_0;
	reg [31:0] b_1295_0;
	reg [31:0] b_1296_0;
	reg [31:0] b_1297_0;
	reg [31:0] b_1298_0;
	reg [31:0] b_1299_0;
	reg [31:0] b_1300_0;
	reg [31:0] b_1301_0;
	reg [31:0] b_1302_0;
	reg [31:0] b_1303_0;
	reg [31:0] b_1304_0;
	reg [31:0] b_1305_0;
	reg [31:0] b_1306_0;
	reg [31:0] b_1307_0;
	reg [31:0] b_1308_0;
	reg [31:0] b_1309_0;
	reg [31:0] b_1310_0;
	reg [31:0] b_1311_0;
	reg [31:0] b_1312_0;
	reg [31:0] b_1313_0;
	reg [31:0] b_1314_0;
	reg [31:0] b_1315_0;
	reg [31:0] b_1316_0;
	reg [31:0] b_1317_0;
	reg [31:0] b_1318_0;
	reg [31:0] b_1319_0;
	reg [31:0] b_1320_0;
	reg [31:0] b_1321_0;
	reg [31:0] b_1322_0;
	reg [31:0] b_1323_0;
	reg [31:0] b_1324_0;
	reg [31:0] b_1325_0;
	reg [31:0] b_1326_0;
	reg [31:0] b_1327_0;
	reg [31:0] b_1328_0;
	reg [31:0] b_1329_0;
	reg [31:0] b_1330_0;
	reg [31:0] b_1331_0;
	reg [31:0] b_1332_0;
	reg [31:0] b_1333_0;
	reg [31:0] b_1334_0;
	reg [31:0] b_1335_0;
	reg [31:0] b_1336_0;
	reg [31:0] b_1337_0;
	reg [31:0] b_1338_0;
	reg [31:0] b_1339_0;
	reg [31:0] b_1340_0;
	reg [31:0] b_1341_0;
	reg [31:0] b_1342_0;
	reg [31:0] b_1343_0;
	reg [31:0] b_1344_0;
	reg [31:0] b_1345_0;
	reg [31:0] b_1346_0;
	reg [31:0] b_1347_0;
	reg [31:0] b_1348_0;
	reg [31:0] b_1349_0;
	reg [31:0] b_1350_0;
	reg [31:0] b_1351_0;
	reg [31:0] b_1352_0;
	reg [31:0] b_1353_0;
	reg [31:0] b_1354_0;
	reg [31:0] b_1355_0;
	reg [31:0] b_1356_0;
	reg [31:0] b_1357_0;
	reg [31:0] b_1358_0;
	reg [31:0] b_1359_0;
	reg [31:0] b_1360_0;
	reg [31:0] b_1361_0;
	reg [31:0] b_1362_0;
	reg [31:0] b_1363_0;
	reg [31:0] b_1364_0;
	reg [31:0] b_1365_0;
	reg [31:0] b_1366_0;
	reg [31:0] b_1367_0;
	reg [31:0] b_1368_0;
	reg [31:0] b_1369_0;
	reg [31:0] b_1370_0;
	reg [31:0] b_1371_0;
	reg [31:0] b_1372_0;
	reg [31:0] b_1373_0;
	reg [31:0] b_1374_0;
	reg [31:0] b_1375_0;
	reg [31:0] b_1376_0;
	reg [31:0] b_1377_0;
	reg [31:0] b_1378_0;
	reg [31:0] b_1379_0;
	reg [31:0] b_1380_0;
	reg [31:0] b_1381_0;
	reg [31:0] b_1382_0;
	reg [31:0] b_1383_0;
	reg [31:0] b_1384_0;
	reg [31:0] b_1385_0;
	reg [31:0] b_1386_0;
	reg [31:0] b_1387_0;
	reg [31:0] b_1388_0;
	reg [31:0] b_1389_0;
	reg [31:0] b_1390_0;
	reg [31:0] b_1391_0;
	reg [31:0] b_1392_0;
	reg [31:0] b_1393_0;
	reg [31:0] b_1394_0;
	reg [31:0] b_1395_0;
	reg [31:0] b_1396_0;
	reg [31:0] b_1397_0;
	reg [31:0] b_1398_0;
	reg [31:0] b_1399_0;
	reg [31:0] b_1400_0;
	reg [31:0] b_1401_0;
	reg [31:0] b_1402_0;
	reg [31:0] b_1403_0;
	reg [31:0] b_1404_0;
	reg [31:0] b_1405_0;
	reg [31:0] b_1406_0;
	reg [31:0] b_1407_0;
	reg [31:0] b_1408_0;
	reg [31:0] b_1409_0;
	reg [31:0] b_1410_0;
	reg [31:0] b_1411_0;
	reg [31:0] b_1412_0;
	reg [31:0] b_1413_0;
	reg [31:0] b_1414_0;
	reg [31:0] b_1415_0;
	reg [31:0] b_1416_0;
	reg [31:0] b_1417_0;
	reg [31:0] b_1418_0;
	reg [31:0] b_1419_0;
	reg [31:0] b_1420_0;
	reg [31:0] b_1421_0;
	reg [31:0] b_1422_0;
	reg [31:0] b_1423_0;
	reg [31:0] b_1424_0;
	reg [31:0] b_1425_0;
	reg [31:0] b_1426_0;
	reg [31:0] b_1427_0;
	reg [31:0] b_1428_0;
	reg [31:0] b_1429_0;
	reg [31:0] b_1430_0;
	reg [31:0] b_1431_0;
	reg [31:0] b_1432_0;
	reg [31:0] b_1433_0;
	reg [31:0] b_1434_0;
	reg [31:0] b_1435_0;
	reg [31:0] b_1436_0;
	reg [31:0] b_1437_0;
	reg [31:0] b_1438_0;
	reg [31:0] b_1439_0;
	reg [31:0] b_1440_0;
	reg [31:0] b_1441_0;
	reg [31:0] b_1442_0;
	reg [31:0] b_1443_0;
	reg [31:0] b_1444_0;
	reg [31:0] b_1445_0;
	reg [31:0] b_1446_0;
	reg [31:0] b_1447_0;
	reg [31:0] b_1448_0;
	reg [31:0] b_1449_0;
	reg [31:0] b_1450_0;
	reg [31:0] b_1451_0;
	reg [31:0] b_1452_0;
	reg [31:0] b_1453_0;
	reg [31:0] b_1454_0;
	reg [31:0] b_1455_0;
	reg [31:0] b_1456_0;
	reg [31:0] b_1457_0;
	reg [31:0] b_1458_0;
	reg [31:0] b_1459_0;
	reg [31:0] b_1460_0;
	reg [31:0] b_1461_0;
	reg [31:0] b_1462_0;
	reg [31:0] b_1463_0;
	reg [31:0] b_1464_0;
	reg [31:0] b_1465_0;
	reg [31:0] b_1466_0;
	reg [31:0] b_1467_0;
	reg [31:0] b_1468_0;
	reg [31:0] b_1469_0;
	reg [31:0] b_1470_0;
	reg [31:0] b_1471_0;
	reg [31:0] b_1472_0;
	reg [31:0] b_1473_0;
	reg [31:0] b_1474_0;
	reg [31:0] b_1475_0;
	reg [31:0] b_1476_0;
	reg [31:0] b_1477_0;
	reg [31:0] b_1478_0;
	reg [31:0] b_1479_0;
	reg [31:0] b_1480_0;
	reg [31:0] b_1481_0;
	reg [31:0] b_1482_0;
	reg [31:0] b_1483_0;
	reg [31:0] b_1484_0;
	reg [31:0] b_1485_0;
	reg [31:0] b_1486_0;
	reg [31:0] b_1487_0;
	reg [31:0] b_1488_0;
	reg [31:0] b_1489_0;
	reg [31:0] b_1490_0;
	reg [31:0] b_1491_0;
	reg [31:0] b_1492_0;
	reg [31:0] b_1493_0;
	reg [31:0] b_1494_0;
	reg [31:0] b_1495_0;
	reg [31:0] b_1496_0;
	reg [31:0] b_1497_0;
	reg [31:0] b_1498_0;
	reg [31:0] b_1499_0;
	reg [31:0] b_1500_0;
	reg [31:0] b_1501_0;
	reg [31:0] b_1502_0;
	reg [31:0] b_1503_0;
	reg [31:0] b_1504_0;
	reg [31:0] b_1505_0;
	reg [31:0] b_1506_0;
	reg [31:0] b_1507_0;
	reg [31:0] b_1508_0;
	reg [31:0] b_1509_0;
	reg [31:0] b_1510_0;
	reg [31:0] b_1511_0;
	reg [31:0] b_1512_0;
	reg [31:0] b_1513_0;
	reg [31:0] b_1514_0;
	reg [31:0] b_1515_0;
	reg [31:0] b_1516_0;
	reg [31:0] b_1517_0;
	reg [31:0] b_1518_0;
	reg [31:0] b_1519_0;
	reg [31:0] b_1520_0;
	reg [31:0] b_1521_0;
	reg [31:0] b_1522_0;
	reg [31:0] b_1523_0;
	reg [31:0] b_1524_0;
	reg [31:0] b_1525_0;
	reg [31:0] b_1526_0;
	reg [31:0] b_1527_0;
	reg [31:0] b_1528_0;
	reg [31:0] b_1529_0;
	reg [31:0] b_1530_0;
	reg [31:0] b_1531_0;
	reg [31:0] b_1532_0;
	reg [31:0] b_1533_0;
	reg [31:0] b_1534_0;
	reg [31:0] b_1535_0;
	reg [31:0] b_1536_0;
	reg [31:0] b_1537_0;
	reg [31:0] b_1538_0;
	reg [31:0] b_1539_0;
	reg [31:0] b_1540_0;
	reg [31:0] b_1541_0;
	reg [31:0] b_1542_0;
	reg [31:0] b_1543_0;
	reg [31:0] b_1544_0;
	reg [31:0] b_1545_0;
	reg [31:0] b_1546_0;
	reg [31:0] b_1547_0;
	reg [31:0] b_1548_0;
	reg [31:0] b_1549_0;
	reg [31:0] b_1550_0;
	reg [31:0] b_1551_0;
	reg [31:0] b_1552_0;
	reg [31:0] b_1553_0;
	reg [31:0] b_1554_0;
	reg [31:0] b_1555_0;
	reg [31:0] b_1556_0;
	reg [31:0] b_1557_0;
	reg [31:0] b_1558_0;
	reg [31:0] b_1559_0;
	reg [31:0] b_1560_0;
	reg [31:0] b_1561_0;
	reg [31:0] b_1562_0;
	reg [31:0] b_1563_0;
	reg [31:0] b_1564_0;
	reg [31:0] b_1565_0;
	reg [31:0] b_1566_0;
	reg [31:0] b_1567_0;
	reg [31:0] b_1568_0;
	reg [31:0] b_1569_0;
	reg [31:0] b_1570_0;
	reg [31:0] b_1571_0;
	reg [31:0] b_1572_0;
	reg [31:0] b_1573_0;
	reg [31:0] b_1574_0;
	reg [31:0] b_1575_0;
	reg [31:0] b_1576_0;
	reg [31:0] b_1577_0;
	reg [31:0] b_1578_0;
	reg [31:0] b_1579_0;
	reg [31:0] b_1580_0;
	reg [31:0] b_1581_0;
	reg [31:0] b_1582_0;
	reg [31:0] b_1583_0;
	reg [31:0] b_1584_0;
	reg [31:0] b_1585_0;
	reg [31:0] b_1586_0;
	reg [31:0] b_1587_0;
	reg [31:0] b_1588_0;
	reg [31:0] b_1589_0;
	reg [31:0] b_1590_0;
	reg [31:0] b_1591_0;
	reg [31:0] b_1592_0;
	reg [31:0] b_1593_0;
	reg [31:0] b_1594_0;
	reg [31:0] b_1595_0;
	reg [31:0] b_1596_0;
	reg [31:0] b_1597_0;
	reg [31:0] b_1598_0;
	reg [31:0] b_1599_0;
	reg [31:0] b_1600_0;
	reg [31:0] b_1601_0;
	reg [31:0] b_1602_0;
	reg [31:0] b_1603_0;
	reg [31:0] b_1604_0;
	reg [31:0] b_1605_0;
	reg [31:0] b_1606_0;
	reg [31:0] b_1607_0;
	reg [31:0] b_1608_0;
	reg [31:0] b_1609_0;
	reg [31:0] b_1610_0;
	reg [31:0] b_1611_0;
	reg [31:0] b_1612_0;
	reg [31:0] b_1613_0;
	reg [31:0] b_1614_0;
	reg [31:0] b_1615_0;
	reg [31:0] b_1616_0;
	reg [31:0] b_1617_0;
	reg [31:0] b_1618_0;
	reg [31:0] b_1619_0;
	reg [31:0] b_1620_0;
	reg [31:0] b_1621_0;
	reg [31:0] b_1622_0;
	reg [31:0] b_1623_0;
	reg [31:0] b_1624_0;
	reg [31:0] b_1625_0;
	reg [31:0] b_1626_0;
	reg [31:0] b_1627_0;
	reg [31:0] b_1628_0;
	reg [31:0] b_1629_0;
	reg [31:0] b_1630_0;
	reg [31:0] b_1631_0;
	reg [31:0] b_1632_0;
	reg [31:0] b_1633_0;
	reg [31:0] b_1634_0;
	reg [31:0] b_1635_0;
	reg [31:0] b_1636_0;
	reg [31:0] b_1637_0;
	reg [31:0] b_1638_0;
	reg [31:0] b_1639_0;
	reg [31:0] b_1640_0;
	reg [31:0] b_1641_0;
	reg [31:0] b_1642_0;
	reg [31:0] b_1643_0;
	reg [31:0] b_1644_0;
	reg [31:0] b_1645_0;
	reg [31:0] b_1646_0;
	reg [31:0] b_1647_0;
	reg [31:0] b_1648_0;
	reg [31:0] b_1649_0;
	reg [31:0] b_1650_0;
	reg [31:0] b_1651_0;
	reg [31:0] b_1652_0;
	reg [31:0] b_1653_0;
	reg [31:0] b_1654_0;
	reg [31:0] b_1655_0;
	reg [31:0] b_1656_0;
	reg [31:0] b_1657_0;
	reg [31:0] b_1658_0;
	reg [31:0] b_1659_0;
	reg [31:0] b_1660_0;
	reg [31:0] b_1661_0;
	reg [31:0] b_1662_0;
	reg [31:0] b_1663_0;
	reg [31:0] b_1664_0;
	reg [31:0] b_1665_0;
	reg [31:0] b_1666_0;
	reg [31:0] b_1667_0;
	reg [31:0] b_1668_0;
	reg [31:0] b_1669_0;
	reg [31:0] b_1670_0;
	reg [31:0] b_1671_0;
	reg [31:0] b_1672_0;
	reg [31:0] b_1673_0;
	reg [31:0] b_1674_0;
	reg [31:0] b_1675_0;
	reg [31:0] b_1676_0;
	reg [31:0] b_1677_0;
	reg [31:0] b_1678_0;
	reg [31:0] b_1679_0;
	reg [31:0] b_1680_0;
	reg [31:0] b_1681_0;
	reg [31:0] b_1682_0;
	reg [31:0] b_1683_0;
	reg [31:0] b_1684_0;
	reg [31:0] b_1685_0;
	reg [31:0] b_1686_0;
	reg [31:0] b_1687_0;
	reg [31:0] b_1688_0;
	reg [31:0] b_1689_0;
	reg [31:0] b_1690_0;
	reg [31:0] b_1691_0;
	reg [31:0] b_1692_0;
	reg [31:0] b_1693_0;
	reg [31:0] b_1694_0;
	reg [31:0] b_1695_0;
	reg [31:0] b_1696_0;
	reg [31:0] b_1697_0;
	reg [31:0] b_1698_0;
	reg [31:0] b_1699_0;
	reg [31:0] b_1700_0;
	reg [31:0] b_1701_0;
	reg [31:0] b_1702_0;
	reg [31:0] b_1703_0;
	reg [31:0] b_1704_0;
	reg [31:0] b_1705_0;
	reg [31:0] b_1706_0;
	reg [31:0] b_1707_0;
	reg [31:0] b_1708_0;
	reg [31:0] b_1709_0;
	reg [31:0] b_1710_0;
	reg [31:0] b_1711_0;
	reg [31:0] b_1712_0;
	reg [31:0] b_1713_0;
	reg [31:0] b_1714_0;
	reg [31:0] b_1715_0;
	reg [31:0] b_1716_0;
	reg [31:0] b_1717_0;
	reg [31:0] b_1718_0;
	reg [31:0] b_1719_0;
	reg [31:0] b_1720_0;
	reg [31:0] b_1721_0;
	reg [31:0] b_1722_0;
	reg [31:0] b_1723_0;
	reg [31:0] b_1724_0;
	reg [31:0] b_1725_0;
	reg [31:0] b_1726_0;
	reg [31:0] b_1727_0;
	reg [31:0] b_1728_0;
	reg [31:0] b_1729_0;
	reg [31:0] b_1730_0;
	reg [31:0] b_1731_0;
	reg [31:0] b_1732_0;
	reg [31:0] b_1733_0;
	reg [31:0] b_1734_0;
	reg [31:0] b_1735_0;
	reg [31:0] b_1736_0;
	reg [31:0] b_1737_0;
	reg [31:0] b_1738_0;
	reg [31:0] b_1739_0;
	reg [31:0] b_1740_0;
	reg [31:0] b_1741_0;
	reg [31:0] b_1742_0;
	reg [31:0] b_1743_0;
	reg [31:0] b_1744_0;
	reg [31:0] b_1745_0;
	reg [31:0] b_1746_0;
	reg [31:0] b_1747_0;
	reg [31:0] b_1748_0;
	reg [31:0] b_1749_0;
	reg [31:0] b_1750_0;
	reg [31:0] b_1751_0;
	reg [31:0] b_1752_0;
	reg [31:0] b_1753_0;
	reg [31:0] b_1754_0;
	reg [31:0] b_1755_0;
	reg [31:0] b_1756_0;
	reg [31:0] b_1757_0;
	reg [31:0] b_1758_0;
	reg [31:0] b_1759_0;
	reg [31:0] b_1760_0;
	reg [31:0] b_1761_0;
	reg [31:0] b_1762_0;
	reg [31:0] b_1763_0;
	reg [31:0] b_1764_0;
	reg [31:0] b_1765_0;
	reg [31:0] b_1766_0;
	reg [31:0] b_1767_0;
	reg [31:0] b_1768_0;
	reg [31:0] b_1769_0;
	reg [31:0] b_1770_0;
	reg [31:0] b_1771_0;
	reg [31:0] b_1772_0;
	reg [31:0] b_1773_0;
	reg [31:0] b_1774_0;
	reg [31:0] b_1775_0;
	reg [31:0] b_1776_0;
	reg [31:0] b_1777_0;
	reg [31:0] b_1778_0;
	reg [31:0] b_1779_0;
	reg [31:0] b_1780_0;
	reg [31:0] b_1781_0;
	reg [31:0] b_1782_0;
	reg [31:0] b_1783_0;
	reg [31:0] b_1784_0;
	reg [31:0] b_1785_0;
	reg [31:0] b_1786_0;
	reg [31:0] b_1787_0;
	reg [31:0] b_1788_0;
	reg [31:0] b_1789_0;
	reg [31:0] b_1790_0;
	reg [31:0] b_1791_0;
	reg [31:0] b_1792_0;
	reg [31:0] b_1793_0;
	reg [31:0] b_1794_0;
	reg [31:0] b_1795_0;
	reg [31:0] b_1796_0;
	reg [31:0] b_1797_0;
	reg [31:0] b_1798_0;
	reg [31:0] b_1799_0;
	reg [31:0] b_1800_0;
	reg [31:0] b_1801_0;
	reg [31:0] b_1802_0;
	reg [31:0] b_1803_0;
	reg [31:0] b_1804_0;
	reg [31:0] b_1805_0;
	reg [31:0] b_1806_0;
	reg [31:0] b_1807_0;
	reg [31:0] b_1808_0;
	reg [31:0] b_1809_0;
	reg [31:0] b_1810_0;
	reg [31:0] b_1811_0;
	reg [31:0] b_1812_0;
	reg [31:0] b_1813_0;
	reg [31:0] b_1814_0;
	reg [31:0] b_1815_0;
	reg [31:0] b_1816_0;
	reg [31:0] b_1817_0;
	reg [31:0] b_1818_0;
	reg [31:0] b_1819_0;
	reg [31:0] b_1820_0;
	reg [31:0] b_1821_0;
	reg [31:0] b_1822_0;
	reg [31:0] b_1823_0;
	reg [31:0] b_1824_0;
	reg [31:0] b_1825_0;
	reg [31:0] b_1826_0;
	reg [31:0] b_1827_0;
	reg [31:0] b_1828_0;
	reg [31:0] b_1829_0;
	reg [31:0] b_1830_0;
	reg [31:0] b_1831_0;
	reg [31:0] b_1832_0;
	reg [31:0] b_1833_0;
	reg [31:0] b_1834_0;
	reg [31:0] b_1835_0;
	reg [31:0] b_1836_0;
	reg [31:0] b_1837_0;
	reg [31:0] b_1838_0;
	reg [31:0] b_1839_0;
	reg [31:0] b_1840_0;
	reg [31:0] b_1841_0;
	reg [31:0] b_1842_0;
	reg [31:0] b_1843_0;
	reg [31:0] b_1844_0;
	reg [31:0] b_1845_0;
	reg [31:0] b_1846_0;
	reg [31:0] b_1847_0;
	reg [31:0] b_1848_0;
	reg [31:0] b_1849_0;
	reg [31:0] b_1850_0;
	reg [31:0] b_1851_0;
	reg [31:0] b_1852_0;
	reg [31:0] b_1853_0;
	reg [31:0] b_1854_0;
	reg [31:0] b_1855_0;
	reg [31:0] b_1856_0;
	reg [31:0] b_1857_0;
	reg [31:0] b_1858_0;
	reg [31:0] b_1859_0;
	reg [31:0] b_1860_0;
	reg [31:0] b_1861_0;
	reg [31:0] b_1862_0;
	reg [31:0] b_1863_0;
	reg [31:0] b_1864_0;
	reg [31:0] b_1865_0;
	reg [31:0] b_1866_0;
	reg [31:0] b_1867_0;
	reg [31:0] b_1868_0;
	reg [31:0] b_1869_0;
	reg [31:0] b_1870_0;
	reg [31:0] b_1871_0;
	reg [31:0] b_1872_0;
	reg [31:0] b_1873_0;
	reg [31:0] b_1874_0;
	reg [31:0] b_1875_0;
	reg [31:0] b_1876_0;
	reg [31:0] b_1877_0;
	reg [31:0] b_1878_0;
	reg [31:0] b_1879_0;
	reg [31:0] b_1880_0;
	reg [31:0] b_1881_0;
	reg [31:0] b_1882_0;
	reg [31:0] b_1883_0;
	reg [31:0] b_1884_0;
	reg [31:0] b_1885_0;
	reg [31:0] b_1886_0;
	reg [31:0] b_1887_0;
	reg [31:0] b_1888_0;
	reg [31:0] b_1889_0;
	reg [31:0] b_1890_0;
	reg [31:0] b_1891_0;
	reg [31:0] b_1892_0;
	reg [31:0] b_1893_0;
	reg [31:0] b_1894_0;
	reg [31:0] b_1895_0;
	reg [31:0] b_1896_0;
	reg [31:0] b_1897_0;
	reg [31:0] b_1898_0;
	reg [31:0] b_1899_0;
	reg [31:0] b_1900_0;
	reg [31:0] b_1901_0;
	reg [31:0] b_1902_0;
	reg [31:0] b_1903_0;
	reg [31:0] b_1904_0;
	reg [31:0] b_1905_0;
	reg [31:0] b_1906_0;
	reg [31:0] b_1907_0;
	reg [31:0] b_1908_0;
	reg [31:0] b_1909_0;
	reg [31:0] b_1910_0;
	reg [31:0] b_1911_0;
	reg [31:0] b_1912_0;
	reg [31:0] b_1913_0;
	reg [31:0] b_1914_0;
	reg [31:0] b_1915_0;
	reg [31:0] b_1916_0;
	reg [31:0] b_1917_0;
	reg [31:0] b_1918_0;
	reg [31:0] b_1919_0;
	reg [31:0] b_1920_0;
	reg [31:0] b_1921_0;
	reg [31:0] b_1922_0;
	reg [31:0] b_1923_0;
	reg [31:0] b_1924_0;
	reg [31:0] b_1925_0;
	reg [31:0] b_1926_0;
	reg [31:0] b_1927_0;
	reg [31:0] b_1928_0;
	reg [31:0] b_1929_0;
	reg [31:0] b_1930_0;
	reg [31:0] b_1931_0;
	reg [31:0] b_1932_0;
	reg [31:0] b_1933_0;
	reg [31:0] b_1934_0;
	reg [31:0] b_1935_0;
	reg [31:0] b_1936_0;
	reg [31:0] b_1937_0;
	reg [31:0] b_1938_0;
	reg [31:0] b_1939_0;
	reg [31:0] b_1940_0;
	reg [31:0] b_1941_0;
	reg [31:0] b_1942_0;
	reg [31:0] b_1943_0;
	reg [31:0] b_1944_0;
	reg [31:0] b_1945_0;
	reg [31:0] b_1946_0;
	reg [31:0] b_1947_0;
	reg [31:0] b_1948_0;
	reg [31:0] b_1949_0;
	reg [31:0] b_1950_0;
	reg [31:0] b_1951_0;
	reg [31:0] b_1952_0;
	reg [31:0] b_1953_0;
	reg [31:0] b_1954_0;
	reg [31:0] b_1955_0;
	reg [31:0] b_1956_0;
	reg [31:0] b_1957_0;
	reg [31:0] b_1958_0;
	reg [31:0] b_1959_0;
	reg [31:0] b_1960_0;
	reg [31:0] b_1961_0;
	reg [31:0] b_1962_0;
	reg [31:0] b_1963_0;
	reg [31:0] b_1964_0;
	reg [31:0] b_1965_0;
	reg [31:0] b_1966_0;
	reg [31:0] b_1967_0;
	reg [31:0] b_1968_0;
	reg [31:0] b_1969_0;
	reg [31:0] b_1970_0;
	reg [31:0] b_1971_0;
	reg [31:0] b_1972_0;
	reg [31:0] b_1973_0;
	reg [31:0] b_1974_0;
	reg [31:0] b_1975_0;
	reg [31:0] b_1976_0;
	reg [31:0] b_1977_0;
	reg [31:0] b_1978_0;
	reg [31:0] b_1979_0;
	reg [31:0] b_1980_0;
	reg [31:0] b_1981_0;
	reg [31:0] b_1982_0;
	reg [31:0] b_1983_0;
	reg [31:0] b_1984_0;
	reg [31:0] b_1985_0;
	reg [31:0] b_1986_0;
	reg [31:0] b_1987_0;
	reg [31:0] b_1988_0;
	reg [31:0] b_1989_0;
	reg [31:0] b_1990_0;
	reg [31:0] b_1991_0;
	reg [31:0] b_1992_0;
	reg [31:0] b_1993_0;
	reg [31:0] b_1994_0;
	reg [31:0] b_1995_0;
	reg [31:0] b_1996_0;
	reg [31:0] b_1997_0;
	reg [31:0] b_1998_0;
	reg [31:0] b_1999_0;
	reg [31:0] b_2000_0;
	reg [31:0] b_2001_0;
	reg [31:0] b_2002_0;
	reg [31:0] b_2003_0;
	reg [31:0] b_2004_0;
	reg [31:0] b_2005_0;
	reg [31:0] b_2006_0;
	reg [31:0] b_2007_0;
	reg [31:0] b_2008_0;
	reg [31:0] b_2009_0;
	reg [31:0] b_2010_0;
	reg [31:0] b_2011_0;
	reg [31:0] b_2012_0;
	reg [31:0] b_2013_0;
	reg [31:0] b_2014_0;
	reg [31:0] b_2015_0;
	reg [31:0] b_2016_0;
	reg [31:0] b_2017_0;
	reg [31:0] b_2018_0;
	reg [31:0] b_2019_0;
	reg [31:0] b_2020_0;
	reg [31:0] b_2021_0;
	reg [31:0] b_2022_0;
	reg [31:0] b_2023_0;
	reg [31:0] b_2024_0;
	reg [31:0] b_2025_0;
	reg [31:0] b_2026_0;
	reg [31:0] b_2027_0;
	reg [31:0] b_2028_0;
	reg [31:0] b_2029_0;
	reg [31:0] b_2030_0;
	reg [31:0] b_2031_0;
	reg [31:0] b_2032_0;
	reg [31:0] b_2033_0;
	reg [31:0] b_2034_0;
	reg [31:0] b_2035_0;
	reg [31:0] b_2036_0;
	reg [31:0] b_2037_0;
	reg [31:0] b_2038_0;
	reg [31:0] b_2039_0;
	reg [31:0] b_2040_0;
	reg [31:0] b_2041_0;
	reg [31:0] b_2042_0;
	reg [31:0] b_2043_0;
	reg [31:0] b_2044_0;
	reg [31:0] b_2045_0;
	reg [31:0] b_2046_0;
	reg [31:0] b_2047_0;
	reg [4:0] mesh_0_0_io_in_control_0_shift_b;
	reg mesh_0_0_io_in_control_0_dataflow_b;
	reg mesh_0_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_0_io_in_control_0_shift_b;
	reg mesh_1_0_io_in_control_0_dataflow_b;
	reg mesh_1_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_0_io_in_control_0_shift_b;
	reg mesh_2_0_io_in_control_0_dataflow_b;
	reg mesh_2_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_0_io_in_control_0_shift_b;
	reg mesh_3_0_io_in_control_0_dataflow_b;
	reg mesh_3_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_0_io_in_control_0_shift_b;
	reg mesh_4_0_io_in_control_0_dataflow_b;
	reg mesh_4_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_0_io_in_control_0_shift_b;
	reg mesh_5_0_io_in_control_0_dataflow_b;
	reg mesh_5_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_0_io_in_control_0_shift_b;
	reg mesh_6_0_io_in_control_0_dataflow_b;
	reg mesh_6_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_0_io_in_control_0_shift_b;
	reg mesh_7_0_io_in_control_0_dataflow_b;
	reg mesh_7_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_0_io_in_control_0_shift_b;
	reg mesh_8_0_io_in_control_0_dataflow_b;
	reg mesh_8_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_0_io_in_control_0_shift_b;
	reg mesh_9_0_io_in_control_0_dataflow_b;
	reg mesh_9_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_0_io_in_control_0_shift_b;
	reg mesh_10_0_io_in_control_0_dataflow_b;
	reg mesh_10_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_0_io_in_control_0_shift_b;
	reg mesh_11_0_io_in_control_0_dataflow_b;
	reg mesh_11_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_0_io_in_control_0_shift_b;
	reg mesh_12_0_io_in_control_0_dataflow_b;
	reg mesh_12_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_0_io_in_control_0_shift_b;
	reg mesh_13_0_io_in_control_0_dataflow_b;
	reg mesh_13_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_0_io_in_control_0_shift_b;
	reg mesh_14_0_io_in_control_0_dataflow_b;
	reg mesh_14_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_0_io_in_control_0_shift_b;
	reg mesh_15_0_io_in_control_0_dataflow_b;
	reg mesh_15_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_0_io_in_control_0_shift_b;
	reg mesh_16_0_io_in_control_0_dataflow_b;
	reg mesh_16_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_0_io_in_control_0_shift_b;
	reg mesh_17_0_io_in_control_0_dataflow_b;
	reg mesh_17_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_0_io_in_control_0_shift_b;
	reg mesh_18_0_io_in_control_0_dataflow_b;
	reg mesh_18_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_0_io_in_control_0_shift_b;
	reg mesh_19_0_io_in_control_0_dataflow_b;
	reg mesh_19_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_0_io_in_control_0_shift_b;
	reg mesh_20_0_io_in_control_0_dataflow_b;
	reg mesh_20_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_0_io_in_control_0_shift_b;
	reg mesh_21_0_io_in_control_0_dataflow_b;
	reg mesh_21_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_0_io_in_control_0_shift_b;
	reg mesh_22_0_io_in_control_0_dataflow_b;
	reg mesh_22_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_0_io_in_control_0_shift_b;
	reg mesh_23_0_io_in_control_0_dataflow_b;
	reg mesh_23_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_0_io_in_control_0_shift_b;
	reg mesh_24_0_io_in_control_0_dataflow_b;
	reg mesh_24_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_0_io_in_control_0_shift_b;
	reg mesh_25_0_io_in_control_0_dataflow_b;
	reg mesh_25_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_0_io_in_control_0_shift_b;
	reg mesh_26_0_io_in_control_0_dataflow_b;
	reg mesh_26_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_0_io_in_control_0_shift_b;
	reg mesh_27_0_io_in_control_0_dataflow_b;
	reg mesh_27_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_0_io_in_control_0_shift_b;
	reg mesh_28_0_io_in_control_0_dataflow_b;
	reg mesh_28_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_0_io_in_control_0_shift_b;
	reg mesh_29_0_io_in_control_0_dataflow_b;
	reg mesh_29_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_0_io_in_control_0_shift_b;
	reg mesh_30_0_io_in_control_0_dataflow_b;
	reg mesh_30_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_0_io_in_control_0_shift_b;
	reg mesh_31_0_io_in_control_0_dataflow_b;
	reg mesh_31_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_1_io_in_control_0_shift_b;
	reg mesh_0_1_io_in_control_0_dataflow_b;
	reg mesh_0_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_1_io_in_control_0_shift_b;
	reg mesh_1_1_io_in_control_0_dataflow_b;
	reg mesh_1_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_1_io_in_control_0_shift_b;
	reg mesh_2_1_io_in_control_0_dataflow_b;
	reg mesh_2_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_1_io_in_control_0_shift_b;
	reg mesh_3_1_io_in_control_0_dataflow_b;
	reg mesh_3_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_1_io_in_control_0_shift_b;
	reg mesh_4_1_io_in_control_0_dataflow_b;
	reg mesh_4_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_1_io_in_control_0_shift_b;
	reg mesh_5_1_io_in_control_0_dataflow_b;
	reg mesh_5_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_1_io_in_control_0_shift_b;
	reg mesh_6_1_io_in_control_0_dataflow_b;
	reg mesh_6_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_1_io_in_control_0_shift_b;
	reg mesh_7_1_io_in_control_0_dataflow_b;
	reg mesh_7_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_1_io_in_control_0_shift_b;
	reg mesh_8_1_io_in_control_0_dataflow_b;
	reg mesh_8_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_1_io_in_control_0_shift_b;
	reg mesh_9_1_io_in_control_0_dataflow_b;
	reg mesh_9_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_1_io_in_control_0_shift_b;
	reg mesh_10_1_io_in_control_0_dataflow_b;
	reg mesh_10_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_1_io_in_control_0_shift_b;
	reg mesh_11_1_io_in_control_0_dataflow_b;
	reg mesh_11_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_1_io_in_control_0_shift_b;
	reg mesh_12_1_io_in_control_0_dataflow_b;
	reg mesh_12_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_1_io_in_control_0_shift_b;
	reg mesh_13_1_io_in_control_0_dataflow_b;
	reg mesh_13_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_1_io_in_control_0_shift_b;
	reg mesh_14_1_io_in_control_0_dataflow_b;
	reg mesh_14_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_1_io_in_control_0_shift_b;
	reg mesh_15_1_io_in_control_0_dataflow_b;
	reg mesh_15_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_1_io_in_control_0_shift_b;
	reg mesh_16_1_io_in_control_0_dataflow_b;
	reg mesh_16_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_1_io_in_control_0_shift_b;
	reg mesh_17_1_io_in_control_0_dataflow_b;
	reg mesh_17_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_1_io_in_control_0_shift_b;
	reg mesh_18_1_io_in_control_0_dataflow_b;
	reg mesh_18_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_1_io_in_control_0_shift_b;
	reg mesh_19_1_io_in_control_0_dataflow_b;
	reg mesh_19_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_1_io_in_control_0_shift_b;
	reg mesh_20_1_io_in_control_0_dataflow_b;
	reg mesh_20_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_1_io_in_control_0_shift_b;
	reg mesh_21_1_io_in_control_0_dataflow_b;
	reg mesh_21_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_1_io_in_control_0_shift_b;
	reg mesh_22_1_io_in_control_0_dataflow_b;
	reg mesh_22_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_1_io_in_control_0_shift_b;
	reg mesh_23_1_io_in_control_0_dataflow_b;
	reg mesh_23_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_1_io_in_control_0_shift_b;
	reg mesh_24_1_io_in_control_0_dataflow_b;
	reg mesh_24_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_1_io_in_control_0_shift_b;
	reg mesh_25_1_io_in_control_0_dataflow_b;
	reg mesh_25_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_1_io_in_control_0_shift_b;
	reg mesh_26_1_io_in_control_0_dataflow_b;
	reg mesh_26_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_1_io_in_control_0_shift_b;
	reg mesh_27_1_io_in_control_0_dataflow_b;
	reg mesh_27_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_1_io_in_control_0_shift_b;
	reg mesh_28_1_io_in_control_0_dataflow_b;
	reg mesh_28_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_1_io_in_control_0_shift_b;
	reg mesh_29_1_io_in_control_0_dataflow_b;
	reg mesh_29_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_1_io_in_control_0_shift_b;
	reg mesh_30_1_io_in_control_0_dataflow_b;
	reg mesh_30_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_1_io_in_control_0_shift_b;
	reg mesh_31_1_io_in_control_0_dataflow_b;
	reg mesh_31_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_2_io_in_control_0_shift_b;
	reg mesh_0_2_io_in_control_0_dataflow_b;
	reg mesh_0_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_2_io_in_control_0_shift_b;
	reg mesh_1_2_io_in_control_0_dataflow_b;
	reg mesh_1_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_2_io_in_control_0_shift_b;
	reg mesh_2_2_io_in_control_0_dataflow_b;
	reg mesh_2_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_2_io_in_control_0_shift_b;
	reg mesh_3_2_io_in_control_0_dataflow_b;
	reg mesh_3_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_2_io_in_control_0_shift_b;
	reg mesh_4_2_io_in_control_0_dataflow_b;
	reg mesh_4_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_2_io_in_control_0_shift_b;
	reg mesh_5_2_io_in_control_0_dataflow_b;
	reg mesh_5_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_2_io_in_control_0_shift_b;
	reg mesh_6_2_io_in_control_0_dataflow_b;
	reg mesh_6_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_2_io_in_control_0_shift_b;
	reg mesh_7_2_io_in_control_0_dataflow_b;
	reg mesh_7_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_2_io_in_control_0_shift_b;
	reg mesh_8_2_io_in_control_0_dataflow_b;
	reg mesh_8_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_2_io_in_control_0_shift_b;
	reg mesh_9_2_io_in_control_0_dataflow_b;
	reg mesh_9_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_2_io_in_control_0_shift_b;
	reg mesh_10_2_io_in_control_0_dataflow_b;
	reg mesh_10_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_2_io_in_control_0_shift_b;
	reg mesh_11_2_io_in_control_0_dataflow_b;
	reg mesh_11_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_2_io_in_control_0_shift_b;
	reg mesh_12_2_io_in_control_0_dataflow_b;
	reg mesh_12_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_2_io_in_control_0_shift_b;
	reg mesh_13_2_io_in_control_0_dataflow_b;
	reg mesh_13_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_2_io_in_control_0_shift_b;
	reg mesh_14_2_io_in_control_0_dataflow_b;
	reg mesh_14_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_2_io_in_control_0_shift_b;
	reg mesh_15_2_io_in_control_0_dataflow_b;
	reg mesh_15_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_2_io_in_control_0_shift_b;
	reg mesh_16_2_io_in_control_0_dataflow_b;
	reg mesh_16_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_2_io_in_control_0_shift_b;
	reg mesh_17_2_io_in_control_0_dataflow_b;
	reg mesh_17_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_2_io_in_control_0_shift_b;
	reg mesh_18_2_io_in_control_0_dataflow_b;
	reg mesh_18_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_2_io_in_control_0_shift_b;
	reg mesh_19_2_io_in_control_0_dataflow_b;
	reg mesh_19_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_2_io_in_control_0_shift_b;
	reg mesh_20_2_io_in_control_0_dataflow_b;
	reg mesh_20_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_2_io_in_control_0_shift_b;
	reg mesh_21_2_io_in_control_0_dataflow_b;
	reg mesh_21_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_2_io_in_control_0_shift_b;
	reg mesh_22_2_io_in_control_0_dataflow_b;
	reg mesh_22_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_2_io_in_control_0_shift_b;
	reg mesh_23_2_io_in_control_0_dataflow_b;
	reg mesh_23_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_2_io_in_control_0_shift_b;
	reg mesh_24_2_io_in_control_0_dataflow_b;
	reg mesh_24_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_2_io_in_control_0_shift_b;
	reg mesh_25_2_io_in_control_0_dataflow_b;
	reg mesh_25_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_2_io_in_control_0_shift_b;
	reg mesh_26_2_io_in_control_0_dataflow_b;
	reg mesh_26_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_2_io_in_control_0_shift_b;
	reg mesh_27_2_io_in_control_0_dataflow_b;
	reg mesh_27_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_2_io_in_control_0_shift_b;
	reg mesh_28_2_io_in_control_0_dataflow_b;
	reg mesh_28_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_2_io_in_control_0_shift_b;
	reg mesh_29_2_io_in_control_0_dataflow_b;
	reg mesh_29_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_2_io_in_control_0_shift_b;
	reg mesh_30_2_io_in_control_0_dataflow_b;
	reg mesh_30_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_2_io_in_control_0_shift_b;
	reg mesh_31_2_io_in_control_0_dataflow_b;
	reg mesh_31_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_3_io_in_control_0_shift_b;
	reg mesh_0_3_io_in_control_0_dataflow_b;
	reg mesh_0_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_3_io_in_control_0_shift_b;
	reg mesh_1_3_io_in_control_0_dataflow_b;
	reg mesh_1_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_3_io_in_control_0_shift_b;
	reg mesh_2_3_io_in_control_0_dataflow_b;
	reg mesh_2_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_3_io_in_control_0_shift_b;
	reg mesh_3_3_io_in_control_0_dataflow_b;
	reg mesh_3_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_3_io_in_control_0_shift_b;
	reg mesh_4_3_io_in_control_0_dataflow_b;
	reg mesh_4_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_3_io_in_control_0_shift_b;
	reg mesh_5_3_io_in_control_0_dataflow_b;
	reg mesh_5_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_3_io_in_control_0_shift_b;
	reg mesh_6_3_io_in_control_0_dataflow_b;
	reg mesh_6_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_3_io_in_control_0_shift_b;
	reg mesh_7_3_io_in_control_0_dataflow_b;
	reg mesh_7_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_3_io_in_control_0_shift_b;
	reg mesh_8_3_io_in_control_0_dataflow_b;
	reg mesh_8_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_3_io_in_control_0_shift_b;
	reg mesh_9_3_io_in_control_0_dataflow_b;
	reg mesh_9_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_3_io_in_control_0_shift_b;
	reg mesh_10_3_io_in_control_0_dataflow_b;
	reg mesh_10_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_3_io_in_control_0_shift_b;
	reg mesh_11_3_io_in_control_0_dataflow_b;
	reg mesh_11_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_3_io_in_control_0_shift_b;
	reg mesh_12_3_io_in_control_0_dataflow_b;
	reg mesh_12_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_3_io_in_control_0_shift_b;
	reg mesh_13_3_io_in_control_0_dataflow_b;
	reg mesh_13_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_3_io_in_control_0_shift_b;
	reg mesh_14_3_io_in_control_0_dataflow_b;
	reg mesh_14_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_3_io_in_control_0_shift_b;
	reg mesh_15_3_io_in_control_0_dataflow_b;
	reg mesh_15_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_3_io_in_control_0_shift_b;
	reg mesh_16_3_io_in_control_0_dataflow_b;
	reg mesh_16_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_3_io_in_control_0_shift_b;
	reg mesh_17_3_io_in_control_0_dataflow_b;
	reg mesh_17_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_3_io_in_control_0_shift_b;
	reg mesh_18_3_io_in_control_0_dataflow_b;
	reg mesh_18_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_3_io_in_control_0_shift_b;
	reg mesh_19_3_io_in_control_0_dataflow_b;
	reg mesh_19_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_3_io_in_control_0_shift_b;
	reg mesh_20_3_io_in_control_0_dataflow_b;
	reg mesh_20_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_3_io_in_control_0_shift_b;
	reg mesh_21_3_io_in_control_0_dataflow_b;
	reg mesh_21_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_3_io_in_control_0_shift_b;
	reg mesh_22_3_io_in_control_0_dataflow_b;
	reg mesh_22_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_3_io_in_control_0_shift_b;
	reg mesh_23_3_io_in_control_0_dataflow_b;
	reg mesh_23_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_3_io_in_control_0_shift_b;
	reg mesh_24_3_io_in_control_0_dataflow_b;
	reg mesh_24_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_3_io_in_control_0_shift_b;
	reg mesh_25_3_io_in_control_0_dataflow_b;
	reg mesh_25_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_3_io_in_control_0_shift_b;
	reg mesh_26_3_io_in_control_0_dataflow_b;
	reg mesh_26_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_3_io_in_control_0_shift_b;
	reg mesh_27_3_io_in_control_0_dataflow_b;
	reg mesh_27_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_3_io_in_control_0_shift_b;
	reg mesh_28_3_io_in_control_0_dataflow_b;
	reg mesh_28_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_3_io_in_control_0_shift_b;
	reg mesh_29_3_io_in_control_0_dataflow_b;
	reg mesh_29_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_3_io_in_control_0_shift_b;
	reg mesh_30_3_io_in_control_0_dataflow_b;
	reg mesh_30_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_3_io_in_control_0_shift_b;
	reg mesh_31_3_io_in_control_0_dataflow_b;
	reg mesh_31_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_4_io_in_control_0_shift_b;
	reg mesh_0_4_io_in_control_0_dataflow_b;
	reg mesh_0_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_4_io_in_control_0_shift_b;
	reg mesh_1_4_io_in_control_0_dataflow_b;
	reg mesh_1_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_4_io_in_control_0_shift_b;
	reg mesh_2_4_io_in_control_0_dataflow_b;
	reg mesh_2_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_4_io_in_control_0_shift_b;
	reg mesh_3_4_io_in_control_0_dataflow_b;
	reg mesh_3_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_4_io_in_control_0_shift_b;
	reg mesh_4_4_io_in_control_0_dataflow_b;
	reg mesh_4_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_4_io_in_control_0_shift_b;
	reg mesh_5_4_io_in_control_0_dataflow_b;
	reg mesh_5_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_4_io_in_control_0_shift_b;
	reg mesh_6_4_io_in_control_0_dataflow_b;
	reg mesh_6_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_4_io_in_control_0_shift_b;
	reg mesh_7_4_io_in_control_0_dataflow_b;
	reg mesh_7_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_4_io_in_control_0_shift_b;
	reg mesh_8_4_io_in_control_0_dataflow_b;
	reg mesh_8_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_4_io_in_control_0_shift_b;
	reg mesh_9_4_io_in_control_0_dataflow_b;
	reg mesh_9_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_4_io_in_control_0_shift_b;
	reg mesh_10_4_io_in_control_0_dataflow_b;
	reg mesh_10_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_4_io_in_control_0_shift_b;
	reg mesh_11_4_io_in_control_0_dataflow_b;
	reg mesh_11_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_4_io_in_control_0_shift_b;
	reg mesh_12_4_io_in_control_0_dataflow_b;
	reg mesh_12_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_4_io_in_control_0_shift_b;
	reg mesh_13_4_io_in_control_0_dataflow_b;
	reg mesh_13_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_4_io_in_control_0_shift_b;
	reg mesh_14_4_io_in_control_0_dataflow_b;
	reg mesh_14_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_4_io_in_control_0_shift_b;
	reg mesh_15_4_io_in_control_0_dataflow_b;
	reg mesh_15_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_4_io_in_control_0_shift_b;
	reg mesh_16_4_io_in_control_0_dataflow_b;
	reg mesh_16_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_4_io_in_control_0_shift_b;
	reg mesh_17_4_io_in_control_0_dataflow_b;
	reg mesh_17_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_4_io_in_control_0_shift_b;
	reg mesh_18_4_io_in_control_0_dataflow_b;
	reg mesh_18_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_4_io_in_control_0_shift_b;
	reg mesh_19_4_io_in_control_0_dataflow_b;
	reg mesh_19_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_4_io_in_control_0_shift_b;
	reg mesh_20_4_io_in_control_0_dataflow_b;
	reg mesh_20_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_4_io_in_control_0_shift_b;
	reg mesh_21_4_io_in_control_0_dataflow_b;
	reg mesh_21_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_4_io_in_control_0_shift_b;
	reg mesh_22_4_io_in_control_0_dataflow_b;
	reg mesh_22_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_4_io_in_control_0_shift_b;
	reg mesh_23_4_io_in_control_0_dataflow_b;
	reg mesh_23_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_4_io_in_control_0_shift_b;
	reg mesh_24_4_io_in_control_0_dataflow_b;
	reg mesh_24_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_4_io_in_control_0_shift_b;
	reg mesh_25_4_io_in_control_0_dataflow_b;
	reg mesh_25_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_4_io_in_control_0_shift_b;
	reg mesh_26_4_io_in_control_0_dataflow_b;
	reg mesh_26_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_4_io_in_control_0_shift_b;
	reg mesh_27_4_io_in_control_0_dataflow_b;
	reg mesh_27_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_4_io_in_control_0_shift_b;
	reg mesh_28_4_io_in_control_0_dataflow_b;
	reg mesh_28_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_4_io_in_control_0_shift_b;
	reg mesh_29_4_io_in_control_0_dataflow_b;
	reg mesh_29_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_4_io_in_control_0_shift_b;
	reg mesh_30_4_io_in_control_0_dataflow_b;
	reg mesh_30_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_4_io_in_control_0_shift_b;
	reg mesh_31_4_io_in_control_0_dataflow_b;
	reg mesh_31_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_5_io_in_control_0_shift_b;
	reg mesh_0_5_io_in_control_0_dataflow_b;
	reg mesh_0_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_5_io_in_control_0_shift_b;
	reg mesh_1_5_io_in_control_0_dataflow_b;
	reg mesh_1_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_5_io_in_control_0_shift_b;
	reg mesh_2_5_io_in_control_0_dataflow_b;
	reg mesh_2_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_5_io_in_control_0_shift_b;
	reg mesh_3_5_io_in_control_0_dataflow_b;
	reg mesh_3_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_5_io_in_control_0_shift_b;
	reg mesh_4_5_io_in_control_0_dataflow_b;
	reg mesh_4_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_5_io_in_control_0_shift_b;
	reg mesh_5_5_io_in_control_0_dataflow_b;
	reg mesh_5_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_5_io_in_control_0_shift_b;
	reg mesh_6_5_io_in_control_0_dataflow_b;
	reg mesh_6_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_5_io_in_control_0_shift_b;
	reg mesh_7_5_io_in_control_0_dataflow_b;
	reg mesh_7_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_5_io_in_control_0_shift_b;
	reg mesh_8_5_io_in_control_0_dataflow_b;
	reg mesh_8_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_5_io_in_control_0_shift_b;
	reg mesh_9_5_io_in_control_0_dataflow_b;
	reg mesh_9_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_5_io_in_control_0_shift_b;
	reg mesh_10_5_io_in_control_0_dataflow_b;
	reg mesh_10_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_5_io_in_control_0_shift_b;
	reg mesh_11_5_io_in_control_0_dataflow_b;
	reg mesh_11_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_5_io_in_control_0_shift_b;
	reg mesh_12_5_io_in_control_0_dataflow_b;
	reg mesh_12_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_5_io_in_control_0_shift_b;
	reg mesh_13_5_io_in_control_0_dataflow_b;
	reg mesh_13_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_5_io_in_control_0_shift_b;
	reg mesh_14_5_io_in_control_0_dataflow_b;
	reg mesh_14_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_5_io_in_control_0_shift_b;
	reg mesh_15_5_io_in_control_0_dataflow_b;
	reg mesh_15_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_5_io_in_control_0_shift_b;
	reg mesh_16_5_io_in_control_0_dataflow_b;
	reg mesh_16_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_5_io_in_control_0_shift_b;
	reg mesh_17_5_io_in_control_0_dataflow_b;
	reg mesh_17_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_5_io_in_control_0_shift_b;
	reg mesh_18_5_io_in_control_0_dataflow_b;
	reg mesh_18_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_5_io_in_control_0_shift_b;
	reg mesh_19_5_io_in_control_0_dataflow_b;
	reg mesh_19_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_5_io_in_control_0_shift_b;
	reg mesh_20_5_io_in_control_0_dataflow_b;
	reg mesh_20_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_5_io_in_control_0_shift_b;
	reg mesh_21_5_io_in_control_0_dataflow_b;
	reg mesh_21_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_5_io_in_control_0_shift_b;
	reg mesh_22_5_io_in_control_0_dataflow_b;
	reg mesh_22_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_5_io_in_control_0_shift_b;
	reg mesh_23_5_io_in_control_0_dataflow_b;
	reg mesh_23_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_5_io_in_control_0_shift_b;
	reg mesh_24_5_io_in_control_0_dataflow_b;
	reg mesh_24_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_5_io_in_control_0_shift_b;
	reg mesh_25_5_io_in_control_0_dataflow_b;
	reg mesh_25_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_5_io_in_control_0_shift_b;
	reg mesh_26_5_io_in_control_0_dataflow_b;
	reg mesh_26_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_5_io_in_control_0_shift_b;
	reg mesh_27_5_io_in_control_0_dataflow_b;
	reg mesh_27_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_5_io_in_control_0_shift_b;
	reg mesh_28_5_io_in_control_0_dataflow_b;
	reg mesh_28_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_5_io_in_control_0_shift_b;
	reg mesh_29_5_io_in_control_0_dataflow_b;
	reg mesh_29_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_5_io_in_control_0_shift_b;
	reg mesh_30_5_io_in_control_0_dataflow_b;
	reg mesh_30_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_5_io_in_control_0_shift_b;
	reg mesh_31_5_io_in_control_0_dataflow_b;
	reg mesh_31_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_6_io_in_control_0_shift_b;
	reg mesh_0_6_io_in_control_0_dataflow_b;
	reg mesh_0_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_6_io_in_control_0_shift_b;
	reg mesh_1_6_io_in_control_0_dataflow_b;
	reg mesh_1_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_6_io_in_control_0_shift_b;
	reg mesh_2_6_io_in_control_0_dataflow_b;
	reg mesh_2_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_6_io_in_control_0_shift_b;
	reg mesh_3_6_io_in_control_0_dataflow_b;
	reg mesh_3_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_6_io_in_control_0_shift_b;
	reg mesh_4_6_io_in_control_0_dataflow_b;
	reg mesh_4_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_6_io_in_control_0_shift_b;
	reg mesh_5_6_io_in_control_0_dataflow_b;
	reg mesh_5_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_6_io_in_control_0_shift_b;
	reg mesh_6_6_io_in_control_0_dataflow_b;
	reg mesh_6_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_6_io_in_control_0_shift_b;
	reg mesh_7_6_io_in_control_0_dataflow_b;
	reg mesh_7_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_6_io_in_control_0_shift_b;
	reg mesh_8_6_io_in_control_0_dataflow_b;
	reg mesh_8_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_6_io_in_control_0_shift_b;
	reg mesh_9_6_io_in_control_0_dataflow_b;
	reg mesh_9_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_6_io_in_control_0_shift_b;
	reg mesh_10_6_io_in_control_0_dataflow_b;
	reg mesh_10_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_6_io_in_control_0_shift_b;
	reg mesh_11_6_io_in_control_0_dataflow_b;
	reg mesh_11_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_6_io_in_control_0_shift_b;
	reg mesh_12_6_io_in_control_0_dataflow_b;
	reg mesh_12_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_6_io_in_control_0_shift_b;
	reg mesh_13_6_io_in_control_0_dataflow_b;
	reg mesh_13_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_6_io_in_control_0_shift_b;
	reg mesh_14_6_io_in_control_0_dataflow_b;
	reg mesh_14_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_6_io_in_control_0_shift_b;
	reg mesh_15_6_io_in_control_0_dataflow_b;
	reg mesh_15_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_6_io_in_control_0_shift_b;
	reg mesh_16_6_io_in_control_0_dataflow_b;
	reg mesh_16_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_6_io_in_control_0_shift_b;
	reg mesh_17_6_io_in_control_0_dataflow_b;
	reg mesh_17_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_6_io_in_control_0_shift_b;
	reg mesh_18_6_io_in_control_0_dataflow_b;
	reg mesh_18_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_6_io_in_control_0_shift_b;
	reg mesh_19_6_io_in_control_0_dataflow_b;
	reg mesh_19_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_6_io_in_control_0_shift_b;
	reg mesh_20_6_io_in_control_0_dataflow_b;
	reg mesh_20_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_6_io_in_control_0_shift_b;
	reg mesh_21_6_io_in_control_0_dataflow_b;
	reg mesh_21_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_6_io_in_control_0_shift_b;
	reg mesh_22_6_io_in_control_0_dataflow_b;
	reg mesh_22_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_6_io_in_control_0_shift_b;
	reg mesh_23_6_io_in_control_0_dataflow_b;
	reg mesh_23_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_6_io_in_control_0_shift_b;
	reg mesh_24_6_io_in_control_0_dataflow_b;
	reg mesh_24_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_6_io_in_control_0_shift_b;
	reg mesh_25_6_io_in_control_0_dataflow_b;
	reg mesh_25_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_6_io_in_control_0_shift_b;
	reg mesh_26_6_io_in_control_0_dataflow_b;
	reg mesh_26_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_6_io_in_control_0_shift_b;
	reg mesh_27_6_io_in_control_0_dataflow_b;
	reg mesh_27_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_6_io_in_control_0_shift_b;
	reg mesh_28_6_io_in_control_0_dataflow_b;
	reg mesh_28_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_6_io_in_control_0_shift_b;
	reg mesh_29_6_io_in_control_0_dataflow_b;
	reg mesh_29_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_6_io_in_control_0_shift_b;
	reg mesh_30_6_io_in_control_0_dataflow_b;
	reg mesh_30_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_6_io_in_control_0_shift_b;
	reg mesh_31_6_io_in_control_0_dataflow_b;
	reg mesh_31_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_7_io_in_control_0_shift_b;
	reg mesh_0_7_io_in_control_0_dataflow_b;
	reg mesh_0_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_7_io_in_control_0_shift_b;
	reg mesh_1_7_io_in_control_0_dataflow_b;
	reg mesh_1_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_7_io_in_control_0_shift_b;
	reg mesh_2_7_io_in_control_0_dataflow_b;
	reg mesh_2_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_7_io_in_control_0_shift_b;
	reg mesh_3_7_io_in_control_0_dataflow_b;
	reg mesh_3_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_7_io_in_control_0_shift_b;
	reg mesh_4_7_io_in_control_0_dataflow_b;
	reg mesh_4_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_7_io_in_control_0_shift_b;
	reg mesh_5_7_io_in_control_0_dataflow_b;
	reg mesh_5_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_7_io_in_control_0_shift_b;
	reg mesh_6_7_io_in_control_0_dataflow_b;
	reg mesh_6_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_7_io_in_control_0_shift_b;
	reg mesh_7_7_io_in_control_0_dataflow_b;
	reg mesh_7_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_7_io_in_control_0_shift_b;
	reg mesh_8_7_io_in_control_0_dataflow_b;
	reg mesh_8_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_7_io_in_control_0_shift_b;
	reg mesh_9_7_io_in_control_0_dataflow_b;
	reg mesh_9_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_7_io_in_control_0_shift_b;
	reg mesh_10_7_io_in_control_0_dataflow_b;
	reg mesh_10_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_7_io_in_control_0_shift_b;
	reg mesh_11_7_io_in_control_0_dataflow_b;
	reg mesh_11_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_7_io_in_control_0_shift_b;
	reg mesh_12_7_io_in_control_0_dataflow_b;
	reg mesh_12_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_7_io_in_control_0_shift_b;
	reg mesh_13_7_io_in_control_0_dataflow_b;
	reg mesh_13_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_7_io_in_control_0_shift_b;
	reg mesh_14_7_io_in_control_0_dataflow_b;
	reg mesh_14_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_7_io_in_control_0_shift_b;
	reg mesh_15_7_io_in_control_0_dataflow_b;
	reg mesh_15_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_7_io_in_control_0_shift_b;
	reg mesh_16_7_io_in_control_0_dataflow_b;
	reg mesh_16_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_7_io_in_control_0_shift_b;
	reg mesh_17_7_io_in_control_0_dataflow_b;
	reg mesh_17_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_7_io_in_control_0_shift_b;
	reg mesh_18_7_io_in_control_0_dataflow_b;
	reg mesh_18_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_7_io_in_control_0_shift_b;
	reg mesh_19_7_io_in_control_0_dataflow_b;
	reg mesh_19_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_7_io_in_control_0_shift_b;
	reg mesh_20_7_io_in_control_0_dataflow_b;
	reg mesh_20_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_7_io_in_control_0_shift_b;
	reg mesh_21_7_io_in_control_0_dataflow_b;
	reg mesh_21_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_7_io_in_control_0_shift_b;
	reg mesh_22_7_io_in_control_0_dataflow_b;
	reg mesh_22_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_7_io_in_control_0_shift_b;
	reg mesh_23_7_io_in_control_0_dataflow_b;
	reg mesh_23_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_7_io_in_control_0_shift_b;
	reg mesh_24_7_io_in_control_0_dataflow_b;
	reg mesh_24_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_7_io_in_control_0_shift_b;
	reg mesh_25_7_io_in_control_0_dataflow_b;
	reg mesh_25_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_7_io_in_control_0_shift_b;
	reg mesh_26_7_io_in_control_0_dataflow_b;
	reg mesh_26_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_7_io_in_control_0_shift_b;
	reg mesh_27_7_io_in_control_0_dataflow_b;
	reg mesh_27_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_7_io_in_control_0_shift_b;
	reg mesh_28_7_io_in_control_0_dataflow_b;
	reg mesh_28_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_7_io_in_control_0_shift_b;
	reg mesh_29_7_io_in_control_0_dataflow_b;
	reg mesh_29_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_7_io_in_control_0_shift_b;
	reg mesh_30_7_io_in_control_0_dataflow_b;
	reg mesh_30_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_7_io_in_control_0_shift_b;
	reg mesh_31_7_io_in_control_0_dataflow_b;
	reg mesh_31_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_8_io_in_control_0_shift_b;
	reg mesh_0_8_io_in_control_0_dataflow_b;
	reg mesh_0_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_8_io_in_control_0_shift_b;
	reg mesh_1_8_io_in_control_0_dataflow_b;
	reg mesh_1_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_8_io_in_control_0_shift_b;
	reg mesh_2_8_io_in_control_0_dataflow_b;
	reg mesh_2_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_8_io_in_control_0_shift_b;
	reg mesh_3_8_io_in_control_0_dataflow_b;
	reg mesh_3_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_8_io_in_control_0_shift_b;
	reg mesh_4_8_io_in_control_0_dataflow_b;
	reg mesh_4_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_8_io_in_control_0_shift_b;
	reg mesh_5_8_io_in_control_0_dataflow_b;
	reg mesh_5_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_8_io_in_control_0_shift_b;
	reg mesh_6_8_io_in_control_0_dataflow_b;
	reg mesh_6_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_8_io_in_control_0_shift_b;
	reg mesh_7_8_io_in_control_0_dataflow_b;
	reg mesh_7_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_8_io_in_control_0_shift_b;
	reg mesh_8_8_io_in_control_0_dataflow_b;
	reg mesh_8_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_8_io_in_control_0_shift_b;
	reg mesh_9_8_io_in_control_0_dataflow_b;
	reg mesh_9_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_8_io_in_control_0_shift_b;
	reg mesh_10_8_io_in_control_0_dataflow_b;
	reg mesh_10_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_8_io_in_control_0_shift_b;
	reg mesh_11_8_io_in_control_0_dataflow_b;
	reg mesh_11_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_8_io_in_control_0_shift_b;
	reg mesh_12_8_io_in_control_0_dataflow_b;
	reg mesh_12_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_8_io_in_control_0_shift_b;
	reg mesh_13_8_io_in_control_0_dataflow_b;
	reg mesh_13_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_8_io_in_control_0_shift_b;
	reg mesh_14_8_io_in_control_0_dataflow_b;
	reg mesh_14_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_8_io_in_control_0_shift_b;
	reg mesh_15_8_io_in_control_0_dataflow_b;
	reg mesh_15_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_8_io_in_control_0_shift_b;
	reg mesh_16_8_io_in_control_0_dataflow_b;
	reg mesh_16_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_8_io_in_control_0_shift_b;
	reg mesh_17_8_io_in_control_0_dataflow_b;
	reg mesh_17_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_8_io_in_control_0_shift_b;
	reg mesh_18_8_io_in_control_0_dataflow_b;
	reg mesh_18_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_8_io_in_control_0_shift_b;
	reg mesh_19_8_io_in_control_0_dataflow_b;
	reg mesh_19_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_8_io_in_control_0_shift_b;
	reg mesh_20_8_io_in_control_0_dataflow_b;
	reg mesh_20_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_8_io_in_control_0_shift_b;
	reg mesh_21_8_io_in_control_0_dataflow_b;
	reg mesh_21_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_8_io_in_control_0_shift_b;
	reg mesh_22_8_io_in_control_0_dataflow_b;
	reg mesh_22_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_8_io_in_control_0_shift_b;
	reg mesh_23_8_io_in_control_0_dataflow_b;
	reg mesh_23_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_8_io_in_control_0_shift_b;
	reg mesh_24_8_io_in_control_0_dataflow_b;
	reg mesh_24_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_8_io_in_control_0_shift_b;
	reg mesh_25_8_io_in_control_0_dataflow_b;
	reg mesh_25_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_8_io_in_control_0_shift_b;
	reg mesh_26_8_io_in_control_0_dataflow_b;
	reg mesh_26_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_8_io_in_control_0_shift_b;
	reg mesh_27_8_io_in_control_0_dataflow_b;
	reg mesh_27_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_8_io_in_control_0_shift_b;
	reg mesh_28_8_io_in_control_0_dataflow_b;
	reg mesh_28_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_8_io_in_control_0_shift_b;
	reg mesh_29_8_io_in_control_0_dataflow_b;
	reg mesh_29_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_8_io_in_control_0_shift_b;
	reg mesh_30_8_io_in_control_0_dataflow_b;
	reg mesh_30_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_8_io_in_control_0_shift_b;
	reg mesh_31_8_io_in_control_0_dataflow_b;
	reg mesh_31_8_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_9_io_in_control_0_shift_b;
	reg mesh_0_9_io_in_control_0_dataflow_b;
	reg mesh_0_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_9_io_in_control_0_shift_b;
	reg mesh_1_9_io_in_control_0_dataflow_b;
	reg mesh_1_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_9_io_in_control_0_shift_b;
	reg mesh_2_9_io_in_control_0_dataflow_b;
	reg mesh_2_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_9_io_in_control_0_shift_b;
	reg mesh_3_9_io_in_control_0_dataflow_b;
	reg mesh_3_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_9_io_in_control_0_shift_b;
	reg mesh_4_9_io_in_control_0_dataflow_b;
	reg mesh_4_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_9_io_in_control_0_shift_b;
	reg mesh_5_9_io_in_control_0_dataflow_b;
	reg mesh_5_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_9_io_in_control_0_shift_b;
	reg mesh_6_9_io_in_control_0_dataflow_b;
	reg mesh_6_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_9_io_in_control_0_shift_b;
	reg mesh_7_9_io_in_control_0_dataflow_b;
	reg mesh_7_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_9_io_in_control_0_shift_b;
	reg mesh_8_9_io_in_control_0_dataflow_b;
	reg mesh_8_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_9_io_in_control_0_shift_b;
	reg mesh_9_9_io_in_control_0_dataflow_b;
	reg mesh_9_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_9_io_in_control_0_shift_b;
	reg mesh_10_9_io_in_control_0_dataflow_b;
	reg mesh_10_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_9_io_in_control_0_shift_b;
	reg mesh_11_9_io_in_control_0_dataflow_b;
	reg mesh_11_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_9_io_in_control_0_shift_b;
	reg mesh_12_9_io_in_control_0_dataflow_b;
	reg mesh_12_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_9_io_in_control_0_shift_b;
	reg mesh_13_9_io_in_control_0_dataflow_b;
	reg mesh_13_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_9_io_in_control_0_shift_b;
	reg mesh_14_9_io_in_control_0_dataflow_b;
	reg mesh_14_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_9_io_in_control_0_shift_b;
	reg mesh_15_9_io_in_control_0_dataflow_b;
	reg mesh_15_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_9_io_in_control_0_shift_b;
	reg mesh_16_9_io_in_control_0_dataflow_b;
	reg mesh_16_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_9_io_in_control_0_shift_b;
	reg mesh_17_9_io_in_control_0_dataflow_b;
	reg mesh_17_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_9_io_in_control_0_shift_b;
	reg mesh_18_9_io_in_control_0_dataflow_b;
	reg mesh_18_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_9_io_in_control_0_shift_b;
	reg mesh_19_9_io_in_control_0_dataflow_b;
	reg mesh_19_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_9_io_in_control_0_shift_b;
	reg mesh_20_9_io_in_control_0_dataflow_b;
	reg mesh_20_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_9_io_in_control_0_shift_b;
	reg mesh_21_9_io_in_control_0_dataflow_b;
	reg mesh_21_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_9_io_in_control_0_shift_b;
	reg mesh_22_9_io_in_control_0_dataflow_b;
	reg mesh_22_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_9_io_in_control_0_shift_b;
	reg mesh_23_9_io_in_control_0_dataflow_b;
	reg mesh_23_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_9_io_in_control_0_shift_b;
	reg mesh_24_9_io_in_control_0_dataflow_b;
	reg mesh_24_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_9_io_in_control_0_shift_b;
	reg mesh_25_9_io_in_control_0_dataflow_b;
	reg mesh_25_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_9_io_in_control_0_shift_b;
	reg mesh_26_9_io_in_control_0_dataflow_b;
	reg mesh_26_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_9_io_in_control_0_shift_b;
	reg mesh_27_9_io_in_control_0_dataflow_b;
	reg mesh_27_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_9_io_in_control_0_shift_b;
	reg mesh_28_9_io_in_control_0_dataflow_b;
	reg mesh_28_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_9_io_in_control_0_shift_b;
	reg mesh_29_9_io_in_control_0_dataflow_b;
	reg mesh_29_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_9_io_in_control_0_shift_b;
	reg mesh_30_9_io_in_control_0_dataflow_b;
	reg mesh_30_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_9_io_in_control_0_shift_b;
	reg mesh_31_9_io_in_control_0_dataflow_b;
	reg mesh_31_9_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_10_io_in_control_0_shift_b;
	reg mesh_0_10_io_in_control_0_dataflow_b;
	reg mesh_0_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_10_io_in_control_0_shift_b;
	reg mesh_1_10_io_in_control_0_dataflow_b;
	reg mesh_1_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_10_io_in_control_0_shift_b;
	reg mesh_2_10_io_in_control_0_dataflow_b;
	reg mesh_2_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_10_io_in_control_0_shift_b;
	reg mesh_3_10_io_in_control_0_dataflow_b;
	reg mesh_3_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_10_io_in_control_0_shift_b;
	reg mesh_4_10_io_in_control_0_dataflow_b;
	reg mesh_4_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_10_io_in_control_0_shift_b;
	reg mesh_5_10_io_in_control_0_dataflow_b;
	reg mesh_5_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_10_io_in_control_0_shift_b;
	reg mesh_6_10_io_in_control_0_dataflow_b;
	reg mesh_6_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_10_io_in_control_0_shift_b;
	reg mesh_7_10_io_in_control_0_dataflow_b;
	reg mesh_7_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_10_io_in_control_0_shift_b;
	reg mesh_8_10_io_in_control_0_dataflow_b;
	reg mesh_8_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_10_io_in_control_0_shift_b;
	reg mesh_9_10_io_in_control_0_dataflow_b;
	reg mesh_9_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_10_io_in_control_0_shift_b;
	reg mesh_10_10_io_in_control_0_dataflow_b;
	reg mesh_10_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_10_io_in_control_0_shift_b;
	reg mesh_11_10_io_in_control_0_dataflow_b;
	reg mesh_11_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_10_io_in_control_0_shift_b;
	reg mesh_12_10_io_in_control_0_dataflow_b;
	reg mesh_12_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_10_io_in_control_0_shift_b;
	reg mesh_13_10_io_in_control_0_dataflow_b;
	reg mesh_13_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_10_io_in_control_0_shift_b;
	reg mesh_14_10_io_in_control_0_dataflow_b;
	reg mesh_14_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_10_io_in_control_0_shift_b;
	reg mesh_15_10_io_in_control_0_dataflow_b;
	reg mesh_15_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_10_io_in_control_0_shift_b;
	reg mesh_16_10_io_in_control_0_dataflow_b;
	reg mesh_16_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_10_io_in_control_0_shift_b;
	reg mesh_17_10_io_in_control_0_dataflow_b;
	reg mesh_17_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_10_io_in_control_0_shift_b;
	reg mesh_18_10_io_in_control_0_dataflow_b;
	reg mesh_18_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_10_io_in_control_0_shift_b;
	reg mesh_19_10_io_in_control_0_dataflow_b;
	reg mesh_19_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_10_io_in_control_0_shift_b;
	reg mesh_20_10_io_in_control_0_dataflow_b;
	reg mesh_20_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_10_io_in_control_0_shift_b;
	reg mesh_21_10_io_in_control_0_dataflow_b;
	reg mesh_21_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_10_io_in_control_0_shift_b;
	reg mesh_22_10_io_in_control_0_dataflow_b;
	reg mesh_22_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_10_io_in_control_0_shift_b;
	reg mesh_23_10_io_in_control_0_dataflow_b;
	reg mesh_23_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_10_io_in_control_0_shift_b;
	reg mesh_24_10_io_in_control_0_dataflow_b;
	reg mesh_24_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_10_io_in_control_0_shift_b;
	reg mesh_25_10_io_in_control_0_dataflow_b;
	reg mesh_25_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_10_io_in_control_0_shift_b;
	reg mesh_26_10_io_in_control_0_dataflow_b;
	reg mesh_26_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_10_io_in_control_0_shift_b;
	reg mesh_27_10_io_in_control_0_dataflow_b;
	reg mesh_27_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_10_io_in_control_0_shift_b;
	reg mesh_28_10_io_in_control_0_dataflow_b;
	reg mesh_28_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_10_io_in_control_0_shift_b;
	reg mesh_29_10_io_in_control_0_dataflow_b;
	reg mesh_29_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_10_io_in_control_0_shift_b;
	reg mesh_30_10_io_in_control_0_dataflow_b;
	reg mesh_30_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_10_io_in_control_0_shift_b;
	reg mesh_31_10_io_in_control_0_dataflow_b;
	reg mesh_31_10_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_11_io_in_control_0_shift_b;
	reg mesh_0_11_io_in_control_0_dataflow_b;
	reg mesh_0_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_11_io_in_control_0_shift_b;
	reg mesh_1_11_io_in_control_0_dataflow_b;
	reg mesh_1_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_11_io_in_control_0_shift_b;
	reg mesh_2_11_io_in_control_0_dataflow_b;
	reg mesh_2_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_11_io_in_control_0_shift_b;
	reg mesh_3_11_io_in_control_0_dataflow_b;
	reg mesh_3_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_11_io_in_control_0_shift_b;
	reg mesh_4_11_io_in_control_0_dataflow_b;
	reg mesh_4_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_11_io_in_control_0_shift_b;
	reg mesh_5_11_io_in_control_0_dataflow_b;
	reg mesh_5_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_11_io_in_control_0_shift_b;
	reg mesh_6_11_io_in_control_0_dataflow_b;
	reg mesh_6_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_11_io_in_control_0_shift_b;
	reg mesh_7_11_io_in_control_0_dataflow_b;
	reg mesh_7_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_11_io_in_control_0_shift_b;
	reg mesh_8_11_io_in_control_0_dataflow_b;
	reg mesh_8_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_11_io_in_control_0_shift_b;
	reg mesh_9_11_io_in_control_0_dataflow_b;
	reg mesh_9_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_11_io_in_control_0_shift_b;
	reg mesh_10_11_io_in_control_0_dataflow_b;
	reg mesh_10_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_11_io_in_control_0_shift_b;
	reg mesh_11_11_io_in_control_0_dataflow_b;
	reg mesh_11_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_11_io_in_control_0_shift_b;
	reg mesh_12_11_io_in_control_0_dataflow_b;
	reg mesh_12_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_11_io_in_control_0_shift_b;
	reg mesh_13_11_io_in_control_0_dataflow_b;
	reg mesh_13_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_11_io_in_control_0_shift_b;
	reg mesh_14_11_io_in_control_0_dataflow_b;
	reg mesh_14_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_11_io_in_control_0_shift_b;
	reg mesh_15_11_io_in_control_0_dataflow_b;
	reg mesh_15_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_11_io_in_control_0_shift_b;
	reg mesh_16_11_io_in_control_0_dataflow_b;
	reg mesh_16_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_11_io_in_control_0_shift_b;
	reg mesh_17_11_io_in_control_0_dataflow_b;
	reg mesh_17_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_11_io_in_control_0_shift_b;
	reg mesh_18_11_io_in_control_0_dataflow_b;
	reg mesh_18_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_11_io_in_control_0_shift_b;
	reg mesh_19_11_io_in_control_0_dataflow_b;
	reg mesh_19_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_11_io_in_control_0_shift_b;
	reg mesh_20_11_io_in_control_0_dataflow_b;
	reg mesh_20_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_11_io_in_control_0_shift_b;
	reg mesh_21_11_io_in_control_0_dataflow_b;
	reg mesh_21_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_11_io_in_control_0_shift_b;
	reg mesh_22_11_io_in_control_0_dataflow_b;
	reg mesh_22_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_11_io_in_control_0_shift_b;
	reg mesh_23_11_io_in_control_0_dataflow_b;
	reg mesh_23_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_11_io_in_control_0_shift_b;
	reg mesh_24_11_io_in_control_0_dataflow_b;
	reg mesh_24_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_11_io_in_control_0_shift_b;
	reg mesh_25_11_io_in_control_0_dataflow_b;
	reg mesh_25_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_11_io_in_control_0_shift_b;
	reg mesh_26_11_io_in_control_0_dataflow_b;
	reg mesh_26_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_11_io_in_control_0_shift_b;
	reg mesh_27_11_io_in_control_0_dataflow_b;
	reg mesh_27_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_11_io_in_control_0_shift_b;
	reg mesh_28_11_io_in_control_0_dataflow_b;
	reg mesh_28_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_11_io_in_control_0_shift_b;
	reg mesh_29_11_io_in_control_0_dataflow_b;
	reg mesh_29_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_11_io_in_control_0_shift_b;
	reg mesh_30_11_io_in_control_0_dataflow_b;
	reg mesh_30_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_11_io_in_control_0_shift_b;
	reg mesh_31_11_io_in_control_0_dataflow_b;
	reg mesh_31_11_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_12_io_in_control_0_shift_b;
	reg mesh_0_12_io_in_control_0_dataflow_b;
	reg mesh_0_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_12_io_in_control_0_shift_b;
	reg mesh_1_12_io_in_control_0_dataflow_b;
	reg mesh_1_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_12_io_in_control_0_shift_b;
	reg mesh_2_12_io_in_control_0_dataflow_b;
	reg mesh_2_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_12_io_in_control_0_shift_b;
	reg mesh_3_12_io_in_control_0_dataflow_b;
	reg mesh_3_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_12_io_in_control_0_shift_b;
	reg mesh_4_12_io_in_control_0_dataflow_b;
	reg mesh_4_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_12_io_in_control_0_shift_b;
	reg mesh_5_12_io_in_control_0_dataflow_b;
	reg mesh_5_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_12_io_in_control_0_shift_b;
	reg mesh_6_12_io_in_control_0_dataflow_b;
	reg mesh_6_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_12_io_in_control_0_shift_b;
	reg mesh_7_12_io_in_control_0_dataflow_b;
	reg mesh_7_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_12_io_in_control_0_shift_b;
	reg mesh_8_12_io_in_control_0_dataflow_b;
	reg mesh_8_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_12_io_in_control_0_shift_b;
	reg mesh_9_12_io_in_control_0_dataflow_b;
	reg mesh_9_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_12_io_in_control_0_shift_b;
	reg mesh_10_12_io_in_control_0_dataflow_b;
	reg mesh_10_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_12_io_in_control_0_shift_b;
	reg mesh_11_12_io_in_control_0_dataflow_b;
	reg mesh_11_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_12_io_in_control_0_shift_b;
	reg mesh_12_12_io_in_control_0_dataflow_b;
	reg mesh_12_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_12_io_in_control_0_shift_b;
	reg mesh_13_12_io_in_control_0_dataflow_b;
	reg mesh_13_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_12_io_in_control_0_shift_b;
	reg mesh_14_12_io_in_control_0_dataflow_b;
	reg mesh_14_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_12_io_in_control_0_shift_b;
	reg mesh_15_12_io_in_control_0_dataflow_b;
	reg mesh_15_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_12_io_in_control_0_shift_b;
	reg mesh_16_12_io_in_control_0_dataflow_b;
	reg mesh_16_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_12_io_in_control_0_shift_b;
	reg mesh_17_12_io_in_control_0_dataflow_b;
	reg mesh_17_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_12_io_in_control_0_shift_b;
	reg mesh_18_12_io_in_control_0_dataflow_b;
	reg mesh_18_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_12_io_in_control_0_shift_b;
	reg mesh_19_12_io_in_control_0_dataflow_b;
	reg mesh_19_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_12_io_in_control_0_shift_b;
	reg mesh_20_12_io_in_control_0_dataflow_b;
	reg mesh_20_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_12_io_in_control_0_shift_b;
	reg mesh_21_12_io_in_control_0_dataflow_b;
	reg mesh_21_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_12_io_in_control_0_shift_b;
	reg mesh_22_12_io_in_control_0_dataflow_b;
	reg mesh_22_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_12_io_in_control_0_shift_b;
	reg mesh_23_12_io_in_control_0_dataflow_b;
	reg mesh_23_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_12_io_in_control_0_shift_b;
	reg mesh_24_12_io_in_control_0_dataflow_b;
	reg mesh_24_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_12_io_in_control_0_shift_b;
	reg mesh_25_12_io_in_control_0_dataflow_b;
	reg mesh_25_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_12_io_in_control_0_shift_b;
	reg mesh_26_12_io_in_control_0_dataflow_b;
	reg mesh_26_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_12_io_in_control_0_shift_b;
	reg mesh_27_12_io_in_control_0_dataflow_b;
	reg mesh_27_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_12_io_in_control_0_shift_b;
	reg mesh_28_12_io_in_control_0_dataflow_b;
	reg mesh_28_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_12_io_in_control_0_shift_b;
	reg mesh_29_12_io_in_control_0_dataflow_b;
	reg mesh_29_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_12_io_in_control_0_shift_b;
	reg mesh_30_12_io_in_control_0_dataflow_b;
	reg mesh_30_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_12_io_in_control_0_shift_b;
	reg mesh_31_12_io_in_control_0_dataflow_b;
	reg mesh_31_12_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_13_io_in_control_0_shift_b;
	reg mesh_0_13_io_in_control_0_dataflow_b;
	reg mesh_0_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_13_io_in_control_0_shift_b;
	reg mesh_1_13_io_in_control_0_dataflow_b;
	reg mesh_1_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_13_io_in_control_0_shift_b;
	reg mesh_2_13_io_in_control_0_dataflow_b;
	reg mesh_2_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_13_io_in_control_0_shift_b;
	reg mesh_3_13_io_in_control_0_dataflow_b;
	reg mesh_3_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_13_io_in_control_0_shift_b;
	reg mesh_4_13_io_in_control_0_dataflow_b;
	reg mesh_4_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_13_io_in_control_0_shift_b;
	reg mesh_5_13_io_in_control_0_dataflow_b;
	reg mesh_5_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_13_io_in_control_0_shift_b;
	reg mesh_6_13_io_in_control_0_dataflow_b;
	reg mesh_6_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_13_io_in_control_0_shift_b;
	reg mesh_7_13_io_in_control_0_dataflow_b;
	reg mesh_7_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_13_io_in_control_0_shift_b;
	reg mesh_8_13_io_in_control_0_dataflow_b;
	reg mesh_8_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_13_io_in_control_0_shift_b;
	reg mesh_9_13_io_in_control_0_dataflow_b;
	reg mesh_9_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_13_io_in_control_0_shift_b;
	reg mesh_10_13_io_in_control_0_dataflow_b;
	reg mesh_10_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_13_io_in_control_0_shift_b;
	reg mesh_11_13_io_in_control_0_dataflow_b;
	reg mesh_11_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_13_io_in_control_0_shift_b;
	reg mesh_12_13_io_in_control_0_dataflow_b;
	reg mesh_12_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_13_io_in_control_0_shift_b;
	reg mesh_13_13_io_in_control_0_dataflow_b;
	reg mesh_13_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_13_io_in_control_0_shift_b;
	reg mesh_14_13_io_in_control_0_dataflow_b;
	reg mesh_14_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_13_io_in_control_0_shift_b;
	reg mesh_15_13_io_in_control_0_dataflow_b;
	reg mesh_15_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_13_io_in_control_0_shift_b;
	reg mesh_16_13_io_in_control_0_dataflow_b;
	reg mesh_16_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_13_io_in_control_0_shift_b;
	reg mesh_17_13_io_in_control_0_dataflow_b;
	reg mesh_17_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_13_io_in_control_0_shift_b;
	reg mesh_18_13_io_in_control_0_dataflow_b;
	reg mesh_18_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_13_io_in_control_0_shift_b;
	reg mesh_19_13_io_in_control_0_dataflow_b;
	reg mesh_19_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_13_io_in_control_0_shift_b;
	reg mesh_20_13_io_in_control_0_dataflow_b;
	reg mesh_20_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_13_io_in_control_0_shift_b;
	reg mesh_21_13_io_in_control_0_dataflow_b;
	reg mesh_21_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_13_io_in_control_0_shift_b;
	reg mesh_22_13_io_in_control_0_dataflow_b;
	reg mesh_22_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_13_io_in_control_0_shift_b;
	reg mesh_23_13_io_in_control_0_dataflow_b;
	reg mesh_23_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_13_io_in_control_0_shift_b;
	reg mesh_24_13_io_in_control_0_dataflow_b;
	reg mesh_24_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_13_io_in_control_0_shift_b;
	reg mesh_25_13_io_in_control_0_dataflow_b;
	reg mesh_25_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_13_io_in_control_0_shift_b;
	reg mesh_26_13_io_in_control_0_dataflow_b;
	reg mesh_26_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_13_io_in_control_0_shift_b;
	reg mesh_27_13_io_in_control_0_dataflow_b;
	reg mesh_27_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_13_io_in_control_0_shift_b;
	reg mesh_28_13_io_in_control_0_dataflow_b;
	reg mesh_28_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_13_io_in_control_0_shift_b;
	reg mesh_29_13_io_in_control_0_dataflow_b;
	reg mesh_29_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_13_io_in_control_0_shift_b;
	reg mesh_30_13_io_in_control_0_dataflow_b;
	reg mesh_30_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_13_io_in_control_0_shift_b;
	reg mesh_31_13_io_in_control_0_dataflow_b;
	reg mesh_31_13_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_14_io_in_control_0_shift_b;
	reg mesh_0_14_io_in_control_0_dataflow_b;
	reg mesh_0_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_14_io_in_control_0_shift_b;
	reg mesh_1_14_io_in_control_0_dataflow_b;
	reg mesh_1_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_14_io_in_control_0_shift_b;
	reg mesh_2_14_io_in_control_0_dataflow_b;
	reg mesh_2_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_14_io_in_control_0_shift_b;
	reg mesh_3_14_io_in_control_0_dataflow_b;
	reg mesh_3_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_14_io_in_control_0_shift_b;
	reg mesh_4_14_io_in_control_0_dataflow_b;
	reg mesh_4_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_14_io_in_control_0_shift_b;
	reg mesh_5_14_io_in_control_0_dataflow_b;
	reg mesh_5_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_14_io_in_control_0_shift_b;
	reg mesh_6_14_io_in_control_0_dataflow_b;
	reg mesh_6_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_14_io_in_control_0_shift_b;
	reg mesh_7_14_io_in_control_0_dataflow_b;
	reg mesh_7_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_14_io_in_control_0_shift_b;
	reg mesh_8_14_io_in_control_0_dataflow_b;
	reg mesh_8_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_14_io_in_control_0_shift_b;
	reg mesh_9_14_io_in_control_0_dataflow_b;
	reg mesh_9_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_14_io_in_control_0_shift_b;
	reg mesh_10_14_io_in_control_0_dataflow_b;
	reg mesh_10_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_14_io_in_control_0_shift_b;
	reg mesh_11_14_io_in_control_0_dataflow_b;
	reg mesh_11_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_14_io_in_control_0_shift_b;
	reg mesh_12_14_io_in_control_0_dataflow_b;
	reg mesh_12_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_14_io_in_control_0_shift_b;
	reg mesh_13_14_io_in_control_0_dataflow_b;
	reg mesh_13_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_14_io_in_control_0_shift_b;
	reg mesh_14_14_io_in_control_0_dataflow_b;
	reg mesh_14_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_14_io_in_control_0_shift_b;
	reg mesh_15_14_io_in_control_0_dataflow_b;
	reg mesh_15_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_14_io_in_control_0_shift_b;
	reg mesh_16_14_io_in_control_0_dataflow_b;
	reg mesh_16_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_14_io_in_control_0_shift_b;
	reg mesh_17_14_io_in_control_0_dataflow_b;
	reg mesh_17_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_14_io_in_control_0_shift_b;
	reg mesh_18_14_io_in_control_0_dataflow_b;
	reg mesh_18_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_14_io_in_control_0_shift_b;
	reg mesh_19_14_io_in_control_0_dataflow_b;
	reg mesh_19_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_14_io_in_control_0_shift_b;
	reg mesh_20_14_io_in_control_0_dataflow_b;
	reg mesh_20_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_14_io_in_control_0_shift_b;
	reg mesh_21_14_io_in_control_0_dataflow_b;
	reg mesh_21_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_14_io_in_control_0_shift_b;
	reg mesh_22_14_io_in_control_0_dataflow_b;
	reg mesh_22_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_14_io_in_control_0_shift_b;
	reg mesh_23_14_io_in_control_0_dataflow_b;
	reg mesh_23_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_14_io_in_control_0_shift_b;
	reg mesh_24_14_io_in_control_0_dataflow_b;
	reg mesh_24_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_14_io_in_control_0_shift_b;
	reg mesh_25_14_io_in_control_0_dataflow_b;
	reg mesh_25_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_14_io_in_control_0_shift_b;
	reg mesh_26_14_io_in_control_0_dataflow_b;
	reg mesh_26_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_14_io_in_control_0_shift_b;
	reg mesh_27_14_io_in_control_0_dataflow_b;
	reg mesh_27_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_14_io_in_control_0_shift_b;
	reg mesh_28_14_io_in_control_0_dataflow_b;
	reg mesh_28_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_14_io_in_control_0_shift_b;
	reg mesh_29_14_io_in_control_0_dataflow_b;
	reg mesh_29_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_14_io_in_control_0_shift_b;
	reg mesh_30_14_io_in_control_0_dataflow_b;
	reg mesh_30_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_14_io_in_control_0_shift_b;
	reg mesh_31_14_io_in_control_0_dataflow_b;
	reg mesh_31_14_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_15_io_in_control_0_shift_b;
	reg mesh_0_15_io_in_control_0_dataflow_b;
	reg mesh_0_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_15_io_in_control_0_shift_b;
	reg mesh_1_15_io_in_control_0_dataflow_b;
	reg mesh_1_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_15_io_in_control_0_shift_b;
	reg mesh_2_15_io_in_control_0_dataflow_b;
	reg mesh_2_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_15_io_in_control_0_shift_b;
	reg mesh_3_15_io_in_control_0_dataflow_b;
	reg mesh_3_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_15_io_in_control_0_shift_b;
	reg mesh_4_15_io_in_control_0_dataflow_b;
	reg mesh_4_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_15_io_in_control_0_shift_b;
	reg mesh_5_15_io_in_control_0_dataflow_b;
	reg mesh_5_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_15_io_in_control_0_shift_b;
	reg mesh_6_15_io_in_control_0_dataflow_b;
	reg mesh_6_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_15_io_in_control_0_shift_b;
	reg mesh_7_15_io_in_control_0_dataflow_b;
	reg mesh_7_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_15_io_in_control_0_shift_b;
	reg mesh_8_15_io_in_control_0_dataflow_b;
	reg mesh_8_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_15_io_in_control_0_shift_b;
	reg mesh_9_15_io_in_control_0_dataflow_b;
	reg mesh_9_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_15_io_in_control_0_shift_b;
	reg mesh_10_15_io_in_control_0_dataflow_b;
	reg mesh_10_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_15_io_in_control_0_shift_b;
	reg mesh_11_15_io_in_control_0_dataflow_b;
	reg mesh_11_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_15_io_in_control_0_shift_b;
	reg mesh_12_15_io_in_control_0_dataflow_b;
	reg mesh_12_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_15_io_in_control_0_shift_b;
	reg mesh_13_15_io_in_control_0_dataflow_b;
	reg mesh_13_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_15_io_in_control_0_shift_b;
	reg mesh_14_15_io_in_control_0_dataflow_b;
	reg mesh_14_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_15_io_in_control_0_shift_b;
	reg mesh_15_15_io_in_control_0_dataflow_b;
	reg mesh_15_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_15_io_in_control_0_shift_b;
	reg mesh_16_15_io_in_control_0_dataflow_b;
	reg mesh_16_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_15_io_in_control_0_shift_b;
	reg mesh_17_15_io_in_control_0_dataflow_b;
	reg mesh_17_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_15_io_in_control_0_shift_b;
	reg mesh_18_15_io_in_control_0_dataflow_b;
	reg mesh_18_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_15_io_in_control_0_shift_b;
	reg mesh_19_15_io_in_control_0_dataflow_b;
	reg mesh_19_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_15_io_in_control_0_shift_b;
	reg mesh_20_15_io_in_control_0_dataflow_b;
	reg mesh_20_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_15_io_in_control_0_shift_b;
	reg mesh_21_15_io_in_control_0_dataflow_b;
	reg mesh_21_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_15_io_in_control_0_shift_b;
	reg mesh_22_15_io_in_control_0_dataflow_b;
	reg mesh_22_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_15_io_in_control_0_shift_b;
	reg mesh_23_15_io_in_control_0_dataflow_b;
	reg mesh_23_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_15_io_in_control_0_shift_b;
	reg mesh_24_15_io_in_control_0_dataflow_b;
	reg mesh_24_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_15_io_in_control_0_shift_b;
	reg mesh_25_15_io_in_control_0_dataflow_b;
	reg mesh_25_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_15_io_in_control_0_shift_b;
	reg mesh_26_15_io_in_control_0_dataflow_b;
	reg mesh_26_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_15_io_in_control_0_shift_b;
	reg mesh_27_15_io_in_control_0_dataflow_b;
	reg mesh_27_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_15_io_in_control_0_shift_b;
	reg mesh_28_15_io_in_control_0_dataflow_b;
	reg mesh_28_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_15_io_in_control_0_shift_b;
	reg mesh_29_15_io_in_control_0_dataflow_b;
	reg mesh_29_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_15_io_in_control_0_shift_b;
	reg mesh_30_15_io_in_control_0_dataflow_b;
	reg mesh_30_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_15_io_in_control_0_shift_b;
	reg mesh_31_15_io_in_control_0_dataflow_b;
	reg mesh_31_15_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_16_io_in_control_0_shift_b;
	reg mesh_0_16_io_in_control_0_dataflow_b;
	reg mesh_0_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_16_io_in_control_0_shift_b;
	reg mesh_1_16_io_in_control_0_dataflow_b;
	reg mesh_1_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_16_io_in_control_0_shift_b;
	reg mesh_2_16_io_in_control_0_dataflow_b;
	reg mesh_2_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_16_io_in_control_0_shift_b;
	reg mesh_3_16_io_in_control_0_dataflow_b;
	reg mesh_3_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_16_io_in_control_0_shift_b;
	reg mesh_4_16_io_in_control_0_dataflow_b;
	reg mesh_4_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_16_io_in_control_0_shift_b;
	reg mesh_5_16_io_in_control_0_dataflow_b;
	reg mesh_5_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_16_io_in_control_0_shift_b;
	reg mesh_6_16_io_in_control_0_dataflow_b;
	reg mesh_6_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_16_io_in_control_0_shift_b;
	reg mesh_7_16_io_in_control_0_dataflow_b;
	reg mesh_7_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_16_io_in_control_0_shift_b;
	reg mesh_8_16_io_in_control_0_dataflow_b;
	reg mesh_8_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_16_io_in_control_0_shift_b;
	reg mesh_9_16_io_in_control_0_dataflow_b;
	reg mesh_9_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_16_io_in_control_0_shift_b;
	reg mesh_10_16_io_in_control_0_dataflow_b;
	reg mesh_10_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_16_io_in_control_0_shift_b;
	reg mesh_11_16_io_in_control_0_dataflow_b;
	reg mesh_11_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_16_io_in_control_0_shift_b;
	reg mesh_12_16_io_in_control_0_dataflow_b;
	reg mesh_12_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_16_io_in_control_0_shift_b;
	reg mesh_13_16_io_in_control_0_dataflow_b;
	reg mesh_13_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_16_io_in_control_0_shift_b;
	reg mesh_14_16_io_in_control_0_dataflow_b;
	reg mesh_14_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_16_io_in_control_0_shift_b;
	reg mesh_15_16_io_in_control_0_dataflow_b;
	reg mesh_15_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_16_io_in_control_0_shift_b;
	reg mesh_16_16_io_in_control_0_dataflow_b;
	reg mesh_16_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_16_io_in_control_0_shift_b;
	reg mesh_17_16_io_in_control_0_dataflow_b;
	reg mesh_17_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_16_io_in_control_0_shift_b;
	reg mesh_18_16_io_in_control_0_dataflow_b;
	reg mesh_18_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_16_io_in_control_0_shift_b;
	reg mesh_19_16_io_in_control_0_dataflow_b;
	reg mesh_19_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_16_io_in_control_0_shift_b;
	reg mesh_20_16_io_in_control_0_dataflow_b;
	reg mesh_20_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_16_io_in_control_0_shift_b;
	reg mesh_21_16_io_in_control_0_dataflow_b;
	reg mesh_21_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_16_io_in_control_0_shift_b;
	reg mesh_22_16_io_in_control_0_dataflow_b;
	reg mesh_22_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_16_io_in_control_0_shift_b;
	reg mesh_23_16_io_in_control_0_dataflow_b;
	reg mesh_23_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_16_io_in_control_0_shift_b;
	reg mesh_24_16_io_in_control_0_dataflow_b;
	reg mesh_24_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_16_io_in_control_0_shift_b;
	reg mesh_25_16_io_in_control_0_dataflow_b;
	reg mesh_25_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_16_io_in_control_0_shift_b;
	reg mesh_26_16_io_in_control_0_dataflow_b;
	reg mesh_26_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_16_io_in_control_0_shift_b;
	reg mesh_27_16_io_in_control_0_dataflow_b;
	reg mesh_27_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_16_io_in_control_0_shift_b;
	reg mesh_28_16_io_in_control_0_dataflow_b;
	reg mesh_28_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_16_io_in_control_0_shift_b;
	reg mesh_29_16_io_in_control_0_dataflow_b;
	reg mesh_29_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_16_io_in_control_0_shift_b;
	reg mesh_30_16_io_in_control_0_dataflow_b;
	reg mesh_30_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_16_io_in_control_0_shift_b;
	reg mesh_31_16_io_in_control_0_dataflow_b;
	reg mesh_31_16_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_17_io_in_control_0_shift_b;
	reg mesh_0_17_io_in_control_0_dataflow_b;
	reg mesh_0_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_17_io_in_control_0_shift_b;
	reg mesh_1_17_io_in_control_0_dataflow_b;
	reg mesh_1_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_17_io_in_control_0_shift_b;
	reg mesh_2_17_io_in_control_0_dataflow_b;
	reg mesh_2_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_17_io_in_control_0_shift_b;
	reg mesh_3_17_io_in_control_0_dataflow_b;
	reg mesh_3_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_17_io_in_control_0_shift_b;
	reg mesh_4_17_io_in_control_0_dataflow_b;
	reg mesh_4_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_17_io_in_control_0_shift_b;
	reg mesh_5_17_io_in_control_0_dataflow_b;
	reg mesh_5_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_17_io_in_control_0_shift_b;
	reg mesh_6_17_io_in_control_0_dataflow_b;
	reg mesh_6_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_17_io_in_control_0_shift_b;
	reg mesh_7_17_io_in_control_0_dataflow_b;
	reg mesh_7_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_17_io_in_control_0_shift_b;
	reg mesh_8_17_io_in_control_0_dataflow_b;
	reg mesh_8_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_17_io_in_control_0_shift_b;
	reg mesh_9_17_io_in_control_0_dataflow_b;
	reg mesh_9_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_17_io_in_control_0_shift_b;
	reg mesh_10_17_io_in_control_0_dataflow_b;
	reg mesh_10_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_17_io_in_control_0_shift_b;
	reg mesh_11_17_io_in_control_0_dataflow_b;
	reg mesh_11_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_17_io_in_control_0_shift_b;
	reg mesh_12_17_io_in_control_0_dataflow_b;
	reg mesh_12_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_17_io_in_control_0_shift_b;
	reg mesh_13_17_io_in_control_0_dataflow_b;
	reg mesh_13_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_17_io_in_control_0_shift_b;
	reg mesh_14_17_io_in_control_0_dataflow_b;
	reg mesh_14_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_17_io_in_control_0_shift_b;
	reg mesh_15_17_io_in_control_0_dataflow_b;
	reg mesh_15_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_17_io_in_control_0_shift_b;
	reg mesh_16_17_io_in_control_0_dataflow_b;
	reg mesh_16_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_17_io_in_control_0_shift_b;
	reg mesh_17_17_io_in_control_0_dataflow_b;
	reg mesh_17_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_17_io_in_control_0_shift_b;
	reg mesh_18_17_io_in_control_0_dataflow_b;
	reg mesh_18_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_17_io_in_control_0_shift_b;
	reg mesh_19_17_io_in_control_0_dataflow_b;
	reg mesh_19_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_17_io_in_control_0_shift_b;
	reg mesh_20_17_io_in_control_0_dataflow_b;
	reg mesh_20_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_17_io_in_control_0_shift_b;
	reg mesh_21_17_io_in_control_0_dataflow_b;
	reg mesh_21_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_17_io_in_control_0_shift_b;
	reg mesh_22_17_io_in_control_0_dataflow_b;
	reg mesh_22_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_17_io_in_control_0_shift_b;
	reg mesh_23_17_io_in_control_0_dataflow_b;
	reg mesh_23_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_17_io_in_control_0_shift_b;
	reg mesh_24_17_io_in_control_0_dataflow_b;
	reg mesh_24_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_17_io_in_control_0_shift_b;
	reg mesh_25_17_io_in_control_0_dataflow_b;
	reg mesh_25_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_17_io_in_control_0_shift_b;
	reg mesh_26_17_io_in_control_0_dataflow_b;
	reg mesh_26_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_17_io_in_control_0_shift_b;
	reg mesh_27_17_io_in_control_0_dataflow_b;
	reg mesh_27_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_17_io_in_control_0_shift_b;
	reg mesh_28_17_io_in_control_0_dataflow_b;
	reg mesh_28_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_17_io_in_control_0_shift_b;
	reg mesh_29_17_io_in_control_0_dataflow_b;
	reg mesh_29_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_17_io_in_control_0_shift_b;
	reg mesh_30_17_io_in_control_0_dataflow_b;
	reg mesh_30_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_17_io_in_control_0_shift_b;
	reg mesh_31_17_io_in_control_0_dataflow_b;
	reg mesh_31_17_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_18_io_in_control_0_shift_b;
	reg mesh_0_18_io_in_control_0_dataflow_b;
	reg mesh_0_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_18_io_in_control_0_shift_b;
	reg mesh_1_18_io_in_control_0_dataflow_b;
	reg mesh_1_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_18_io_in_control_0_shift_b;
	reg mesh_2_18_io_in_control_0_dataflow_b;
	reg mesh_2_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_18_io_in_control_0_shift_b;
	reg mesh_3_18_io_in_control_0_dataflow_b;
	reg mesh_3_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_18_io_in_control_0_shift_b;
	reg mesh_4_18_io_in_control_0_dataflow_b;
	reg mesh_4_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_18_io_in_control_0_shift_b;
	reg mesh_5_18_io_in_control_0_dataflow_b;
	reg mesh_5_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_18_io_in_control_0_shift_b;
	reg mesh_6_18_io_in_control_0_dataflow_b;
	reg mesh_6_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_18_io_in_control_0_shift_b;
	reg mesh_7_18_io_in_control_0_dataflow_b;
	reg mesh_7_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_18_io_in_control_0_shift_b;
	reg mesh_8_18_io_in_control_0_dataflow_b;
	reg mesh_8_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_18_io_in_control_0_shift_b;
	reg mesh_9_18_io_in_control_0_dataflow_b;
	reg mesh_9_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_18_io_in_control_0_shift_b;
	reg mesh_10_18_io_in_control_0_dataflow_b;
	reg mesh_10_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_18_io_in_control_0_shift_b;
	reg mesh_11_18_io_in_control_0_dataflow_b;
	reg mesh_11_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_18_io_in_control_0_shift_b;
	reg mesh_12_18_io_in_control_0_dataflow_b;
	reg mesh_12_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_18_io_in_control_0_shift_b;
	reg mesh_13_18_io_in_control_0_dataflow_b;
	reg mesh_13_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_18_io_in_control_0_shift_b;
	reg mesh_14_18_io_in_control_0_dataflow_b;
	reg mesh_14_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_18_io_in_control_0_shift_b;
	reg mesh_15_18_io_in_control_0_dataflow_b;
	reg mesh_15_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_18_io_in_control_0_shift_b;
	reg mesh_16_18_io_in_control_0_dataflow_b;
	reg mesh_16_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_18_io_in_control_0_shift_b;
	reg mesh_17_18_io_in_control_0_dataflow_b;
	reg mesh_17_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_18_io_in_control_0_shift_b;
	reg mesh_18_18_io_in_control_0_dataflow_b;
	reg mesh_18_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_18_io_in_control_0_shift_b;
	reg mesh_19_18_io_in_control_0_dataflow_b;
	reg mesh_19_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_18_io_in_control_0_shift_b;
	reg mesh_20_18_io_in_control_0_dataflow_b;
	reg mesh_20_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_18_io_in_control_0_shift_b;
	reg mesh_21_18_io_in_control_0_dataflow_b;
	reg mesh_21_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_18_io_in_control_0_shift_b;
	reg mesh_22_18_io_in_control_0_dataflow_b;
	reg mesh_22_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_18_io_in_control_0_shift_b;
	reg mesh_23_18_io_in_control_0_dataflow_b;
	reg mesh_23_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_18_io_in_control_0_shift_b;
	reg mesh_24_18_io_in_control_0_dataflow_b;
	reg mesh_24_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_18_io_in_control_0_shift_b;
	reg mesh_25_18_io_in_control_0_dataflow_b;
	reg mesh_25_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_18_io_in_control_0_shift_b;
	reg mesh_26_18_io_in_control_0_dataflow_b;
	reg mesh_26_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_18_io_in_control_0_shift_b;
	reg mesh_27_18_io_in_control_0_dataflow_b;
	reg mesh_27_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_18_io_in_control_0_shift_b;
	reg mesh_28_18_io_in_control_0_dataflow_b;
	reg mesh_28_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_18_io_in_control_0_shift_b;
	reg mesh_29_18_io_in_control_0_dataflow_b;
	reg mesh_29_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_18_io_in_control_0_shift_b;
	reg mesh_30_18_io_in_control_0_dataflow_b;
	reg mesh_30_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_18_io_in_control_0_shift_b;
	reg mesh_31_18_io_in_control_0_dataflow_b;
	reg mesh_31_18_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_19_io_in_control_0_shift_b;
	reg mesh_0_19_io_in_control_0_dataflow_b;
	reg mesh_0_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_19_io_in_control_0_shift_b;
	reg mesh_1_19_io_in_control_0_dataflow_b;
	reg mesh_1_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_19_io_in_control_0_shift_b;
	reg mesh_2_19_io_in_control_0_dataflow_b;
	reg mesh_2_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_19_io_in_control_0_shift_b;
	reg mesh_3_19_io_in_control_0_dataflow_b;
	reg mesh_3_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_19_io_in_control_0_shift_b;
	reg mesh_4_19_io_in_control_0_dataflow_b;
	reg mesh_4_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_19_io_in_control_0_shift_b;
	reg mesh_5_19_io_in_control_0_dataflow_b;
	reg mesh_5_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_19_io_in_control_0_shift_b;
	reg mesh_6_19_io_in_control_0_dataflow_b;
	reg mesh_6_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_19_io_in_control_0_shift_b;
	reg mesh_7_19_io_in_control_0_dataflow_b;
	reg mesh_7_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_19_io_in_control_0_shift_b;
	reg mesh_8_19_io_in_control_0_dataflow_b;
	reg mesh_8_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_19_io_in_control_0_shift_b;
	reg mesh_9_19_io_in_control_0_dataflow_b;
	reg mesh_9_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_19_io_in_control_0_shift_b;
	reg mesh_10_19_io_in_control_0_dataflow_b;
	reg mesh_10_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_19_io_in_control_0_shift_b;
	reg mesh_11_19_io_in_control_0_dataflow_b;
	reg mesh_11_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_19_io_in_control_0_shift_b;
	reg mesh_12_19_io_in_control_0_dataflow_b;
	reg mesh_12_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_19_io_in_control_0_shift_b;
	reg mesh_13_19_io_in_control_0_dataflow_b;
	reg mesh_13_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_19_io_in_control_0_shift_b;
	reg mesh_14_19_io_in_control_0_dataflow_b;
	reg mesh_14_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_19_io_in_control_0_shift_b;
	reg mesh_15_19_io_in_control_0_dataflow_b;
	reg mesh_15_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_19_io_in_control_0_shift_b;
	reg mesh_16_19_io_in_control_0_dataflow_b;
	reg mesh_16_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_19_io_in_control_0_shift_b;
	reg mesh_17_19_io_in_control_0_dataflow_b;
	reg mesh_17_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_19_io_in_control_0_shift_b;
	reg mesh_18_19_io_in_control_0_dataflow_b;
	reg mesh_18_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_19_io_in_control_0_shift_b;
	reg mesh_19_19_io_in_control_0_dataflow_b;
	reg mesh_19_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_19_io_in_control_0_shift_b;
	reg mesh_20_19_io_in_control_0_dataflow_b;
	reg mesh_20_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_19_io_in_control_0_shift_b;
	reg mesh_21_19_io_in_control_0_dataflow_b;
	reg mesh_21_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_19_io_in_control_0_shift_b;
	reg mesh_22_19_io_in_control_0_dataflow_b;
	reg mesh_22_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_19_io_in_control_0_shift_b;
	reg mesh_23_19_io_in_control_0_dataflow_b;
	reg mesh_23_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_19_io_in_control_0_shift_b;
	reg mesh_24_19_io_in_control_0_dataflow_b;
	reg mesh_24_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_19_io_in_control_0_shift_b;
	reg mesh_25_19_io_in_control_0_dataflow_b;
	reg mesh_25_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_19_io_in_control_0_shift_b;
	reg mesh_26_19_io_in_control_0_dataflow_b;
	reg mesh_26_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_19_io_in_control_0_shift_b;
	reg mesh_27_19_io_in_control_0_dataflow_b;
	reg mesh_27_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_19_io_in_control_0_shift_b;
	reg mesh_28_19_io_in_control_0_dataflow_b;
	reg mesh_28_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_19_io_in_control_0_shift_b;
	reg mesh_29_19_io_in_control_0_dataflow_b;
	reg mesh_29_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_19_io_in_control_0_shift_b;
	reg mesh_30_19_io_in_control_0_dataflow_b;
	reg mesh_30_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_19_io_in_control_0_shift_b;
	reg mesh_31_19_io_in_control_0_dataflow_b;
	reg mesh_31_19_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_20_io_in_control_0_shift_b;
	reg mesh_0_20_io_in_control_0_dataflow_b;
	reg mesh_0_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_20_io_in_control_0_shift_b;
	reg mesh_1_20_io_in_control_0_dataflow_b;
	reg mesh_1_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_20_io_in_control_0_shift_b;
	reg mesh_2_20_io_in_control_0_dataflow_b;
	reg mesh_2_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_20_io_in_control_0_shift_b;
	reg mesh_3_20_io_in_control_0_dataflow_b;
	reg mesh_3_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_20_io_in_control_0_shift_b;
	reg mesh_4_20_io_in_control_0_dataflow_b;
	reg mesh_4_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_20_io_in_control_0_shift_b;
	reg mesh_5_20_io_in_control_0_dataflow_b;
	reg mesh_5_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_20_io_in_control_0_shift_b;
	reg mesh_6_20_io_in_control_0_dataflow_b;
	reg mesh_6_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_20_io_in_control_0_shift_b;
	reg mesh_7_20_io_in_control_0_dataflow_b;
	reg mesh_7_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_20_io_in_control_0_shift_b;
	reg mesh_8_20_io_in_control_0_dataflow_b;
	reg mesh_8_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_20_io_in_control_0_shift_b;
	reg mesh_9_20_io_in_control_0_dataflow_b;
	reg mesh_9_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_20_io_in_control_0_shift_b;
	reg mesh_10_20_io_in_control_0_dataflow_b;
	reg mesh_10_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_20_io_in_control_0_shift_b;
	reg mesh_11_20_io_in_control_0_dataflow_b;
	reg mesh_11_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_20_io_in_control_0_shift_b;
	reg mesh_12_20_io_in_control_0_dataflow_b;
	reg mesh_12_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_20_io_in_control_0_shift_b;
	reg mesh_13_20_io_in_control_0_dataflow_b;
	reg mesh_13_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_20_io_in_control_0_shift_b;
	reg mesh_14_20_io_in_control_0_dataflow_b;
	reg mesh_14_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_20_io_in_control_0_shift_b;
	reg mesh_15_20_io_in_control_0_dataflow_b;
	reg mesh_15_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_20_io_in_control_0_shift_b;
	reg mesh_16_20_io_in_control_0_dataflow_b;
	reg mesh_16_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_20_io_in_control_0_shift_b;
	reg mesh_17_20_io_in_control_0_dataflow_b;
	reg mesh_17_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_20_io_in_control_0_shift_b;
	reg mesh_18_20_io_in_control_0_dataflow_b;
	reg mesh_18_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_20_io_in_control_0_shift_b;
	reg mesh_19_20_io_in_control_0_dataflow_b;
	reg mesh_19_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_20_io_in_control_0_shift_b;
	reg mesh_20_20_io_in_control_0_dataflow_b;
	reg mesh_20_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_20_io_in_control_0_shift_b;
	reg mesh_21_20_io_in_control_0_dataflow_b;
	reg mesh_21_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_20_io_in_control_0_shift_b;
	reg mesh_22_20_io_in_control_0_dataflow_b;
	reg mesh_22_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_20_io_in_control_0_shift_b;
	reg mesh_23_20_io_in_control_0_dataflow_b;
	reg mesh_23_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_20_io_in_control_0_shift_b;
	reg mesh_24_20_io_in_control_0_dataflow_b;
	reg mesh_24_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_20_io_in_control_0_shift_b;
	reg mesh_25_20_io_in_control_0_dataflow_b;
	reg mesh_25_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_20_io_in_control_0_shift_b;
	reg mesh_26_20_io_in_control_0_dataflow_b;
	reg mesh_26_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_20_io_in_control_0_shift_b;
	reg mesh_27_20_io_in_control_0_dataflow_b;
	reg mesh_27_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_20_io_in_control_0_shift_b;
	reg mesh_28_20_io_in_control_0_dataflow_b;
	reg mesh_28_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_20_io_in_control_0_shift_b;
	reg mesh_29_20_io_in_control_0_dataflow_b;
	reg mesh_29_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_20_io_in_control_0_shift_b;
	reg mesh_30_20_io_in_control_0_dataflow_b;
	reg mesh_30_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_20_io_in_control_0_shift_b;
	reg mesh_31_20_io_in_control_0_dataflow_b;
	reg mesh_31_20_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_21_io_in_control_0_shift_b;
	reg mesh_0_21_io_in_control_0_dataflow_b;
	reg mesh_0_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_21_io_in_control_0_shift_b;
	reg mesh_1_21_io_in_control_0_dataflow_b;
	reg mesh_1_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_21_io_in_control_0_shift_b;
	reg mesh_2_21_io_in_control_0_dataflow_b;
	reg mesh_2_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_21_io_in_control_0_shift_b;
	reg mesh_3_21_io_in_control_0_dataflow_b;
	reg mesh_3_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_21_io_in_control_0_shift_b;
	reg mesh_4_21_io_in_control_0_dataflow_b;
	reg mesh_4_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_21_io_in_control_0_shift_b;
	reg mesh_5_21_io_in_control_0_dataflow_b;
	reg mesh_5_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_21_io_in_control_0_shift_b;
	reg mesh_6_21_io_in_control_0_dataflow_b;
	reg mesh_6_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_21_io_in_control_0_shift_b;
	reg mesh_7_21_io_in_control_0_dataflow_b;
	reg mesh_7_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_21_io_in_control_0_shift_b;
	reg mesh_8_21_io_in_control_0_dataflow_b;
	reg mesh_8_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_21_io_in_control_0_shift_b;
	reg mesh_9_21_io_in_control_0_dataflow_b;
	reg mesh_9_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_21_io_in_control_0_shift_b;
	reg mesh_10_21_io_in_control_0_dataflow_b;
	reg mesh_10_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_21_io_in_control_0_shift_b;
	reg mesh_11_21_io_in_control_0_dataflow_b;
	reg mesh_11_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_21_io_in_control_0_shift_b;
	reg mesh_12_21_io_in_control_0_dataflow_b;
	reg mesh_12_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_21_io_in_control_0_shift_b;
	reg mesh_13_21_io_in_control_0_dataflow_b;
	reg mesh_13_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_21_io_in_control_0_shift_b;
	reg mesh_14_21_io_in_control_0_dataflow_b;
	reg mesh_14_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_21_io_in_control_0_shift_b;
	reg mesh_15_21_io_in_control_0_dataflow_b;
	reg mesh_15_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_21_io_in_control_0_shift_b;
	reg mesh_16_21_io_in_control_0_dataflow_b;
	reg mesh_16_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_21_io_in_control_0_shift_b;
	reg mesh_17_21_io_in_control_0_dataflow_b;
	reg mesh_17_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_21_io_in_control_0_shift_b;
	reg mesh_18_21_io_in_control_0_dataflow_b;
	reg mesh_18_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_21_io_in_control_0_shift_b;
	reg mesh_19_21_io_in_control_0_dataflow_b;
	reg mesh_19_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_21_io_in_control_0_shift_b;
	reg mesh_20_21_io_in_control_0_dataflow_b;
	reg mesh_20_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_21_io_in_control_0_shift_b;
	reg mesh_21_21_io_in_control_0_dataflow_b;
	reg mesh_21_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_21_io_in_control_0_shift_b;
	reg mesh_22_21_io_in_control_0_dataflow_b;
	reg mesh_22_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_21_io_in_control_0_shift_b;
	reg mesh_23_21_io_in_control_0_dataflow_b;
	reg mesh_23_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_21_io_in_control_0_shift_b;
	reg mesh_24_21_io_in_control_0_dataflow_b;
	reg mesh_24_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_21_io_in_control_0_shift_b;
	reg mesh_25_21_io_in_control_0_dataflow_b;
	reg mesh_25_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_21_io_in_control_0_shift_b;
	reg mesh_26_21_io_in_control_0_dataflow_b;
	reg mesh_26_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_21_io_in_control_0_shift_b;
	reg mesh_27_21_io_in_control_0_dataflow_b;
	reg mesh_27_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_21_io_in_control_0_shift_b;
	reg mesh_28_21_io_in_control_0_dataflow_b;
	reg mesh_28_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_21_io_in_control_0_shift_b;
	reg mesh_29_21_io_in_control_0_dataflow_b;
	reg mesh_29_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_21_io_in_control_0_shift_b;
	reg mesh_30_21_io_in_control_0_dataflow_b;
	reg mesh_30_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_21_io_in_control_0_shift_b;
	reg mesh_31_21_io_in_control_0_dataflow_b;
	reg mesh_31_21_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_22_io_in_control_0_shift_b;
	reg mesh_0_22_io_in_control_0_dataflow_b;
	reg mesh_0_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_22_io_in_control_0_shift_b;
	reg mesh_1_22_io_in_control_0_dataflow_b;
	reg mesh_1_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_22_io_in_control_0_shift_b;
	reg mesh_2_22_io_in_control_0_dataflow_b;
	reg mesh_2_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_22_io_in_control_0_shift_b;
	reg mesh_3_22_io_in_control_0_dataflow_b;
	reg mesh_3_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_22_io_in_control_0_shift_b;
	reg mesh_4_22_io_in_control_0_dataflow_b;
	reg mesh_4_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_22_io_in_control_0_shift_b;
	reg mesh_5_22_io_in_control_0_dataflow_b;
	reg mesh_5_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_22_io_in_control_0_shift_b;
	reg mesh_6_22_io_in_control_0_dataflow_b;
	reg mesh_6_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_22_io_in_control_0_shift_b;
	reg mesh_7_22_io_in_control_0_dataflow_b;
	reg mesh_7_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_22_io_in_control_0_shift_b;
	reg mesh_8_22_io_in_control_0_dataflow_b;
	reg mesh_8_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_22_io_in_control_0_shift_b;
	reg mesh_9_22_io_in_control_0_dataflow_b;
	reg mesh_9_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_22_io_in_control_0_shift_b;
	reg mesh_10_22_io_in_control_0_dataflow_b;
	reg mesh_10_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_22_io_in_control_0_shift_b;
	reg mesh_11_22_io_in_control_0_dataflow_b;
	reg mesh_11_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_22_io_in_control_0_shift_b;
	reg mesh_12_22_io_in_control_0_dataflow_b;
	reg mesh_12_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_22_io_in_control_0_shift_b;
	reg mesh_13_22_io_in_control_0_dataflow_b;
	reg mesh_13_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_22_io_in_control_0_shift_b;
	reg mesh_14_22_io_in_control_0_dataflow_b;
	reg mesh_14_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_22_io_in_control_0_shift_b;
	reg mesh_15_22_io_in_control_0_dataflow_b;
	reg mesh_15_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_22_io_in_control_0_shift_b;
	reg mesh_16_22_io_in_control_0_dataflow_b;
	reg mesh_16_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_22_io_in_control_0_shift_b;
	reg mesh_17_22_io_in_control_0_dataflow_b;
	reg mesh_17_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_22_io_in_control_0_shift_b;
	reg mesh_18_22_io_in_control_0_dataflow_b;
	reg mesh_18_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_22_io_in_control_0_shift_b;
	reg mesh_19_22_io_in_control_0_dataflow_b;
	reg mesh_19_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_22_io_in_control_0_shift_b;
	reg mesh_20_22_io_in_control_0_dataflow_b;
	reg mesh_20_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_22_io_in_control_0_shift_b;
	reg mesh_21_22_io_in_control_0_dataflow_b;
	reg mesh_21_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_22_io_in_control_0_shift_b;
	reg mesh_22_22_io_in_control_0_dataflow_b;
	reg mesh_22_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_22_io_in_control_0_shift_b;
	reg mesh_23_22_io_in_control_0_dataflow_b;
	reg mesh_23_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_22_io_in_control_0_shift_b;
	reg mesh_24_22_io_in_control_0_dataflow_b;
	reg mesh_24_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_22_io_in_control_0_shift_b;
	reg mesh_25_22_io_in_control_0_dataflow_b;
	reg mesh_25_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_22_io_in_control_0_shift_b;
	reg mesh_26_22_io_in_control_0_dataflow_b;
	reg mesh_26_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_22_io_in_control_0_shift_b;
	reg mesh_27_22_io_in_control_0_dataflow_b;
	reg mesh_27_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_22_io_in_control_0_shift_b;
	reg mesh_28_22_io_in_control_0_dataflow_b;
	reg mesh_28_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_22_io_in_control_0_shift_b;
	reg mesh_29_22_io_in_control_0_dataflow_b;
	reg mesh_29_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_22_io_in_control_0_shift_b;
	reg mesh_30_22_io_in_control_0_dataflow_b;
	reg mesh_30_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_22_io_in_control_0_shift_b;
	reg mesh_31_22_io_in_control_0_dataflow_b;
	reg mesh_31_22_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_23_io_in_control_0_shift_b;
	reg mesh_0_23_io_in_control_0_dataflow_b;
	reg mesh_0_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_23_io_in_control_0_shift_b;
	reg mesh_1_23_io_in_control_0_dataflow_b;
	reg mesh_1_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_23_io_in_control_0_shift_b;
	reg mesh_2_23_io_in_control_0_dataflow_b;
	reg mesh_2_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_23_io_in_control_0_shift_b;
	reg mesh_3_23_io_in_control_0_dataflow_b;
	reg mesh_3_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_23_io_in_control_0_shift_b;
	reg mesh_4_23_io_in_control_0_dataflow_b;
	reg mesh_4_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_23_io_in_control_0_shift_b;
	reg mesh_5_23_io_in_control_0_dataflow_b;
	reg mesh_5_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_23_io_in_control_0_shift_b;
	reg mesh_6_23_io_in_control_0_dataflow_b;
	reg mesh_6_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_23_io_in_control_0_shift_b;
	reg mesh_7_23_io_in_control_0_dataflow_b;
	reg mesh_7_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_23_io_in_control_0_shift_b;
	reg mesh_8_23_io_in_control_0_dataflow_b;
	reg mesh_8_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_23_io_in_control_0_shift_b;
	reg mesh_9_23_io_in_control_0_dataflow_b;
	reg mesh_9_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_23_io_in_control_0_shift_b;
	reg mesh_10_23_io_in_control_0_dataflow_b;
	reg mesh_10_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_23_io_in_control_0_shift_b;
	reg mesh_11_23_io_in_control_0_dataflow_b;
	reg mesh_11_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_23_io_in_control_0_shift_b;
	reg mesh_12_23_io_in_control_0_dataflow_b;
	reg mesh_12_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_23_io_in_control_0_shift_b;
	reg mesh_13_23_io_in_control_0_dataflow_b;
	reg mesh_13_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_23_io_in_control_0_shift_b;
	reg mesh_14_23_io_in_control_0_dataflow_b;
	reg mesh_14_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_23_io_in_control_0_shift_b;
	reg mesh_15_23_io_in_control_0_dataflow_b;
	reg mesh_15_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_23_io_in_control_0_shift_b;
	reg mesh_16_23_io_in_control_0_dataflow_b;
	reg mesh_16_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_23_io_in_control_0_shift_b;
	reg mesh_17_23_io_in_control_0_dataflow_b;
	reg mesh_17_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_23_io_in_control_0_shift_b;
	reg mesh_18_23_io_in_control_0_dataflow_b;
	reg mesh_18_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_23_io_in_control_0_shift_b;
	reg mesh_19_23_io_in_control_0_dataflow_b;
	reg mesh_19_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_23_io_in_control_0_shift_b;
	reg mesh_20_23_io_in_control_0_dataflow_b;
	reg mesh_20_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_23_io_in_control_0_shift_b;
	reg mesh_21_23_io_in_control_0_dataflow_b;
	reg mesh_21_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_23_io_in_control_0_shift_b;
	reg mesh_22_23_io_in_control_0_dataflow_b;
	reg mesh_22_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_23_io_in_control_0_shift_b;
	reg mesh_23_23_io_in_control_0_dataflow_b;
	reg mesh_23_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_23_io_in_control_0_shift_b;
	reg mesh_24_23_io_in_control_0_dataflow_b;
	reg mesh_24_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_23_io_in_control_0_shift_b;
	reg mesh_25_23_io_in_control_0_dataflow_b;
	reg mesh_25_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_23_io_in_control_0_shift_b;
	reg mesh_26_23_io_in_control_0_dataflow_b;
	reg mesh_26_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_23_io_in_control_0_shift_b;
	reg mesh_27_23_io_in_control_0_dataflow_b;
	reg mesh_27_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_23_io_in_control_0_shift_b;
	reg mesh_28_23_io_in_control_0_dataflow_b;
	reg mesh_28_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_23_io_in_control_0_shift_b;
	reg mesh_29_23_io_in_control_0_dataflow_b;
	reg mesh_29_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_23_io_in_control_0_shift_b;
	reg mesh_30_23_io_in_control_0_dataflow_b;
	reg mesh_30_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_23_io_in_control_0_shift_b;
	reg mesh_31_23_io_in_control_0_dataflow_b;
	reg mesh_31_23_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_24_io_in_control_0_shift_b;
	reg mesh_0_24_io_in_control_0_dataflow_b;
	reg mesh_0_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_24_io_in_control_0_shift_b;
	reg mesh_1_24_io_in_control_0_dataflow_b;
	reg mesh_1_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_24_io_in_control_0_shift_b;
	reg mesh_2_24_io_in_control_0_dataflow_b;
	reg mesh_2_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_24_io_in_control_0_shift_b;
	reg mesh_3_24_io_in_control_0_dataflow_b;
	reg mesh_3_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_24_io_in_control_0_shift_b;
	reg mesh_4_24_io_in_control_0_dataflow_b;
	reg mesh_4_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_24_io_in_control_0_shift_b;
	reg mesh_5_24_io_in_control_0_dataflow_b;
	reg mesh_5_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_24_io_in_control_0_shift_b;
	reg mesh_6_24_io_in_control_0_dataflow_b;
	reg mesh_6_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_24_io_in_control_0_shift_b;
	reg mesh_7_24_io_in_control_0_dataflow_b;
	reg mesh_7_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_24_io_in_control_0_shift_b;
	reg mesh_8_24_io_in_control_0_dataflow_b;
	reg mesh_8_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_24_io_in_control_0_shift_b;
	reg mesh_9_24_io_in_control_0_dataflow_b;
	reg mesh_9_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_24_io_in_control_0_shift_b;
	reg mesh_10_24_io_in_control_0_dataflow_b;
	reg mesh_10_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_24_io_in_control_0_shift_b;
	reg mesh_11_24_io_in_control_0_dataflow_b;
	reg mesh_11_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_24_io_in_control_0_shift_b;
	reg mesh_12_24_io_in_control_0_dataflow_b;
	reg mesh_12_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_24_io_in_control_0_shift_b;
	reg mesh_13_24_io_in_control_0_dataflow_b;
	reg mesh_13_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_24_io_in_control_0_shift_b;
	reg mesh_14_24_io_in_control_0_dataflow_b;
	reg mesh_14_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_24_io_in_control_0_shift_b;
	reg mesh_15_24_io_in_control_0_dataflow_b;
	reg mesh_15_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_24_io_in_control_0_shift_b;
	reg mesh_16_24_io_in_control_0_dataflow_b;
	reg mesh_16_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_24_io_in_control_0_shift_b;
	reg mesh_17_24_io_in_control_0_dataflow_b;
	reg mesh_17_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_24_io_in_control_0_shift_b;
	reg mesh_18_24_io_in_control_0_dataflow_b;
	reg mesh_18_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_24_io_in_control_0_shift_b;
	reg mesh_19_24_io_in_control_0_dataflow_b;
	reg mesh_19_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_24_io_in_control_0_shift_b;
	reg mesh_20_24_io_in_control_0_dataflow_b;
	reg mesh_20_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_24_io_in_control_0_shift_b;
	reg mesh_21_24_io_in_control_0_dataflow_b;
	reg mesh_21_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_24_io_in_control_0_shift_b;
	reg mesh_22_24_io_in_control_0_dataflow_b;
	reg mesh_22_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_24_io_in_control_0_shift_b;
	reg mesh_23_24_io_in_control_0_dataflow_b;
	reg mesh_23_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_24_io_in_control_0_shift_b;
	reg mesh_24_24_io_in_control_0_dataflow_b;
	reg mesh_24_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_24_io_in_control_0_shift_b;
	reg mesh_25_24_io_in_control_0_dataflow_b;
	reg mesh_25_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_24_io_in_control_0_shift_b;
	reg mesh_26_24_io_in_control_0_dataflow_b;
	reg mesh_26_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_24_io_in_control_0_shift_b;
	reg mesh_27_24_io_in_control_0_dataflow_b;
	reg mesh_27_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_24_io_in_control_0_shift_b;
	reg mesh_28_24_io_in_control_0_dataflow_b;
	reg mesh_28_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_24_io_in_control_0_shift_b;
	reg mesh_29_24_io_in_control_0_dataflow_b;
	reg mesh_29_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_24_io_in_control_0_shift_b;
	reg mesh_30_24_io_in_control_0_dataflow_b;
	reg mesh_30_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_24_io_in_control_0_shift_b;
	reg mesh_31_24_io_in_control_0_dataflow_b;
	reg mesh_31_24_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_25_io_in_control_0_shift_b;
	reg mesh_0_25_io_in_control_0_dataflow_b;
	reg mesh_0_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_25_io_in_control_0_shift_b;
	reg mesh_1_25_io_in_control_0_dataflow_b;
	reg mesh_1_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_25_io_in_control_0_shift_b;
	reg mesh_2_25_io_in_control_0_dataflow_b;
	reg mesh_2_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_25_io_in_control_0_shift_b;
	reg mesh_3_25_io_in_control_0_dataflow_b;
	reg mesh_3_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_25_io_in_control_0_shift_b;
	reg mesh_4_25_io_in_control_0_dataflow_b;
	reg mesh_4_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_25_io_in_control_0_shift_b;
	reg mesh_5_25_io_in_control_0_dataflow_b;
	reg mesh_5_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_25_io_in_control_0_shift_b;
	reg mesh_6_25_io_in_control_0_dataflow_b;
	reg mesh_6_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_25_io_in_control_0_shift_b;
	reg mesh_7_25_io_in_control_0_dataflow_b;
	reg mesh_7_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_25_io_in_control_0_shift_b;
	reg mesh_8_25_io_in_control_0_dataflow_b;
	reg mesh_8_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_25_io_in_control_0_shift_b;
	reg mesh_9_25_io_in_control_0_dataflow_b;
	reg mesh_9_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_25_io_in_control_0_shift_b;
	reg mesh_10_25_io_in_control_0_dataflow_b;
	reg mesh_10_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_25_io_in_control_0_shift_b;
	reg mesh_11_25_io_in_control_0_dataflow_b;
	reg mesh_11_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_25_io_in_control_0_shift_b;
	reg mesh_12_25_io_in_control_0_dataflow_b;
	reg mesh_12_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_25_io_in_control_0_shift_b;
	reg mesh_13_25_io_in_control_0_dataflow_b;
	reg mesh_13_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_25_io_in_control_0_shift_b;
	reg mesh_14_25_io_in_control_0_dataflow_b;
	reg mesh_14_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_25_io_in_control_0_shift_b;
	reg mesh_15_25_io_in_control_0_dataflow_b;
	reg mesh_15_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_25_io_in_control_0_shift_b;
	reg mesh_16_25_io_in_control_0_dataflow_b;
	reg mesh_16_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_25_io_in_control_0_shift_b;
	reg mesh_17_25_io_in_control_0_dataflow_b;
	reg mesh_17_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_25_io_in_control_0_shift_b;
	reg mesh_18_25_io_in_control_0_dataflow_b;
	reg mesh_18_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_25_io_in_control_0_shift_b;
	reg mesh_19_25_io_in_control_0_dataflow_b;
	reg mesh_19_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_25_io_in_control_0_shift_b;
	reg mesh_20_25_io_in_control_0_dataflow_b;
	reg mesh_20_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_25_io_in_control_0_shift_b;
	reg mesh_21_25_io_in_control_0_dataflow_b;
	reg mesh_21_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_25_io_in_control_0_shift_b;
	reg mesh_22_25_io_in_control_0_dataflow_b;
	reg mesh_22_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_25_io_in_control_0_shift_b;
	reg mesh_23_25_io_in_control_0_dataflow_b;
	reg mesh_23_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_25_io_in_control_0_shift_b;
	reg mesh_24_25_io_in_control_0_dataflow_b;
	reg mesh_24_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_25_io_in_control_0_shift_b;
	reg mesh_25_25_io_in_control_0_dataflow_b;
	reg mesh_25_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_25_io_in_control_0_shift_b;
	reg mesh_26_25_io_in_control_0_dataflow_b;
	reg mesh_26_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_25_io_in_control_0_shift_b;
	reg mesh_27_25_io_in_control_0_dataflow_b;
	reg mesh_27_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_25_io_in_control_0_shift_b;
	reg mesh_28_25_io_in_control_0_dataflow_b;
	reg mesh_28_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_25_io_in_control_0_shift_b;
	reg mesh_29_25_io_in_control_0_dataflow_b;
	reg mesh_29_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_25_io_in_control_0_shift_b;
	reg mesh_30_25_io_in_control_0_dataflow_b;
	reg mesh_30_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_25_io_in_control_0_shift_b;
	reg mesh_31_25_io_in_control_0_dataflow_b;
	reg mesh_31_25_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_26_io_in_control_0_shift_b;
	reg mesh_0_26_io_in_control_0_dataflow_b;
	reg mesh_0_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_26_io_in_control_0_shift_b;
	reg mesh_1_26_io_in_control_0_dataflow_b;
	reg mesh_1_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_26_io_in_control_0_shift_b;
	reg mesh_2_26_io_in_control_0_dataflow_b;
	reg mesh_2_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_26_io_in_control_0_shift_b;
	reg mesh_3_26_io_in_control_0_dataflow_b;
	reg mesh_3_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_26_io_in_control_0_shift_b;
	reg mesh_4_26_io_in_control_0_dataflow_b;
	reg mesh_4_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_26_io_in_control_0_shift_b;
	reg mesh_5_26_io_in_control_0_dataflow_b;
	reg mesh_5_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_26_io_in_control_0_shift_b;
	reg mesh_6_26_io_in_control_0_dataflow_b;
	reg mesh_6_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_26_io_in_control_0_shift_b;
	reg mesh_7_26_io_in_control_0_dataflow_b;
	reg mesh_7_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_26_io_in_control_0_shift_b;
	reg mesh_8_26_io_in_control_0_dataflow_b;
	reg mesh_8_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_26_io_in_control_0_shift_b;
	reg mesh_9_26_io_in_control_0_dataflow_b;
	reg mesh_9_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_26_io_in_control_0_shift_b;
	reg mesh_10_26_io_in_control_0_dataflow_b;
	reg mesh_10_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_26_io_in_control_0_shift_b;
	reg mesh_11_26_io_in_control_0_dataflow_b;
	reg mesh_11_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_26_io_in_control_0_shift_b;
	reg mesh_12_26_io_in_control_0_dataflow_b;
	reg mesh_12_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_26_io_in_control_0_shift_b;
	reg mesh_13_26_io_in_control_0_dataflow_b;
	reg mesh_13_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_26_io_in_control_0_shift_b;
	reg mesh_14_26_io_in_control_0_dataflow_b;
	reg mesh_14_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_26_io_in_control_0_shift_b;
	reg mesh_15_26_io_in_control_0_dataflow_b;
	reg mesh_15_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_26_io_in_control_0_shift_b;
	reg mesh_16_26_io_in_control_0_dataflow_b;
	reg mesh_16_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_26_io_in_control_0_shift_b;
	reg mesh_17_26_io_in_control_0_dataflow_b;
	reg mesh_17_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_26_io_in_control_0_shift_b;
	reg mesh_18_26_io_in_control_0_dataflow_b;
	reg mesh_18_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_26_io_in_control_0_shift_b;
	reg mesh_19_26_io_in_control_0_dataflow_b;
	reg mesh_19_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_26_io_in_control_0_shift_b;
	reg mesh_20_26_io_in_control_0_dataflow_b;
	reg mesh_20_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_26_io_in_control_0_shift_b;
	reg mesh_21_26_io_in_control_0_dataflow_b;
	reg mesh_21_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_26_io_in_control_0_shift_b;
	reg mesh_22_26_io_in_control_0_dataflow_b;
	reg mesh_22_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_26_io_in_control_0_shift_b;
	reg mesh_23_26_io_in_control_0_dataflow_b;
	reg mesh_23_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_26_io_in_control_0_shift_b;
	reg mesh_24_26_io_in_control_0_dataflow_b;
	reg mesh_24_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_26_io_in_control_0_shift_b;
	reg mesh_25_26_io_in_control_0_dataflow_b;
	reg mesh_25_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_26_io_in_control_0_shift_b;
	reg mesh_26_26_io_in_control_0_dataflow_b;
	reg mesh_26_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_26_io_in_control_0_shift_b;
	reg mesh_27_26_io_in_control_0_dataflow_b;
	reg mesh_27_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_26_io_in_control_0_shift_b;
	reg mesh_28_26_io_in_control_0_dataflow_b;
	reg mesh_28_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_26_io_in_control_0_shift_b;
	reg mesh_29_26_io_in_control_0_dataflow_b;
	reg mesh_29_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_26_io_in_control_0_shift_b;
	reg mesh_30_26_io_in_control_0_dataflow_b;
	reg mesh_30_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_26_io_in_control_0_shift_b;
	reg mesh_31_26_io_in_control_0_dataflow_b;
	reg mesh_31_26_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_27_io_in_control_0_shift_b;
	reg mesh_0_27_io_in_control_0_dataflow_b;
	reg mesh_0_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_27_io_in_control_0_shift_b;
	reg mesh_1_27_io_in_control_0_dataflow_b;
	reg mesh_1_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_27_io_in_control_0_shift_b;
	reg mesh_2_27_io_in_control_0_dataflow_b;
	reg mesh_2_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_27_io_in_control_0_shift_b;
	reg mesh_3_27_io_in_control_0_dataflow_b;
	reg mesh_3_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_27_io_in_control_0_shift_b;
	reg mesh_4_27_io_in_control_0_dataflow_b;
	reg mesh_4_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_27_io_in_control_0_shift_b;
	reg mesh_5_27_io_in_control_0_dataflow_b;
	reg mesh_5_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_27_io_in_control_0_shift_b;
	reg mesh_6_27_io_in_control_0_dataflow_b;
	reg mesh_6_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_27_io_in_control_0_shift_b;
	reg mesh_7_27_io_in_control_0_dataflow_b;
	reg mesh_7_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_27_io_in_control_0_shift_b;
	reg mesh_8_27_io_in_control_0_dataflow_b;
	reg mesh_8_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_27_io_in_control_0_shift_b;
	reg mesh_9_27_io_in_control_0_dataflow_b;
	reg mesh_9_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_27_io_in_control_0_shift_b;
	reg mesh_10_27_io_in_control_0_dataflow_b;
	reg mesh_10_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_27_io_in_control_0_shift_b;
	reg mesh_11_27_io_in_control_0_dataflow_b;
	reg mesh_11_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_27_io_in_control_0_shift_b;
	reg mesh_12_27_io_in_control_0_dataflow_b;
	reg mesh_12_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_27_io_in_control_0_shift_b;
	reg mesh_13_27_io_in_control_0_dataflow_b;
	reg mesh_13_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_27_io_in_control_0_shift_b;
	reg mesh_14_27_io_in_control_0_dataflow_b;
	reg mesh_14_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_27_io_in_control_0_shift_b;
	reg mesh_15_27_io_in_control_0_dataflow_b;
	reg mesh_15_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_27_io_in_control_0_shift_b;
	reg mesh_16_27_io_in_control_0_dataflow_b;
	reg mesh_16_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_27_io_in_control_0_shift_b;
	reg mesh_17_27_io_in_control_0_dataflow_b;
	reg mesh_17_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_27_io_in_control_0_shift_b;
	reg mesh_18_27_io_in_control_0_dataflow_b;
	reg mesh_18_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_27_io_in_control_0_shift_b;
	reg mesh_19_27_io_in_control_0_dataflow_b;
	reg mesh_19_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_27_io_in_control_0_shift_b;
	reg mesh_20_27_io_in_control_0_dataflow_b;
	reg mesh_20_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_27_io_in_control_0_shift_b;
	reg mesh_21_27_io_in_control_0_dataflow_b;
	reg mesh_21_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_27_io_in_control_0_shift_b;
	reg mesh_22_27_io_in_control_0_dataflow_b;
	reg mesh_22_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_27_io_in_control_0_shift_b;
	reg mesh_23_27_io_in_control_0_dataflow_b;
	reg mesh_23_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_27_io_in_control_0_shift_b;
	reg mesh_24_27_io_in_control_0_dataflow_b;
	reg mesh_24_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_27_io_in_control_0_shift_b;
	reg mesh_25_27_io_in_control_0_dataflow_b;
	reg mesh_25_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_27_io_in_control_0_shift_b;
	reg mesh_26_27_io_in_control_0_dataflow_b;
	reg mesh_26_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_27_io_in_control_0_shift_b;
	reg mesh_27_27_io_in_control_0_dataflow_b;
	reg mesh_27_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_27_io_in_control_0_shift_b;
	reg mesh_28_27_io_in_control_0_dataflow_b;
	reg mesh_28_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_27_io_in_control_0_shift_b;
	reg mesh_29_27_io_in_control_0_dataflow_b;
	reg mesh_29_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_27_io_in_control_0_shift_b;
	reg mesh_30_27_io_in_control_0_dataflow_b;
	reg mesh_30_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_27_io_in_control_0_shift_b;
	reg mesh_31_27_io_in_control_0_dataflow_b;
	reg mesh_31_27_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_28_io_in_control_0_shift_b;
	reg mesh_0_28_io_in_control_0_dataflow_b;
	reg mesh_0_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_28_io_in_control_0_shift_b;
	reg mesh_1_28_io_in_control_0_dataflow_b;
	reg mesh_1_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_28_io_in_control_0_shift_b;
	reg mesh_2_28_io_in_control_0_dataflow_b;
	reg mesh_2_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_28_io_in_control_0_shift_b;
	reg mesh_3_28_io_in_control_0_dataflow_b;
	reg mesh_3_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_28_io_in_control_0_shift_b;
	reg mesh_4_28_io_in_control_0_dataflow_b;
	reg mesh_4_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_28_io_in_control_0_shift_b;
	reg mesh_5_28_io_in_control_0_dataflow_b;
	reg mesh_5_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_28_io_in_control_0_shift_b;
	reg mesh_6_28_io_in_control_0_dataflow_b;
	reg mesh_6_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_28_io_in_control_0_shift_b;
	reg mesh_7_28_io_in_control_0_dataflow_b;
	reg mesh_7_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_28_io_in_control_0_shift_b;
	reg mesh_8_28_io_in_control_0_dataflow_b;
	reg mesh_8_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_28_io_in_control_0_shift_b;
	reg mesh_9_28_io_in_control_0_dataflow_b;
	reg mesh_9_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_28_io_in_control_0_shift_b;
	reg mesh_10_28_io_in_control_0_dataflow_b;
	reg mesh_10_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_28_io_in_control_0_shift_b;
	reg mesh_11_28_io_in_control_0_dataflow_b;
	reg mesh_11_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_28_io_in_control_0_shift_b;
	reg mesh_12_28_io_in_control_0_dataflow_b;
	reg mesh_12_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_28_io_in_control_0_shift_b;
	reg mesh_13_28_io_in_control_0_dataflow_b;
	reg mesh_13_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_28_io_in_control_0_shift_b;
	reg mesh_14_28_io_in_control_0_dataflow_b;
	reg mesh_14_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_28_io_in_control_0_shift_b;
	reg mesh_15_28_io_in_control_0_dataflow_b;
	reg mesh_15_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_28_io_in_control_0_shift_b;
	reg mesh_16_28_io_in_control_0_dataflow_b;
	reg mesh_16_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_28_io_in_control_0_shift_b;
	reg mesh_17_28_io_in_control_0_dataflow_b;
	reg mesh_17_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_28_io_in_control_0_shift_b;
	reg mesh_18_28_io_in_control_0_dataflow_b;
	reg mesh_18_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_28_io_in_control_0_shift_b;
	reg mesh_19_28_io_in_control_0_dataflow_b;
	reg mesh_19_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_28_io_in_control_0_shift_b;
	reg mesh_20_28_io_in_control_0_dataflow_b;
	reg mesh_20_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_28_io_in_control_0_shift_b;
	reg mesh_21_28_io_in_control_0_dataflow_b;
	reg mesh_21_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_28_io_in_control_0_shift_b;
	reg mesh_22_28_io_in_control_0_dataflow_b;
	reg mesh_22_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_28_io_in_control_0_shift_b;
	reg mesh_23_28_io_in_control_0_dataflow_b;
	reg mesh_23_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_28_io_in_control_0_shift_b;
	reg mesh_24_28_io_in_control_0_dataflow_b;
	reg mesh_24_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_28_io_in_control_0_shift_b;
	reg mesh_25_28_io_in_control_0_dataflow_b;
	reg mesh_25_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_28_io_in_control_0_shift_b;
	reg mesh_26_28_io_in_control_0_dataflow_b;
	reg mesh_26_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_28_io_in_control_0_shift_b;
	reg mesh_27_28_io_in_control_0_dataflow_b;
	reg mesh_27_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_28_io_in_control_0_shift_b;
	reg mesh_28_28_io_in_control_0_dataflow_b;
	reg mesh_28_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_28_io_in_control_0_shift_b;
	reg mesh_29_28_io_in_control_0_dataflow_b;
	reg mesh_29_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_28_io_in_control_0_shift_b;
	reg mesh_30_28_io_in_control_0_dataflow_b;
	reg mesh_30_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_28_io_in_control_0_shift_b;
	reg mesh_31_28_io_in_control_0_dataflow_b;
	reg mesh_31_28_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_29_io_in_control_0_shift_b;
	reg mesh_0_29_io_in_control_0_dataflow_b;
	reg mesh_0_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_29_io_in_control_0_shift_b;
	reg mesh_1_29_io_in_control_0_dataflow_b;
	reg mesh_1_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_29_io_in_control_0_shift_b;
	reg mesh_2_29_io_in_control_0_dataflow_b;
	reg mesh_2_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_29_io_in_control_0_shift_b;
	reg mesh_3_29_io_in_control_0_dataflow_b;
	reg mesh_3_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_29_io_in_control_0_shift_b;
	reg mesh_4_29_io_in_control_0_dataflow_b;
	reg mesh_4_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_29_io_in_control_0_shift_b;
	reg mesh_5_29_io_in_control_0_dataflow_b;
	reg mesh_5_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_29_io_in_control_0_shift_b;
	reg mesh_6_29_io_in_control_0_dataflow_b;
	reg mesh_6_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_29_io_in_control_0_shift_b;
	reg mesh_7_29_io_in_control_0_dataflow_b;
	reg mesh_7_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_29_io_in_control_0_shift_b;
	reg mesh_8_29_io_in_control_0_dataflow_b;
	reg mesh_8_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_29_io_in_control_0_shift_b;
	reg mesh_9_29_io_in_control_0_dataflow_b;
	reg mesh_9_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_29_io_in_control_0_shift_b;
	reg mesh_10_29_io_in_control_0_dataflow_b;
	reg mesh_10_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_29_io_in_control_0_shift_b;
	reg mesh_11_29_io_in_control_0_dataflow_b;
	reg mesh_11_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_29_io_in_control_0_shift_b;
	reg mesh_12_29_io_in_control_0_dataflow_b;
	reg mesh_12_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_29_io_in_control_0_shift_b;
	reg mesh_13_29_io_in_control_0_dataflow_b;
	reg mesh_13_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_29_io_in_control_0_shift_b;
	reg mesh_14_29_io_in_control_0_dataflow_b;
	reg mesh_14_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_29_io_in_control_0_shift_b;
	reg mesh_15_29_io_in_control_0_dataflow_b;
	reg mesh_15_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_29_io_in_control_0_shift_b;
	reg mesh_16_29_io_in_control_0_dataflow_b;
	reg mesh_16_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_29_io_in_control_0_shift_b;
	reg mesh_17_29_io_in_control_0_dataflow_b;
	reg mesh_17_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_29_io_in_control_0_shift_b;
	reg mesh_18_29_io_in_control_0_dataflow_b;
	reg mesh_18_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_29_io_in_control_0_shift_b;
	reg mesh_19_29_io_in_control_0_dataflow_b;
	reg mesh_19_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_29_io_in_control_0_shift_b;
	reg mesh_20_29_io_in_control_0_dataflow_b;
	reg mesh_20_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_29_io_in_control_0_shift_b;
	reg mesh_21_29_io_in_control_0_dataflow_b;
	reg mesh_21_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_29_io_in_control_0_shift_b;
	reg mesh_22_29_io_in_control_0_dataflow_b;
	reg mesh_22_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_29_io_in_control_0_shift_b;
	reg mesh_23_29_io_in_control_0_dataflow_b;
	reg mesh_23_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_29_io_in_control_0_shift_b;
	reg mesh_24_29_io_in_control_0_dataflow_b;
	reg mesh_24_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_29_io_in_control_0_shift_b;
	reg mesh_25_29_io_in_control_0_dataflow_b;
	reg mesh_25_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_29_io_in_control_0_shift_b;
	reg mesh_26_29_io_in_control_0_dataflow_b;
	reg mesh_26_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_29_io_in_control_0_shift_b;
	reg mesh_27_29_io_in_control_0_dataflow_b;
	reg mesh_27_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_29_io_in_control_0_shift_b;
	reg mesh_28_29_io_in_control_0_dataflow_b;
	reg mesh_28_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_29_io_in_control_0_shift_b;
	reg mesh_29_29_io_in_control_0_dataflow_b;
	reg mesh_29_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_29_io_in_control_0_shift_b;
	reg mesh_30_29_io_in_control_0_dataflow_b;
	reg mesh_30_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_29_io_in_control_0_shift_b;
	reg mesh_31_29_io_in_control_0_dataflow_b;
	reg mesh_31_29_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_30_io_in_control_0_shift_b;
	reg mesh_0_30_io_in_control_0_dataflow_b;
	reg mesh_0_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_30_io_in_control_0_shift_b;
	reg mesh_1_30_io_in_control_0_dataflow_b;
	reg mesh_1_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_30_io_in_control_0_shift_b;
	reg mesh_2_30_io_in_control_0_dataflow_b;
	reg mesh_2_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_30_io_in_control_0_shift_b;
	reg mesh_3_30_io_in_control_0_dataflow_b;
	reg mesh_3_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_30_io_in_control_0_shift_b;
	reg mesh_4_30_io_in_control_0_dataflow_b;
	reg mesh_4_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_30_io_in_control_0_shift_b;
	reg mesh_5_30_io_in_control_0_dataflow_b;
	reg mesh_5_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_30_io_in_control_0_shift_b;
	reg mesh_6_30_io_in_control_0_dataflow_b;
	reg mesh_6_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_30_io_in_control_0_shift_b;
	reg mesh_7_30_io_in_control_0_dataflow_b;
	reg mesh_7_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_30_io_in_control_0_shift_b;
	reg mesh_8_30_io_in_control_0_dataflow_b;
	reg mesh_8_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_30_io_in_control_0_shift_b;
	reg mesh_9_30_io_in_control_0_dataflow_b;
	reg mesh_9_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_30_io_in_control_0_shift_b;
	reg mesh_10_30_io_in_control_0_dataflow_b;
	reg mesh_10_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_30_io_in_control_0_shift_b;
	reg mesh_11_30_io_in_control_0_dataflow_b;
	reg mesh_11_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_30_io_in_control_0_shift_b;
	reg mesh_12_30_io_in_control_0_dataflow_b;
	reg mesh_12_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_30_io_in_control_0_shift_b;
	reg mesh_13_30_io_in_control_0_dataflow_b;
	reg mesh_13_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_30_io_in_control_0_shift_b;
	reg mesh_14_30_io_in_control_0_dataflow_b;
	reg mesh_14_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_30_io_in_control_0_shift_b;
	reg mesh_15_30_io_in_control_0_dataflow_b;
	reg mesh_15_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_30_io_in_control_0_shift_b;
	reg mesh_16_30_io_in_control_0_dataflow_b;
	reg mesh_16_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_30_io_in_control_0_shift_b;
	reg mesh_17_30_io_in_control_0_dataflow_b;
	reg mesh_17_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_30_io_in_control_0_shift_b;
	reg mesh_18_30_io_in_control_0_dataflow_b;
	reg mesh_18_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_30_io_in_control_0_shift_b;
	reg mesh_19_30_io_in_control_0_dataflow_b;
	reg mesh_19_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_30_io_in_control_0_shift_b;
	reg mesh_20_30_io_in_control_0_dataflow_b;
	reg mesh_20_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_30_io_in_control_0_shift_b;
	reg mesh_21_30_io_in_control_0_dataflow_b;
	reg mesh_21_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_30_io_in_control_0_shift_b;
	reg mesh_22_30_io_in_control_0_dataflow_b;
	reg mesh_22_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_30_io_in_control_0_shift_b;
	reg mesh_23_30_io_in_control_0_dataflow_b;
	reg mesh_23_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_30_io_in_control_0_shift_b;
	reg mesh_24_30_io_in_control_0_dataflow_b;
	reg mesh_24_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_30_io_in_control_0_shift_b;
	reg mesh_25_30_io_in_control_0_dataflow_b;
	reg mesh_25_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_30_io_in_control_0_shift_b;
	reg mesh_26_30_io_in_control_0_dataflow_b;
	reg mesh_26_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_30_io_in_control_0_shift_b;
	reg mesh_27_30_io_in_control_0_dataflow_b;
	reg mesh_27_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_30_io_in_control_0_shift_b;
	reg mesh_28_30_io_in_control_0_dataflow_b;
	reg mesh_28_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_30_io_in_control_0_shift_b;
	reg mesh_29_30_io_in_control_0_dataflow_b;
	reg mesh_29_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_30_io_in_control_0_shift_b;
	reg mesh_30_30_io_in_control_0_dataflow_b;
	reg mesh_30_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_30_io_in_control_0_shift_b;
	reg mesh_31_30_io_in_control_0_dataflow_b;
	reg mesh_31_30_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_31_io_in_control_0_shift_b;
	reg mesh_0_31_io_in_control_0_dataflow_b;
	reg mesh_0_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_31_io_in_control_0_shift_b;
	reg mesh_1_31_io_in_control_0_dataflow_b;
	reg mesh_1_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_31_io_in_control_0_shift_b;
	reg mesh_2_31_io_in_control_0_dataflow_b;
	reg mesh_2_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_31_io_in_control_0_shift_b;
	reg mesh_3_31_io_in_control_0_dataflow_b;
	reg mesh_3_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_31_io_in_control_0_shift_b;
	reg mesh_4_31_io_in_control_0_dataflow_b;
	reg mesh_4_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_31_io_in_control_0_shift_b;
	reg mesh_5_31_io_in_control_0_dataflow_b;
	reg mesh_5_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_31_io_in_control_0_shift_b;
	reg mesh_6_31_io_in_control_0_dataflow_b;
	reg mesh_6_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_31_io_in_control_0_shift_b;
	reg mesh_7_31_io_in_control_0_dataflow_b;
	reg mesh_7_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_8_31_io_in_control_0_shift_b;
	reg mesh_8_31_io_in_control_0_dataflow_b;
	reg mesh_8_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_9_31_io_in_control_0_shift_b;
	reg mesh_9_31_io_in_control_0_dataflow_b;
	reg mesh_9_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_10_31_io_in_control_0_shift_b;
	reg mesh_10_31_io_in_control_0_dataflow_b;
	reg mesh_10_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_11_31_io_in_control_0_shift_b;
	reg mesh_11_31_io_in_control_0_dataflow_b;
	reg mesh_11_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_12_31_io_in_control_0_shift_b;
	reg mesh_12_31_io_in_control_0_dataflow_b;
	reg mesh_12_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_13_31_io_in_control_0_shift_b;
	reg mesh_13_31_io_in_control_0_dataflow_b;
	reg mesh_13_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_14_31_io_in_control_0_shift_b;
	reg mesh_14_31_io_in_control_0_dataflow_b;
	reg mesh_14_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_15_31_io_in_control_0_shift_b;
	reg mesh_15_31_io_in_control_0_dataflow_b;
	reg mesh_15_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_16_31_io_in_control_0_shift_b;
	reg mesh_16_31_io_in_control_0_dataflow_b;
	reg mesh_16_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_17_31_io_in_control_0_shift_b;
	reg mesh_17_31_io_in_control_0_dataflow_b;
	reg mesh_17_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_18_31_io_in_control_0_shift_b;
	reg mesh_18_31_io_in_control_0_dataflow_b;
	reg mesh_18_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_19_31_io_in_control_0_shift_b;
	reg mesh_19_31_io_in_control_0_dataflow_b;
	reg mesh_19_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_20_31_io_in_control_0_shift_b;
	reg mesh_20_31_io_in_control_0_dataflow_b;
	reg mesh_20_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_21_31_io_in_control_0_shift_b;
	reg mesh_21_31_io_in_control_0_dataflow_b;
	reg mesh_21_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_22_31_io_in_control_0_shift_b;
	reg mesh_22_31_io_in_control_0_dataflow_b;
	reg mesh_22_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_23_31_io_in_control_0_shift_b;
	reg mesh_23_31_io_in_control_0_dataflow_b;
	reg mesh_23_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_24_31_io_in_control_0_shift_b;
	reg mesh_24_31_io_in_control_0_dataflow_b;
	reg mesh_24_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_25_31_io_in_control_0_shift_b;
	reg mesh_25_31_io_in_control_0_dataflow_b;
	reg mesh_25_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_26_31_io_in_control_0_shift_b;
	reg mesh_26_31_io_in_control_0_dataflow_b;
	reg mesh_26_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_27_31_io_in_control_0_shift_b;
	reg mesh_27_31_io_in_control_0_dataflow_b;
	reg mesh_27_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_28_31_io_in_control_0_shift_b;
	reg mesh_28_31_io_in_control_0_dataflow_b;
	reg mesh_28_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_29_31_io_in_control_0_shift_b;
	reg mesh_29_31_io_in_control_0_dataflow_b;
	reg mesh_29_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_30_31_io_in_control_0_shift_b;
	reg mesh_30_31_io_in_control_0_dataflow_b;
	reg mesh_30_31_io_in_control_0_propagate_b;
	reg [4:0] mesh_31_31_io_in_control_0_shift_b;
	reg mesh_31_31_io_in_control_0_dataflow_b;
	reg mesh_31_31_io_in_control_0_propagate_b;
	reg r_1024_0;
	reg r_1025_0;
	reg r_1026_0;
	reg r_1027_0;
	reg r_1028_0;
	reg r_1029_0;
	reg r_1030_0;
	reg r_1031_0;
	reg r_1032_0;
	reg r_1033_0;
	reg r_1034_0;
	reg r_1035_0;
	reg r_1036_0;
	reg r_1037_0;
	reg r_1038_0;
	reg r_1039_0;
	reg r_1040_0;
	reg r_1041_0;
	reg r_1042_0;
	reg r_1043_0;
	reg r_1044_0;
	reg r_1045_0;
	reg r_1046_0;
	reg r_1047_0;
	reg r_1048_0;
	reg r_1049_0;
	reg r_1050_0;
	reg r_1051_0;
	reg r_1052_0;
	reg r_1053_0;
	reg r_1054_0;
	reg r_1055_0;
	reg r_1056_0;
	reg r_1057_0;
	reg r_1058_0;
	reg r_1059_0;
	reg r_1060_0;
	reg r_1061_0;
	reg r_1062_0;
	reg r_1063_0;
	reg r_1064_0;
	reg r_1065_0;
	reg r_1066_0;
	reg r_1067_0;
	reg r_1068_0;
	reg r_1069_0;
	reg r_1070_0;
	reg r_1071_0;
	reg r_1072_0;
	reg r_1073_0;
	reg r_1074_0;
	reg r_1075_0;
	reg r_1076_0;
	reg r_1077_0;
	reg r_1078_0;
	reg r_1079_0;
	reg r_1080_0;
	reg r_1081_0;
	reg r_1082_0;
	reg r_1083_0;
	reg r_1084_0;
	reg r_1085_0;
	reg r_1086_0;
	reg r_1087_0;
	reg r_1088_0;
	reg r_1089_0;
	reg r_1090_0;
	reg r_1091_0;
	reg r_1092_0;
	reg r_1093_0;
	reg r_1094_0;
	reg r_1095_0;
	reg r_1096_0;
	reg r_1097_0;
	reg r_1098_0;
	reg r_1099_0;
	reg r_1100_0;
	reg r_1101_0;
	reg r_1102_0;
	reg r_1103_0;
	reg r_1104_0;
	reg r_1105_0;
	reg r_1106_0;
	reg r_1107_0;
	reg r_1108_0;
	reg r_1109_0;
	reg r_1110_0;
	reg r_1111_0;
	reg r_1112_0;
	reg r_1113_0;
	reg r_1114_0;
	reg r_1115_0;
	reg r_1116_0;
	reg r_1117_0;
	reg r_1118_0;
	reg r_1119_0;
	reg r_1120_0;
	reg r_1121_0;
	reg r_1122_0;
	reg r_1123_0;
	reg r_1124_0;
	reg r_1125_0;
	reg r_1126_0;
	reg r_1127_0;
	reg r_1128_0;
	reg r_1129_0;
	reg r_1130_0;
	reg r_1131_0;
	reg r_1132_0;
	reg r_1133_0;
	reg r_1134_0;
	reg r_1135_0;
	reg r_1136_0;
	reg r_1137_0;
	reg r_1138_0;
	reg r_1139_0;
	reg r_1140_0;
	reg r_1141_0;
	reg r_1142_0;
	reg r_1143_0;
	reg r_1144_0;
	reg r_1145_0;
	reg r_1146_0;
	reg r_1147_0;
	reg r_1148_0;
	reg r_1149_0;
	reg r_1150_0;
	reg r_1151_0;
	reg r_1152_0;
	reg r_1153_0;
	reg r_1154_0;
	reg r_1155_0;
	reg r_1156_0;
	reg r_1157_0;
	reg r_1158_0;
	reg r_1159_0;
	reg r_1160_0;
	reg r_1161_0;
	reg r_1162_0;
	reg r_1163_0;
	reg r_1164_0;
	reg r_1165_0;
	reg r_1166_0;
	reg r_1167_0;
	reg r_1168_0;
	reg r_1169_0;
	reg r_1170_0;
	reg r_1171_0;
	reg r_1172_0;
	reg r_1173_0;
	reg r_1174_0;
	reg r_1175_0;
	reg r_1176_0;
	reg r_1177_0;
	reg r_1178_0;
	reg r_1179_0;
	reg r_1180_0;
	reg r_1181_0;
	reg r_1182_0;
	reg r_1183_0;
	reg r_1184_0;
	reg r_1185_0;
	reg r_1186_0;
	reg r_1187_0;
	reg r_1188_0;
	reg r_1189_0;
	reg r_1190_0;
	reg r_1191_0;
	reg r_1192_0;
	reg r_1193_0;
	reg r_1194_0;
	reg r_1195_0;
	reg r_1196_0;
	reg r_1197_0;
	reg r_1198_0;
	reg r_1199_0;
	reg r_1200_0;
	reg r_1201_0;
	reg r_1202_0;
	reg r_1203_0;
	reg r_1204_0;
	reg r_1205_0;
	reg r_1206_0;
	reg r_1207_0;
	reg r_1208_0;
	reg r_1209_0;
	reg r_1210_0;
	reg r_1211_0;
	reg r_1212_0;
	reg r_1213_0;
	reg r_1214_0;
	reg r_1215_0;
	reg r_1216_0;
	reg r_1217_0;
	reg r_1218_0;
	reg r_1219_0;
	reg r_1220_0;
	reg r_1221_0;
	reg r_1222_0;
	reg r_1223_0;
	reg r_1224_0;
	reg r_1225_0;
	reg r_1226_0;
	reg r_1227_0;
	reg r_1228_0;
	reg r_1229_0;
	reg r_1230_0;
	reg r_1231_0;
	reg r_1232_0;
	reg r_1233_0;
	reg r_1234_0;
	reg r_1235_0;
	reg r_1236_0;
	reg r_1237_0;
	reg r_1238_0;
	reg r_1239_0;
	reg r_1240_0;
	reg r_1241_0;
	reg r_1242_0;
	reg r_1243_0;
	reg r_1244_0;
	reg r_1245_0;
	reg r_1246_0;
	reg r_1247_0;
	reg r_1248_0;
	reg r_1249_0;
	reg r_1250_0;
	reg r_1251_0;
	reg r_1252_0;
	reg r_1253_0;
	reg r_1254_0;
	reg r_1255_0;
	reg r_1256_0;
	reg r_1257_0;
	reg r_1258_0;
	reg r_1259_0;
	reg r_1260_0;
	reg r_1261_0;
	reg r_1262_0;
	reg r_1263_0;
	reg r_1264_0;
	reg r_1265_0;
	reg r_1266_0;
	reg r_1267_0;
	reg r_1268_0;
	reg r_1269_0;
	reg r_1270_0;
	reg r_1271_0;
	reg r_1272_0;
	reg r_1273_0;
	reg r_1274_0;
	reg r_1275_0;
	reg r_1276_0;
	reg r_1277_0;
	reg r_1278_0;
	reg r_1279_0;
	reg r_1280_0;
	reg r_1281_0;
	reg r_1282_0;
	reg r_1283_0;
	reg r_1284_0;
	reg r_1285_0;
	reg r_1286_0;
	reg r_1287_0;
	reg r_1288_0;
	reg r_1289_0;
	reg r_1290_0;
	reg r_1291_0;
	reg r_1292_0;
	reg r_1293_0;
	reg r_1294_0;
	reg r_1295_0;
	reg r_1296_0;
	reg r_1297_0;
	reg r_1298_0;
	reg r_1299_0;
	reg r_1300_0;
	reg r_1301_0;
	reg r_1302_0;
	reg r_1303_0;
	reg r_1304_0;
	reg r_1305_0;
	reg r_1306_0;
	reg r_1307_0;
	reg r_1308_0;
	reg r_1309_0;
	reg r_1310_0;
	reg r_1311_0;
	reg r_1312_0;
	reg r_1313_0;
	reg r_1314_0;
	reg r_1315_0;
	reg r_1316_0;
	reg r_1317_0;
	reg r_1318_0;
	reg r_1319_0;
	reg r_1320_0;
	reg r_1321_0;
	reg r_1322_0;
	reg r_1323_0;
	reg r_1324_0;
	reg r_1325_0;
	reg r_1326_0;
	reg r_1327_0;
	reg r_1328_0;
	reg r_1329_0;
	reg r_1330_0;
	reg r_1331_0;
	reg r_1332_0;
	reg r_1333_0;
	reg r_1334_0;
	reg r_1335_0;
	reg r_1336_0;
	reg r_1337_0;
	reg r_1338_0;
	reg r_1339_0;
	reg r_1340_0;
	reg r_1341_0;
	reg r_1342_0;
	reg r_1343_0;
	reg r_1344_0;
	reg r_1345_0;
	reg r_1346_0;
	reg r_1347_0;
	reg r_1348_0;
	reg r_1349_0;
	reg r_1350_0;
	reg r_1351_0;
	reg r_1352_0;
	reg r_1353_0;
	reg r_1354_0;
	reg r_1355_0;
	reg r_1356_0;
	reg r_1357_0;
	reg r_1358_0;
	reg r_1359_0;
	reg r_1360_0;
	reg r_1361_0;
	reg r_1362_0;
	reg r_1363_0;
	reg r_1364_0;
	reg r_1365_0;
	reg r_1366_0;
	reg r_1367_0;
	reg r_1368_0;
	reg r_1369_0;
	reg r_1370_0;
	reg r_1371_0;
	reg r_1372_0;
	reg r_1373_0;
	reg r_1374_0;
	reg r_1375_0;
	reg r_1376_0;
	reg r_1377_0;
	reg r_1378_0;
	reg r_1379_0;
	reg r_1380_0;
	reg r_1381_0;
	reg r_1382_0;
	reg r_1383_0;
	reg r_1384_0;
	reg r_1385_0;
	reg r_1386_0;
	reg r_1387_0;
	reg r_1388_0;
	reg r_1389_0;
	reg r_1390_0;
	reg r_1391_0;
	reg r_1392_0;
	reg r_1393_0;
	reg r_1394_0;
	reg r_1395_0;
	reg r_1396_0;
	reg r_1397_0;
	reg r_1398_0;
	reg r_1399_0;
	reg r_1400_0;
	reg r_1401_0;
	reg r_1402_0;
	reg r_1403_0;
	reg r_1404_0;
	reg r_1405_0;
	reg r_1406_0;
	reg r_1407_0;
	reg r_1408_0;
	reg r_1409_0;
	reg r_1410_0;
	reg r_1411_0;
	reg r_1412_0;
	reg r_1413_0;
	reg r_1414_0;
	reg r_1415_0;
	reg r_1416_0;
	reg r_1417_0;
	reg r_1418_0;
	reg r_1419_0;
	reg r_1420_0;
	reg r_1421_0;
	reg r_1422_0;
	reg r_1423_0;
	reg r_1424_0;
	reg r_1425_0;
	reg r_1426_0;
	reg r_1427_0;
	reg r_1428_0;
	reg r_1429_0;
	reg r_1430_0;
	reg r_1431_0;
	reg r_1432_0;
	reg r_1433_0;
	reg r_1434_0;
	reg r_1435_0;
	reg r_1436_0;
	reg r_1437_0;
	reg r_1438_0;
	reg r_1439_0;
	reg r_1440_0;
	reg r_1441_0;
	reg r_1442_0;
	reg r_1443_0;
	reg r_1444_0;
	reg r_1445_0;
	reg r_1446_0;
	reg r_1447_0;
	reg r_1448_0;
	reg r_1449_0;
	reg r_1450_0;
	reg r_1451_0;
	reg r_1452_0;
	reg r_1453_0;
	reg r_1454_0;
	reg r_1455_0;
	reg r_1456_0;
	reg r_1457_0;
	reg r_1458_0;
	reg r_1459_0;
	reg r_1460_0;
	reg r_1461_0;
	reg r_1462_0;
	reg r_1463_0;
	reg r_1464_0;
	reg r_1465_0;
	reg r_1466_0;
	reg r_1467_0;
	reg r_1468_0;
	reg r_1469_0;
	reg r_1470_0;
	reg r_1471_0;
	reg r_1472_0;
	reg r_1473_0;
	reg r_1474_0;
	reg r_1475_0;
	reg r_1476_0;
	reg r_1477_0;
	reg r_1478_0;
	reg r_1479_0;
	reg r_1480_0;
	reg r_1481_0;
	reg r_1482_0;
	reg r_1483_0;
	reg r_1484_0;
	reg r_1485_0;
	reg r_1486_0;
	reg r_1487_0;
	reg r_1488_0;
	reg r_1489_0;
	reg r_1490_0;
	reg r_1491_0;
	reg r_1492_0;
	reg r_1493_0;
	reg r_1494_0;
	reg r_1495_0;
	reg r_1496_0;
	reg r_1497_0;
	reg r_1498_0;
	reg r_1499_0;
	reg r_1500_0;
	reg r_1501_0;
	reg r_1502_0;
	reg r_1503_0;
	reg r_1504_0;
	reg r_1505_0;
	reg r_1506_0;
	reg r_1507_0;
	reg r_1508_0;
	reg r_1509_0;
	reg r_1510_0;
	reg r_1511_0;
	reg r_1512_0;
	reg r_1513_0;
	reg r_1514_0;
	reg r_1515_0;
	reg r_1516_0;
	reg r_1517_0;
	reg r_1518_0;
	reg r_1519_0;
	reg r_1520_0;
	reg r_1521_0;
	reg r_1522_0;
	reg r_1523_0;
	reg r_1524_0;
	reg r_1525_0;
	reg r_1526_0;
	reg r_1527_0;
	reg r_1528_0;
	reg r_1529_0;
	reg r_1530_0;
	reg r_1531_0;
	reg r_1532_0;
	reg r_1533_0;
	reg r_1534_0;
	reg r_1535_0;
	reg r_1536_0;
	reg r_1537_0;
	reg r_1538_0;
	reg r_1539_0;
	reg r_1540_0;
	reg r_1541_0;
	reg r_1542_0;
	reg r_1543_0;
	reg r_1544_0;
	reg r_1545_0;
	reg r_1546_0;
	reg r_1547_0;
	reg r_1548_0;
	reg r_1549_0;
	reg r_1550_0;
	reg r_1551_0;
	reg r_1552_0;
	reg r_1553_0;
	reg r_1554_0;
	reg r_1555_0;
	reg r_1556_0;
	reg r_1557_0;
	reg r_1558_0;
	reg r_1559_0;
	reg r_1560_0;
	reg r_1561_0;
	reg r_1562_0;
	reg r_1563_0;
	reg r_1564_0;
	reg r_1565_0;
	reg r_1566_0;
	reg r_1567_0;
	reg r_1568_0;
	reg r_1569_0;
	reg r_1570_0;
	reg r_1571_0;
	reg r_1572_0;
	reg r_1573_0;
	reg r_1574_0;
	reg r_1575_0;
	reg r_1576_0;
	reg r_1577_0;
	reg r_1578_0;
	reg r_1579_0;
	reg r_1580_0;
	reg r_1581_0;
	reg r_1582_0;
	reg r_1583_0;
	reg r_1584_0;
	reg r_1585_0;
	reg r_1586_0;
	reg r_1587_0;
	reg r_1588_0;
	reg r_1589_0;
	reg r_1590_0;
	reg r_1591_0;
	reg r_1592_0;
	reg r_1593_0;
	reg r_1594_0;
	reg r_1595_0;
	reg r_1596_0;
	reg r_1597_0;
	reg r_1598_0;
	reg r_1599_0;
	reg r_1600_0;
	reg r_1601_0;
	reg r_1602_0;
	reg r_1603_0;
	reg r_1604_0;
	reg r_1605_0;
	reg r_1606_0;
	reg r_1607_0;
	reg r_1608_0;
	reg r_1609_0;
	reg r_1610_0;
	reg r_1611_0;
	reg r_1612_0;
	reg r_1613_0;
	reg r_1614_0;
	reg r_1615_0;
	reg r_1616_0;
	reg r_1617_0;
	reg r_1618_0;
	reg r_1619_0;
	reg r_1620_0;
	reg r_1621_0;
	reg r_1622_0;
	reg r_1623_0;
	reg r_1624_0;
	reg r_1625_0;
	reg r_1626_0;
	reg r_1627_0;
	reg r_1628_0;
	reg r_1629_0;
	reg r_1630_0;
	reg r_1631_0;
	reg r_1632_0;
	reg r_1633_0;
	reg r_1634_0;
	reg r_1635_0;
	reg r_1636_0;
	reg r_1637_0;
	reg r_1638_0;
	reg r_1639_0;
	reg r_1640_0;
	reg r_1641_0;
	reg r_1642_0;
	reg r_1643_0;
	reg r_1644_0;
	reg r_1645_0;
	reg r_1646_0;
	reg r_1647_0;
	reg r_1648_0;
	reg r_1649_0;
	reg r_1650_0;
	reg r_1651_0;
	reg r_1652_0;
	reg r_1653_0;
	reg r_1654_0;
	reg r_1655_0;
	reg r_1656_0;
	reg r_1657_0;
	reg r_1658_0;
	reg r_1659_0;
	reg r_1660_0;
	reg r_1661_0;
	reg r_1662_0;
	reg r_1663_0;
	reg r_1664_0;
	reg r_1665_0;
	reg r_1666_0;
	reg r_1667_0;
	reg r_1668_0;
	reg r_1669_0;
	reg r_1670_0;
	reg r_1671_0;
	reg r_1672_0;
	reg r_1673_0;
	reg r_1674_0;
	reg r_1675_0;
	reg r_1676_0;
	reg r_1677_0;
	reg r_1678_0;
	reg r_1679_0;
	reg r_1680_0;
	reg r_1681_0;
	reg r_1682_0;
	reg r_1683_0;
	reg r_1684_0;
	reg r_1685_0;
	reg r_1686_0;
	reg r_1687_0;
	reg r_1688_0;
	reg r_1689_0;
	reg r_1690_0;
	reg r_1691_0;
	reg r_1692_0;
	reg r_1693_0;
	reg r_1694_0;
	reg r_1695_0;
	reg r_1696_0;
	reg r_1697_0;
	reg r_1698_0;
	reg r_1699_0;
	reg r_1700_0;
	reg r_1701_0;
	reg r_1702_0;
	reg r_1703_0;
	reg r_1704_0;
	reg r_1705_0;
	reg r_1706_0;
	reg r_1707_0;
	reg r_1708_0;
	reg r_1709_0;
	reg r_1710_0;
	reg r_1711_0;
	reg r_1712_0;
	reg r_1713_0;
	reg r_1714_0;
	reg r_1715_0;
	reg r_1716_0;
	reg r_1717_0;
	reg r_1718_0;
	reg r_1719_0;
	reg r_1720_0;
	reg r_1721_0;
	reg r_1722_0;
	reg r_1723_0;
	reg r_1724_0;
	reg r_1725_0;
	reg r_1726_0;
	reg r_1727_0;
	reg r_1728_0;
	reg r_1729_0;
	reg r_1730_0;
	reg r_1731_0;
	reg r_1732_0;
	reg r_1733_0;
	reg r_1734_0;
	reg r_1735_0;
	reg r_1736_0;
	reg r_1737_0;
	reg r_1738_0;
	reg r_1739_0;
	reg r_1740_0;
	reg r_1741_0;
	reg r_1742_0;
	reg r_1743_0;
	reg r_1744_0;
	reg r_1745_0;
	reg r_1746_0;
	reg r_1747_0;
	reg r_1748_0;
	reg r_1749_0;
	reg r_1750_0;
	reg r_1751_0;
	reg r_1752_0;
	reg r_1753_0;
	reg r_1754_0;
	reg r_1755_0;
	reg r_1756_0;
	reg r_1757_0;
	reg r_1758_0;
	reg r_1759_0;
	reg r_1760_0;
	reg r_1761_0;
	reg r_1762_0;
	reg r_1763_0;
	reg r_1764_0;
	reg r_1765_0;
	reg r_1766_0;
	reg r_1767_0;
	reg r_1768_0;
	reg r_1769_0;
	reg r_1770_0;
	reg r_1771_0;
	reg r_1772_0;
	reg r_1773_0;
	reg r_1774_0;
	reg r_1775_0;
	reg r_1776_0;
	reg r_1777_0;
	reg r_1778_0;
	reg r_1779_0;
	reg r_1780_0;
	reg r_1781_0;
	reg r_1782_0;
	reg r_1783_0;
	reg r_1784_0;
	reg r_1785_0;
	reg r_1786_0;
	reg r_1787_0;
	reg r_1788_0;
	reg r_1789_0;
	reg r_1790_0;
	reg r_1791_0;
	reg r_1792_0;
	reg r_1793_0;
	reg r_1794_0;
	reg r_1795_0;
	reg r_1796_0;
	reg r_1797_0;
	reg r_1798_0;
	reg r_1799_0;
	reg r_1800_0;
	reg r_1801_0;
	reg r_1802_0;
	reg r_1803_0;
	reg r_1804_0;
	reg r_1805_0;
	reg r_1806_0;
	reg r_1807_0;
	reg r_1808_0;
	reg r_1809_0;
	reg r_1810_0;
	reg r_1811_0;
	reg r_1812_0;
	reg r_1813_0;
	reg r_1814_0;
	reg r_1815_0;
	reg r_1816_0;
	reg r_1817_0;
	reg r_1818_0;
	reg r_1819_0;
	reg r_1820_0;
	reg r_1821_0;
	reg r_1822_0;
	reg r_1823_0;
	reg r_1824_0;
	reg r_1825_0;
	reg r_1826_0;
	reg r_1827_0;
	reg r_1828_0;
	reg r_1829_0;
	reg r_1830_0;
	reg r_1831_0;
	reg r_1832_0;
	reg r_1833_0;
	reg r_1834_0;
	reg r_1835_0;
	reg r_1836_0;
	reg r_1837_0;
	reg r_1838_0;
	reg r_1839_0;
	reg r_1840_0;
	reg r_1841_0;
	reg r_1842_0;
	reg r_1843_0;
	reg r_1844_0;
	reg r_1845_0;
	reg r_1846_0;
	reg r_1847_0;
	reg r_1848_0;
	reg r_1849_0;
	reg r_1850_0;
	reg r_1851_0;
	reg r_1852_0;
	reg r_1853_0;
	reg r_1854_0;
	reg r_1855_0;
	reg r_1856_0;
	reg r_1857_0;
	reg r_1858_0;
	reg r_1859_0;
	reg r_1860_0;
	reg r_1861_0;
	reg r_1862_0;
	reg r_1863_0;
	reg r_1864_0;
	reg r_1865_0;
	reg r_1866_0;
	reg r_1867_0;
	reg r_1868_0;
	reg r_1869_0;
	reg r_1870_0;
	reg r_1871_0;
	reg r_1872_0;
	reg r_1873_0;
	reg r_1874_0;
	reg r_1875_0;
	reg r_1876_0;
	reg r_1877_0;
	reg r_1878_0;
	reg r_1879_0;
	reg r_1880_0;
	reg r_1881_0;
	reg r_1882_0;
	reg r_1883_0;
	reg r_1884_0;
	reg r_1885_0;
	reg r_1886_0;
	reg r_1887_0;
	reg r_1888_0;
	reg r_1889_0;
	reg r_1890_0;
	reg r_1891_0;
	reg r_1892_0;
	reg r_1893_0;
	reg r_1894_0;
	reg r_1895_0;
	reg r_1896_0;
	reg r_1897_0;
	reg r_1898_0;
	reg r_1899_0;
	reg r_1900_0;
	reg r_1901_0;
	reg r_1902_0;
	reg r_1903_0;
	reg r_1904_0;
	reg r_1905_0;
	reg r_1906_0;
	reg r_1907_0;
	reg r_1908_0;
	reg r_1909_0;
	reg r_1910_0;
	reg r_1911_0;
	reg r_1912_0;
	reg r_1913_0;
	reg r_1914_0;
	reg r_1915_0;
	reg r_1916_0;
	reg r_1917_0;
	reg r_1918_0;
	reg r_1919_0;
	reg r_1920_0;
	reg r_1921_0;
	reg r_1922_0;
	reg r_1923_0;
	reg r_1924_0;
	reg r_1925_0;
	reg r_1926_0;
	reg r_1927_0;
	reg r_1928_0;
	reg r_1929_0;
	reg r_1930_0;
	reg r_1931_0;
	reg r_1932_0;
	reg r_1933_0;
	reg r_1934_0;
	reg r_1935_0;
	reg r_1936_0;
	reg r_1937_0;
	reg r_1938_0;
	reg r_1939_0;
	reg r_1940_0;
	reg r_1941_0;
	reg r_1942_0;
	reg r_1943_0;
	reg r_1944_0;
	reg r_1945_0;
	reg r_1946_0;
	reg r_1947_0;
	reg r_1948_0;
	reg r_1949_0;
	reg r_1950_0;
	reg r_1951_0;
	reg r_1952_0;
	reg r_1953_0;
	reg r_1954_0;
	reg r_1955_0;
	reg r_1956_0;
	reg r_1957_0;
	reg r_1958_0;
	reg r_1959_0;
	reg r_1960_0;
	reg r_1961_0;
	reg r_1962_0;
	reg r_1963_0;
	reg r_1964_0;
	reg r_1965_0;
	reg r_1966_0;
	reg r_1967_0;
	reg r_1968_0;
	reg r_1969_0;
	reg r_1970_0;
	reg r_1971_0;
	reg r_1972_0;
	reg r_1973_0;
	reg r_1974_0;
	reg r_1975_0;
	reg r_1976_0;
	reg r_1977_0;
	reg r_1978_0;
	reg r_1979_0;
	reg r_1980_0;
	reg r_1981_0;
	reg r_1982_0;
	reg r_1983_0;
	reg r_1984_0;
	reg r_1985_0;
	reg r_1986_0;
	reg r_1987_0;
	reg r_1988_0;
	reg r_1989_0;
	reg r_1990_0;
	reg r_1991_0;
	reg r_1992_0;
	reg r_1993_0;
	reg r_1994_0;
	reg r_1995_0;
	reg r_1996_0;
	reg r_1997_0;
	reg r_1998_0;
	reg r_1999_0;
	reg r_2000_0;
	reg r_2001_0;
	reg r_2002_0;
	reg r_2003_0;
	reg r_2004_0;
	reg r_2005_0;
	reg r_2006_0;
	reg r_2007_0;
	reg r_2008_0;
	reg r_2009_0;
	reg r_2010_0;
	reg r_2011_0;
	reg r_2012_0;
	reg r_2013_0;
	reg r_2014_0;
	reg r_2015_0;
	reg r_2016_0;
	reg r_2017_0;
	reg r_2018_0;
	reg r_2019_0;
	reg r_2020_0;
	reg r_2021_0;
	reg r_2022_0;
	reg r_2023_0;
	reg r_2024_0;
	reg r_2025_0;
	reg r_2026_0;
	reg r_2027_0;
	reg r_2028_0;
	reg r_2029_0;
	reg r_2030_0;
	reg r_2031_0;
	reg r_2032_0;
	reg r_2033_0;
	reg r_2034_0;
	reg r_2035_0;
	reg r_2036_0;
	reg r_2037_0;
	reg r_2038_0;
	reg r_2039_0;
	reg r_2040_0;
	reg r_2041_0;
	reg r_2042_0;
	reg r_2043_0;
	reg r_2044_0;
	reg r_2045_0;
	reg r_2046_0;
	reg r_2047_0;
	reg [2:0] r_2048_0;
	reg [2:0] r_2049_0;
	reg [2:0] r_2050_0;
	reg [2:0] r_2051_0;
	reg [2:0] r_2052_0;
	reg [2:0] r_2053_0;
	reg [2:0] r_2054_0;
	reg [2:0] r_2055_0;
	reg [2:0] r_2056_0;
	reg [2:0] r_2057_0;
	reg [2:0] r_2058_0;
	reg [2:0] r_2059_0;
	reg [2:0] r_2060_0;
	reg [2:0] r_2061_0;
	reg [2:0] r_2062_0;
	reg [2:0] r_2063_0;
	reg [2:0] r_2064_0;
	reg [2:0] r_2065_0;
	reg [2:0] r_2066_0;
	reg [2:0] r_2067_0;
	reg [2:0] r_2068_0;
	reg [2:0] r_2069_0;
	reg [2:0] r_2070_0;
	reg [2:0] r_2071_0;
	reg [2:0] r_2072_0;
	reg [2:0] r_2073_0;
	reg [2:0] r_2074_0;
	reg [2:0] r_2075_0;
	reg [2:0] r_2076_0;
	reg [2:0] r_2077_0;
	reg [2:0] r_2078_0;
	reg [2:0] r_2079_0;
	reg [2:0] r_2080_0;
	reg [2:0] r_2081_0;
	reg [2:0] r_2082_0;
	reg [2:0] r_2083_0;
	reg [2:0] r_2084_0;
	reg [2:0] r_2085_0;
	reg [2:0] r_2086_0;
	reg [2:0] r_2087_0;
	reg [2:0] r_2088_0;
	reg [2:0] r_2089_0;
	reg [2:0] r_2090_0;
	reg [2:0] r_2091_0;
	reg [2:0] r_2092_0;
	reg [2:0] r_2093_0;
	reg [2:0] r_2094_0;
	reg [2:0] r_2095_0;
	reg [2:0] r_2096_0;
	reg [2:0] r_2097_0;
	reg [2:0] r_2098_0;
	reg [2:0] r_2099_0;
	reg [2:0] r_2100_0;
	reg [2:0] r_2101_0;
	reg [2:0] r_2102_0;
	reg [2:0] r_2103_0;
	reg [2:0] r_2104_0;
	reg [2:0] r_2105_0;
	reg [2:0] r_2106_0;
	reg [2:0] r_2107_0;
	reg [2:0] r_2108_0;
	reg [2:0] r_2109_0;
	reg [2:0] r_2110_0;
	reg [2:0] r_2111_0;
	reg [2:0] r_2112_0;
	reg [2:0] r_2113_0;
	reg [2:0] r_2114_0;
	reg [2:0] r_2115_0;
	reg [2:0] r_2116_0;
	reg [2:0] r_2117_0;
	reg [2:0] r_2118_0;
	reg [2:0] r_2119_0;
	reg [2:0] r_2120_0;
	reg [2:0] r_2121_0;
	reg [2:0] r_2122_0;
	reg [2:0] r_2123_0;
	reg [2:0] r_2124_0;
	reg [2:0] r_2125_0;
	reg [2:0] r_2126_0;
	reg [2:0] r_2127_0;
	reg [2:0] r_2128_0;
	reg [2:0] r_2129_0;
	reg [2:0] r_2130_0;
	reg [2:0] r_2131_0;
	reg [2:0] r_2132_0;
	reg [2:0] r_2133_0;
	reg [2:0] r_2134_0;
	reg [2:0] r_2135_0;
	reg [2:0] r_2136_0;
	reg [2:0] r_2137_0;
	reg [2:0] r_2138_0;
	reg [2:0] r_2139_0;
	reg [2:0] r_2140_0;
	reg [2:0] r_2141_0;
	reg [2:0] r_2142_0;
	reg [2:0] r_2143_0;
	reg [2:0] r_2144_0;
	reg [2:0] r_2145_0;
	reg [2:0] r_2146_0;
	reg [2:0] r_2147_0;
	reg [2:0] r_2148_0;
	reg [2:0] r_2149_0;
	reg [2:0] r_2150_0;
	reg [2:0] r_2151_0;
	reg [2:0] r_2152_0;
	reg [2:0] r_2153_0;
	reg [2:0] r_2154_0;
	reg [2:0] r_2155_0;
	reg [2:0] r_2156_0;
	reg [2:0] r_2157_0;
	reg [2:0] r_2158_0;
	reg [2:0] r_2159_0;
	reg [2:0] r_2160_0;
	reg [2:0] r_2161_0;
	reg [2:0] r_2162_0;
	reg [2:0] r_2163_0;
	reg [2:0] r_2164_0;
	reg [2:0] r_2165_0;
	reg [2:0] r_2166_0;
	reg [2:0] r_2167_0;
	reg [2:0] r_2168_0;
	reg [2:0] r_2169_0;
	reg [2:0] r_2170_0;
	reg [2:0] r_2171_0;
	reg [2:0] r_2172_0;
	reg [2:0] r_2173_0;
	reg [2:0] r_2174_0;
	reg [2:0] r_2175_0;
	reg [2:0] r_2176_0;
	reg [2:0] r_2177_0;
	reg [2:0] r_2178_0;
	reg [2:0] r_2179_0;
	reg [2:0] r_2180_0;
	reg [2:0] r_2181_0;
	reg [2:0] r_2182_0;
	reg [2:0] r_2183_0;
	reg [2:0] r_2184_0;
	reg [2:0] r_2185_0;
	reg [2:0] r_2186_0;
	reg [2:0] r_2187_0;
	reg [2:0] r_2188_0;
	reg [2:0] r_2189_0;
	reg [2:0] r_2190_0;
	reg [2:0] r_2191_0;
	reg [2:0] r_2192_0;
	reg [2:0] r_2193_0;
	reg [2:0] r_2194_0;
	reg [2:0] r_2195_0;
	reg [2:0] r_2196_0;
	reg [2:0] r_2197_0;
	reg [2:0] r_2198_0;
	reg [2:0] r_2199_0;
	reg [2:0] r_2200_0;
	reg [2:0] r_2201_0;
	reg [2:0] r_2202_0;
	reg [2:0] r_2203_0;
	reg [2:0] r_2204_0;
	reg [2:0] r_2205_0;
	reg [2:0] r_2206_0;
	reg [2:0] r_2207_0;
	reg [2:0] r_2208_0;
	reg [2:0] r_2209_0;
	reg [2:0] r_2210_0;
	reg [2:0] r_2211_0;
	reg [2:0] r_2212_0;
	reg [2:0] r_2213_0;
	reg [2:0] r_2214_0;
	reg [2:0] r_2215_0;
	reg [2:0] r_2216_0;
	reg [2:0] r_2217_0;
	reg [2:0] r_2218_0;
	reg [2:0] r_2219_0;
	reg [2:0] r_2220_0;
	reg [2:0] r_2221_0;
	reg [2:0] r_2222_0;
	reg [2:0] r_2223_0;
	reg [2:0] r_2224_0;
	reg [2:0] r_2225_0;
	reg [2:0] r_2226_0;
	reg [2:0] r_2227_0;
	reg [2:0] r_2228_0;
	reg [2:0] r_2229_0;
	reg [2:0] r_2230_0;
	reg [2:0] r_2231_0;
	reg [2:0] r_2232_0;
	reg [2:0] r_2233_0;
	reg [2:0] r_2234_0;
	reg [2:0] r_2235_0;
	reg [2:0] r_2236_0;
	reg [2:0] r_2237_0;
	reg [2:0] r_2238_0;
	reg [2:0] r_2239_0;
	reg [2:0] r_2240_0;
	reg [2:0] r_2241_0;
	reg [2:0] r_2242_0;
	reg [2:0] r_2243_0;
	reg [2:0] r_2244_0;
	reg [2:0] r_2245_0;
	reg [2:0] r_2246_0;
	reg [2:0] r_2247_0;
	reg [2:0] r_2248_0;
	reg [2:0] r_2249_0;
	reg [2:0] r_2250_0;
	reg [2:0] r_2251_0;
	reg [2:0] r_2252_0;
	reg [2:0] r_2253_0;
	reg [2:0] r_2254_0;
	reg [2:0] r_2255_0;
	reg [2:0] r_2256_0;
	reg [2:0] r_2257_0;
	reg [2:0] r_2258_0;
	reg [2:0] r_2259_0;
	reg [2:0] r_2260_0;
	reg [2:0] r_2261_0;
	reg [2:0] r_2262_0;
	reg [2:0] r_2263_0;
	reg [2:0] r_2264_0;
	reg [2:0] r_2265_0;
	reg [2:0] r_2266_0;
	reg [2:0] r_2267_0;
	reg [2:0] r_2268_0;
	reg [2:0] r_2269_0;
	reg [2:0] r_2270_0;
	reg [2:0] r_2271_0;
	reg [2:0] r_2272_0;
	reg [2:0] r_2273_0;
	reg [2:0] r_2274_0;
	reg [2:0] r_2275_0;
	reg [2:0] r_2276_0;
	reg [2:0] r_2277_0;
	reg [2:0] r_2278_0;
	reg [2:0] r_2279_0;
	reg [2:0] r_2280_0;
	reg [2:0] r_2281_0;
	reg [2:0] r_2282_0;
	reg [2:0] r_2283_0;
	reg [2:0] r_2284_0;
	reg [2:0] r_2285_0;
	reg [2:0] r_2286_0;
	reg [2:0] r_2287_0;
	reg [2:0] r_2288_0;
	reg [2:0] r_2289_0;
	reg [2:0] r_2290_0;
	reg [2:0] r_2291_0;
	reg [2:0] r_2292_0;
	reg [2:0] r_2293_0;
	reg [2:0] r_2294_0;
	reg [2:0] r_2295_0;
	reg [2:0] r_2296_0;
	reg [2:0] r_2297_0;
	reg [2:0] r_2298_0;
	reg [2:0] r_2299_0;
	reg [2:0] r_2300_0;
	reg [2:0] r_2301_0;
	reg [2:0] r_2302_0;
	reg [2:0] r_2303_0;
	reg [2:0] r_2304_0;
	reg [2:0] r_2305_0;
	reg [2:0] r_2306_0;
	reg [2:0] r_2307_0;
	reg [2:0] r_2308_0;
	reg [2:0] r_2309_0;
	reg [2:0] r_2310_0;
	reg [2:0] r_2311_0;
	reg [2:0] r_2312_0;
	reg [2:0] r_2313_0;
	reg [2:0] r_2314_0;
	reg [2:0] r_2315_0;
	reg [2:0] r_2316_0;
	reg [2:0] r_2317_0;
	reg [2:0] r_2318_0;
	reg [2:0] r_2319_0;
	reg [2:0] r_2320_0;
	reg [2:0] r_2321_0;
	reg [2:0] r_2322_0;
	reg [2:0] r_2323_0;
	reg [2:0] r_2324_0;
	reg [2:0] r_2325_0;
	reg [2:0] r_2326_0;
	reg [2:0] r_2327_0;
	reg [2:0] r_2328_0;
	reg [2:0] r_2329_0;
	reg [2:0] r_2330_0;
	reg [2:0] r_2331_0;
	reg [2:0] r_2332_0;
	reg [2:0] r_2333_0;
	reg [2:0] r_2334_0;
	reg [2:0] r_2335_0;
	reg [2:0] r_2336_0;
	reg [2:0] r_2337_0;
	reg [2:0] r_2338_0;
	reg [2:0] r_2339_0;
	reg [2:0] r_2340_0;
	reg [2:0] r_2341_0;
	reg [2:0] r_2342_0;
	reg [2:0] r_2343_0;
	reg [2:0] r_2344_0;
	reg [2:0] r_2345_0;
	reg [2:0] r_2346_0;
	reg [2:0] r_2347_0;
	reg [2:0] r_2348_0;
	reg [2:0] r_2349_0;
	reg [2:0] r_2350_0;
	reg [2:0] r_2351_0;
	reg [2:0] r_2352_0;
	reg [2:0] r_2353_0;
	reg [2:0] r_2354_0;
	reg [2:0] r_2355_0;
	reg [2:0] r_2356_0;
	reg [2:0] r_2357_0;
	reg [2:0] r_2358_0;
	reg [2:0] r_2359_0;
	reg [2:0] r_2360_0;
	reg [2:0] r_2361_0;
	reg [2:0] r_2362_0;
	reg [2:0] r_2363_0;
	reg [2:0] r_2364_0;
	reg [2:0] r_2365_0;
	reg [2:0] r_2366_0;
	reg [2:0] r_2367_0;
	reg [2:0] r_2368_0;
	reg [2:0] r_2369_0;
	reg [2:0] r_2370_0;
	reg [2:0] r_2371_0;
	reg [2:0] r_2372_0;
	reg [2:0] r_2373_0;
	reg [2:0] r_2374_0;
	reg [2:0] r_2375_0;
	reg [2:0] r_2376_0;
	reg [2:0] r_2377_0;
	reg [2:0] r_2378_0;
	reg [2:0] r_2379_0;
	reg [2:0] r_2380_0;
	reg [2:0] r_2381_0;
	reg [2:0] r_2382_0;
	reg [2:0] r_2383_0;
	reg [2:0] r_2384_0;
	reg [2:0] r_2385_0;
	reg [2:0] r_2386_0;
	reg [2:0] r_2387_0;
	reg [2:0] r_2388_0;
	reg [2:0] r_2389_0;
	reg [2:0] r_2390_0;
	reg [2:0] r_2391_0;
	reg [2:0] r_2392_0;
	reg [2:0] r_2393_0;
	reg [2:0] r_2394_0;
	reg [2:0] r_2395_0;
	reg [2:0] r_2396_0;
	reg [2:0] r_2397_0;
	reg [2:0] r_2398_0;
	reg [2:0] r_2399_0;
	reg [2:0] r_2400_0;
	reg [2:0] r_2401_0;
	reg [2:0] r_2402_0;
	reg [2:0] r_2403_0;
	reg [2:0] r_2404_0;
	reg [2:0] r_2405_0;
	reg [2:0] r_2406_0;
	reg [2:0] r_2407_0;
	reg [2:0] r_2408_0;
	reg [2:0] r_2409_0;
	reg [2:0] r_2410_0;
	reg [2:0] r_2411_0;
	reg [2:0] r_2412_0;
	reg [2:0] r_2413_0;
	reg [2:0] r_2414_0;
	reg [2:0] r_2415_0;
	reg [2:0] r_2416_0;
	reg [2:0] r_2417_0;
	reg [2:0] r_2418_0;
	reg [2:0] r_2419_0;
	reg [2:0] r_2420_0;
	reg [2:0] r_2421_0;
	reg [2:0] r_2422_0;
	reg [2:0] r_2423_0;
	reg [2:0] r_2424_0;
	reg [2:0] r_2425_0;
	reg [2:0] r_2426_0;
	reg [2:0] r_2427_0;
	reg [2:0] r_2428_0;
	reg [2:0] r_2429_0;
	reg [2:0] r_2430_0;
	reg [2:0] r_2431_0;
	reg [2:0] r_2432_0;
	reg [2:0] r_2433_0;
	reg [2:0] r_2434_0;
	reg [2:0] r_2435_0;
	reg [2:0] r_2436_0;
	reg [2:0] r_2437_0;
	reg [2:0] r_2438_0;
	reg [2:0] r_2439_0;
	reg [2:0] r_2440_0;
	reg [2:0] r_2441_0;
	reg [2:0] r_2442_0;
	reg [2:0] r_2443_0;
	reg [2:0] r_2444_0;
	reg [2:0] r_2445_0;
	reg [2:0] r_2446_0;
	reg [2:0] r_2447_0;
	reg [2:0] r_2448_0;
	reg [2:0] r_2449_0;
	reg [2:0] r_2450_0;
	reg [2:0] r_2451_0;
	reg [2:0] r_2452_0;
	reg [2:0] r_2453_0;
	reg [2:0] r_2454_0;
	reg [2:0] r_2455_0;
	reg [2:0] r_2456_0;
	reg [2:0] r_2457_0;
	reg [2:0] r_2458_0;
	reg [2:0] r_2459_0;
	reg [2:0] r_2460_0;
	reg [2:0] r_2461_0;
	reg [2:0] r_2462_0;
	reg [2:0] r_2463_0;
	reg [2:0] r_2464_0;
	reg [2:0] r_2465_0;
	reg [2:0] r_2466_0;
	reg [2:0] r_2467_0;
	reg [2:0] r_2468_0;
	reg [2:0] r_2469_0;
	reg [2:0] r_2470_0;
	reg [2:0] r_2471_0;
	reg [2:0] r_2472_0;
	reg [2:0] r_2473_0;
	reg [2:0] r_2474_0;
	reg [2:0] r_2475_0;
	reg [2:0] r_2476_0;
	reg [2:0] r_2477_0;
	reg [2:0] r_2478_0;
	reg [2:0] r_2479_0;
	reg [2:0] r_2480_0;
	reg [2:0] r_2481_0;
	reg [2:0] r_2482_0;
	reg [2:0] r_2483_0;
	reg [2:0] r_2484_0;
	reg [2:0] r_2485_0;
	reg [2:0] r_2486_0;
	reg [2:0] r_2487_0;
	reg [2:0] r_2488_0;
	reg [2:0] r_2489_0;
	reg [2:0] r_2490_0;
	reg [2:0] r_2491_0;
	reg [2:0] r_2492_0;
	reg [2:0] r_2493_0;
	reg [2:0] r_2494_0;
	reg [2:0] r_2495_0;
	reg [2:0] r_2496_0;
	reg [2:0] r_2497_0;
	reg [2:0] r_2498_0;
	reg [2:0] r_2499_0;
	reg [2:0] r_2500_0;
	reg [2:0] r_2501_0;
	reg [2:0] r_2502_0;
	reg [2:0] r_2503_0;
	reg [2:0] r_2504_0;
	reg [2:0] r_2505_0;
	reg [2:0] r_2506_0;
	reg [2:0] r_2507_0;
	reg [2:0] r_2508_0;
	reg [2:0] r_2509_0;
	reg [2:0] r_2510_0;
	reg [2:0] r_2511_0;
	reg [2:0] r_2512_0;
	reg [2:0] r_2513_0;
	reg [2:0] r_2514_0;
	reg [2:0] r_2515_0;
	reg [2:0] r_2516_0;
	reg [2:0] r_2517_0;
	reg [2:0] r_2518_0;
	reg [2:0] r_2519_0;
	reg [2:0] r_2520_0;
	reg [2:0] r_2521_0;
	reg [2:0] r_2522_0;
	reg [2:0] r_2523_0;
	reg [2:0] r_2524_0;
	reg [2:0] r_2525_0;
	reg [2:0] r_2526_0;
	reg [2:0] r_2527_0;
	reg [2:0] r_2528_0;
	reg [2:0] r_2529_0;
	reg [2:0] r_2530_0;
	reg [2:0] r_2531_0;
	reg [2:0] r_2532_0;
	reg [2:0] r_2533_0;
	reg [2:0] r_2534_0;
	reg [2:0] r_2535_0;
	reg [2:0] r_2536_0;
	reg [2:0] r_2537_0;
	reg [2:0] r_2538_0;
	reg [2:0] r_2539_0;
	reg [2:0] r_2540_0;
	reg [2:0] r_2541_0;
	reg [2:0] r_2542_0;
	reg [2:0] r_2543_0;
	reg [2:0] r_2544_0;
	reg [2:0] r_2545_0;
	reg [2:0] r_2546_0;
	reg [2:0] r_2547_0;
	reg [2:0] r_2548_0;
	reg [2:0] r_2549_0;
	reg [2:0] r_2550_0;
	reg [2:0] r_2551_0;
	reg [2:0] r_2552_0;
	reg [2:0] r_2553_0;
	reg [2:0] r_2554_0;
	reg [2:0] r_2555_0;
	reg [2:0] r_2556_0;
	reg [2:0] r_2557_0;
	reg [2:0] r_2558_0;
	reg [2:0] r_2559_0;
	reg [2:0] r_2560_0;
	reg [2:0] r_2561_0;
	reg [2:0] r_2562_0;
	reg [2:0] r_2563_0;
	reg [2:0] r_2564_0;
	reg [2:0] r_2565_0;
	reg [2:0] r_2566_0;
	reg [2:0] r_2567_0;
	reg [2:0] r_2568_0;
	reg [2:0] r_2569_0;
	reg [2:0] r_2570_0;
	reg [2:0] r_2571_0;
	reg [2:0] r_2572_0;
	reg [2:0] r_2573_0;
	reg [2:0] r_2574_0;
	reg [2:0] r_2575_0;
	reg [2:0] r_2576_0;
	reg [2:0] r_2577_0;
	reg [2:0] r_2578_0;
	reg [2:0] r_2579_0;
	reg [2:0] r_2580_0;
	reg [2:0] r_2581_0;
	reg [2:0] r_2582_0;
	reg [2:0] r_2583_0;
	reg [2:0] r_2584_0;
	reg [2:0] r_2585_0;
	reg [2:0] r_2586_0;
	reg [2:0] r_2587_0;
	reg [2:0] r_2588_0;
	reg [2:0] r_2589_0;
	reg [2:0] r_2590_0;
	reg [2:0] r_2591_0;
	reg [2:0] r_2592_0;
	reg [2:0] r_2593_0;
	reg [2:0] r_2594_0;
	reg [2:0] r_2595_0;
	reg [2:0] r_2596_0;
	reg [2:0] r_2597_0;
	reg [2:0] r_2598_0;
	reg [2:0] r_2599_0;
	reg [2:0] r_2600_0;
	reg [2:0] r_2601_0;
	reg [2:0] r_2602_0;
	reg [2:0] r_2603_0;
	reg [2:0] r_2604_0;
	reg [2:0] r_2605_0;
	reg [2:0] r_2606_0;
	reg [2:0] r_2607_0;
	reg [2:0] r_2608_0;
	reg [2:0] r_2609_0;
	reg [2:0] r_2610_0;
	reg [2:0] r_2611_0;
	reg [2:0] r_2612_0;
	reg [2:0] r_2613_0;
	reg [2:0] r_2614_0;
	reg [2:0] r_2615_0;
	reg [2:0] r_2616_0;
	reg [2:0] r_2617_0;
	reg [2:0] r_2618_0;
	reg [2:0] r_2619_0;
	reg [2:0] r_2620_0;
	reg [2:0] r_2621_0;
	reg [2:0] r_2622_0;
	reg [2:0] r_2623_0;
	reg [2:0] r_2624_0;
	reg [2:0] r_2625_0;
	reg [2:0] r_2626_0;
	reg [2:0] r_2627_0;
	reg [2:0] r_2628_0;
	reg [2:0] r_2629_0;
	reg [2:0] r_2630_0;
	reg [2:0] r_2631_0;
	reg [2:0] r_2632_0;
	reg [2:0] r_2633_0;
	reg [2:0] r_2634_0;
	reg [2:0] r_2635_0;
	reg [2:0] r_2636_0;
	reg [2:0] r_2637_0;
	reg [2:0] r_2638_0;
	reg [2:0] r_2639_0;
	reg [2:0] r_2640_0;
	reg [2:0] r_2641_0;
	reg [2:0] r_2642_0;
	reg [2:0] r_2643_0;
	reg [2:0] r_2644_0;
	reg [2:0] r_2645_0;
	reg [2:0] r_2646_0;
	reg [2:0] r_2647_0;
	reg [2:0] r_2648_0;
	reg [2:0] r_2649_0;
	reg [2:0] r_2650_0;
	reg [2:0] r_2651_0;
	reg [2:0] r_2652_0;
	reg [2:0] r_2653_0;
	reg [2:0] r_2654_0;
	reg [2:0] r_2655_0;
	reg [2:0] r_2656_0;
	reg [2:0] r_2657_0;
	reg [2:0] r_2658_0;
	reg [2:0] r_2659_0;
	reg [2:0] r_2660_0;
	reg [2:0] r_2661_0;
	reg [2:0] r_2662_0;
	reg [2:0] r_2663_0;
	reg [2:0] r_2664_0;
	reg [2:0] r_2665_0;
	reg [2:0] r_2666_0;
	reg [2:0] r_2667_0;
	reg [2:0] r_2668_0;
	reg [2:0] r_2669_0;
	reg [2:0] r_2670_0;
	reg [2:0] r_2671_0;
	reg [2:0] r_2672_0;
	reg [2:0] r_2673_0;
	reg [2:0] r_2674_0;
	reg [2:0] r_2675_0;
	reg [2:0] r_2676_0;
	reg [2:0] r_2677_0;
	reg [2:0] r_2678_0;
	reg [2:0] r_2679_0;
	reg [2:0] r_2680_0;
	reg [2:0] r_2681_0;
	reg [2:0] r_2682_0;
	reg [2:0] r_2683_0;
	reg [2:0] r_2684_0;
	reg [2:0] r_2685_0;
	reg [2:0] r_2686_0;
	reg [2:0] r_2687_0;
	reg [2:0] r_2688_0;
	reg [2:0] r_2689_0;
	reg [2:0] r_2690_0;
	reg [2:0] r_2691_0;
	reg [2:0] r_2692_0;
	reg [2:0] r_2693_0;
	reg [2:0] r_2694_0;
	reg [2:0] r_2695_0;
	reg [2:0] r_2696_0;
	reg [2:0] r_2697_0;
	reg [2:0] r_2698_0;
	reg [2:0] r_2699_0;
	reg [2:0] r_2700_0;
	reg [2:0] r_2701_0;
	reg [2:0] r_2702_0;
	reg [2:0] r_2703_0;
	reg [2:0] r_2704_0;
	reg [2:0] r_2705_0;
	reg [2:0] r_2706_0;
	reg [2:0] r_2707_0;
	reg [2:0] r_2708_0;
	reg [2:0] r_2709_0;
	reg [2:0] r_2710_0;
	reg [2:0] r_2711_0;
	reg [2:0] r_2712_0;
	reg [2:0] r_2713_0;
	reg [2:0] r_2714_0;
	reg [2:0] r_2715_0;
	reg [2:0] r_2716_0;
	reg [2:0] r_2717_0;
	reg [2:0] r_2718_0;
	reg [2:0] r_2719_0;
	reg [2:0] r_2720_0;
	reg [2:0] r_2721_0;
	reg [2:0] r_2722_0;
	reg [2:0] r_2723_0;
	reg [2:0] r_2724_0;
	reg [2:0] r_2725_0;
	reg [2:0] r_2726_0;
	reg [2:0] r_2727_0;
	reg [2:0] r_2728_0;
	reg [2:0] r_2729_0;
	reg [2:0] r_2730_0;
	reg [2:0] r_2731_0;
	reg [2:0] r_2732_0;
	reg [2:0] r_2733_0;
	reg [2:0] r_2734_0;
	reg [2:0] r_2735_0;
	reg [2:0] r_2736_0;
	reg [2:0] r_2737_0;
	reg [2:0] r_2738_0;
	reg [2:0] r_2739_0;
	reg [2:0] r_2740_0;
	reg [2:0] r_2741_0;
	reg [2:0] r_2742_0;
	reg [2:0] r_2743_0;
	reg [2:0] r_2744_0;
	reg [2:0] r_2745_0;
	reg [2:0] r_2746_0;
	reg [2:0] r_2747_0;
	reg [2:0] r_2748_0;
	reg [2:0] r_2749_0;
	reg [2:0] r_2750_0;
	reg [2:0] r_2751_0;
	reg [2:0] r_2752_0;
	reg [2:0] r_2753_0;
	reg [2:0] r_2754_0;
	reg [2:0] r_2755_0;
	reg [2:0] r_2756_0;
	reg [2:0] r_2757_0;
	reg [2:0] r_2758_0;
	reg [2:0] r_2759_0;
	reg [2:0] r_2760_0;
	reg [2:0] r_2761_0;
	reg [2:0] r_2762_0;
	reg [2:0] r_2763_0;
	reg [2:0] r_2764_0;
	reg [2:0] r_2765_0;
	reg [2:0] r_2766_0;
	reg [2:0] r_2767_0;
	reg [2:0] r_2768_0;
	reg [2:0] r_2769_0;
	reg [2:0] r_2770_0;
	reg [2:0] r_2771_0;
	reg [2:0] r_2772_0;
	reg [2:0] r_2773_0;
	reg [2:0] r_2774_0;
	reg [2:0] r_2775_0;
	reg [2:0] r_2776_0;
	reg [2:0] r_2777_0;
	reg [2:0] r_2778_0;
	reg [2:0] r_2779_0;
	reg [2:0] r_2780_0;
	reg [2:0] r_2781_0;
	reg [2:0] r_2782_0;
	reg [2:0] r_2783_0;
	reg [2:0] r_2784_0;
	reg [2:0] r_2785_0;
	reg [2:0] r_2786_0;
	reg [2:0] r_2787_0;
	reg [2:0] r_2788_0;
	reg [2:0] r_2789_0;
	reg [2:0] r_2790_0;
	reg [2:0] r_2791_0;
	reg [2:0] r_2792_0;
	reg [2:0] r_2793_0;
	reg [2:0] r_2794_0;
	reg [2:0] r_2795_0;
	reg [2:0] r_2796_0;
	reg [2:0] r_2797_0;
	reg [2:0] r_2798_0;
	reg [2:0] r_2799_0;
	reg [2:0] r_2800_0;
	reg [2:0] r_2801_0;
	reg [2:0] r_2802_0;
	reg [2:0] r_2803_0;
	reg [2:0] r_2804_0;
	reg [2:0] r_2805_0;
	reg [2:0] r_2806_0;
	reg [2:0] r_2807_0;
	reg [2:0] r_2808_0;
	reg [2:0] r_2809_0;
	reg [2:0] r_2810_0;
	reg [2:0] r_2811_0;
	reg [2:0] r_2812_0;
	reg [2:0] r_2813_0;
	reg [2:0] r_2814_0;
	reg [2:0] r_2815_0;
	reg [2:0] r_2816_0;
	reg [2:0] r_2817_0;
	reg [2:0] r_2818_0;
	reg [2:0] r_2819_0;
	reg [2:0] r_2820_0;
	reg [2:0] r_2821_0;
	reg [2:0] r_2822_0;
	reg [2:0] r_2823_0;
	reg [2:0] r_2824_0;
	reg [2:0] r_2825_0;
	reg [2:0] r_2826_0;
	reg [2:0] r_2827_0;
	reg [2:0] r_2828_0;
	reg [2:0] r_2829_0;
	reg [2:0] r_2830_0;
	reg [2:0] r_2831_0;
	reg [2:0] r_2832_0;
	reg [2:0] r_2833_0;
	reg [2:0] r_2834_0;
	reg [2:0] r_2835_0;
	reg [2:0] r_2836_0;
	reg [2:0] r_2837_0;
	reg [2:0] r_2838_0;
	reg [2:0] r_2839_0;
	reg [2:0] r_2840_0;
	reg [2:0] r_2841_0;
	reg [2:0] r_2842_0;
	reg [2:0] r_2843_0;
	reg [2:0] r_2844_0;
	reg [2:0] r_2845_0;
	reg [2:0] r_2846_0;
	reg [2:0] r_2847_0;
	reg [2:0] r_2848_0;
	reg [2:0] r_2849_0;
	reg [2:0] r_2850_0;
	reg [2:0] r_2851_0;
	reg [2:0] r_2852_0;
	reg [2:0] r_2853_0;
	reg [2:0] r_2854_0;
	reg [2:0] r_2855_0;
	reg [2:0] r_2856_0;
	reg [2:0] r_2857_0;
	reg [2:0] r_2858_0;
	reg [2:0] r_2859_0;
	reg [2:0] r_2860_0;
	reg [2:0] r_2861_0;
	reg [2:0] r_2862_0;
	reg [2:0] r_2863_0;
	reg [2:0] r_2864_0;
	reg [2:0] r_2865_0;
	reg [2:0] r_2866_0;
	reg [2:0] r_2867_0;
	reg [2:0] r_2868_0;
	reg [2:0] r_2869_0;
	reg [2:0] r_2870_0;
	reg [2:0] r_2871_0;
	reg [2:0] r_2872_0;
	reg [2:0] r_2873_0;
	reg [2:0] r_2874_0;
	reg [2:0] r_2875_0;
	reg [2:0] r_2876_0;
	reg [2:0] r_2877_0;
	reg [2:0] r_2878_0;
	reg [2:0] r_2879_0;
	reg [2:0] r_2880_0;
	reg [2:0] r_2881_0;
	reg [2:0] r_2882_0;
	reg [2:0] r_2883_0;
	reg [2:0] r_2884_0;
	reg [2:0] r_2885_0;
	reg [2:0] r_2886_0;
	reg [2:0] r_2887_0;
	reg [2:0] r_2888_0;
	reg [2:0] r_2889_0;
	reg [2:0] r_2890_0;
	reg [2:0] r_2891_0;
	reg [2:0] r_2892_0;
	reg [2:0] r_2893_0;
	reg [2:0] r_2894_0;
	reg [2:0] r_2895_0;
	reg [2:0] r_2896_0;
	reg [2:0] r_2897_0;
	reg [2:0] r_2898_0;
	reg [2:0] r_2899_0;
	reg [2:0] r_2900_0;
	reg [2:0] r_2901_0;
	reg [2:0] r_2902_0;
	reg [2:0] r_2903_0;
	reg [2:0] r_2904_0;
	reg [2:0] r_2905_0;
	reg [2:0] r_2906_0;
	reg [2:0] r_2907_0;
	reg [2:0] r_2908_0;
	reg [2:0] r_2909_0;
	reg [2:0] r_2910_0;
	reg [2:0] r_2911_0;
	reg [2:0] r_2912_0;
	reg [2:0] r_2913_0;
	reg [2:0] r_2914_0;
	reg [2:0] r_2915_0;
	reg [2:0] r_2916_0;
	reg [2:0] r_2917_0;
	reg [2:0] r_2918_0;
	reg [2:0] r_2919_0;
	reg [2:0] r_2920_0;
	reg [2:0] r_2921_0;
	reg [2:0] r_2922_0;
	reg [2:0] r_2923_0;
	reg [2:0] r_2924_0;
	reg [2:0] r_2925_0;
	reg [2:0] r_2926_0;
	reg [2:0] r_2927_0;
	reg [2:0] r_2928_0;
	reg [2:0] r_2929_0;
	reg [2:0] r_2930_0;
	reg [2:0] r_2931_0;
	reg [2:0] r_2932_0;
	reg [2:0] r_2933_0;
	reg [2:0] r_2934_0;
	reg [2:0] r_2935_0;
	reg [2:0] r_2936_0;
	reg [2:0] r_2937_0;
	reg [2:0] r_2938_0;
	reg [2:0] r_2939_0;
	reg [2:0] r_2940_0;
	reg [2:0] r_2941_0;
	reg [2:0] r_2942_0;
	reg [2:0] r_2943_0;
	reg [2:0] r_2944_0;
	reg [2:0] r_2945_0;
	reg [2:0] r_2946_0;
	reg [2:0] r_2947_0;
	reg [2:0] r_2948_0;
	reg [2:0] r_2949_0;
	reg [2:0] r_2950_0;
	reg [2:0] r_2951_0;
	reg [2:0] r_2952_0;
	reg [2:0] r_2953_0;
	reg [2:0] r_2954_0;
	reg [2:0] r_2955_0;
	reg [2:0] r_2956_0;
	reg [2:0] r_2957_0;
	reg [2:0] r_2958_0;
	reg [2:0] r_2959_0;
	reg [2:0] r_2960_0;
	reg [2:0] r_2961_0;
	reg [2:0] r_2962_0;
	reg [2:0] r_2963_0;
	reg [2:0] r_2964_0;
	reg [2:0] r_2965_0;
	reg [2:0] r_2966_0;
	reg [2:0] r_2967_0;
	reg [2:0] r_2968_0;
	reg [2:0] r_2969_0;
	reg [2:0] r_2970_0;
	reg [2:0] r_2971_0;
	reg [2:0] r_2972_0;
	reg [2:0] r_2973_0;
	reg [2:0] r_2974_0;
	reg [2:0] r_2975_0;
	reg [2:0] r_2976_0;
	reg [2:0] r_2977_0;
	reg [2:0] r_2978_0;
	reg [2:0] r_2979_0;
	reg [2:0] r_2980_0;
	reg [2:0] r_2981_0;
	reg [2:0] r_2982_0;
	reg [2:0] r_2983_0;
	reg [2:0] r_2984_0;
	reg [2:0] r_2985_0;
	reg [2:0] r_2986_0;
	reg [2:0] r_2987_0;
	reg [2:0] r_2988_0;
	reg [2:0] r_2989_0;
	reg [2:0] r_2990_0;
	reg [2:0] r_2991_0;
	reg [2:0] r_2992_0;
	reg [2:0] r_2993_0;
	reg [2:0] r_2994_0;
	reg [2:0] r_2995_0;
	reg [2:0] r_2996_0;
	reg [2:0] r_2997_0;
	reg [2:0] r_2998_0;
	reg [2:0] r_2999_0;
	reg [2:0] r_3000_0;
	reg [2:0] r_3001_0;
	reg [2:0] r_3002_0;
	reg [2:0] r_3003_0;
	reg [2:0] r_3004_0;
	reg [2:0] r_3005_0;
	reg [2:0] r_3006_0;
	reg [2:0] r_3007_0;
	reg [2:0] r_3008_0;
	reg [2:0] r_3009_0;
	reg [2:0] r_3010_0;
	reg [2:0] r_3011_0;
	reg [2:0] r_3012_0;
	reg [2:0] r_3013_0;
	reg [2:0] r_3014_0;
	reg [2:0] r_3015_0;
	reg [2:0] r_3016_0;
	reg [2:0] r_3017_0;
	reg [2:0] r_3018_0;
	reg [2:0] r_3019_0;
	reg [2:0] r_3020_0;
	reg [2:0] r_3021_0;
	reg [2:0] r_3022_0;
	reg [2:0] r_3023_0;
	reg [2:0] r_3024_0;
	reg [2:0] r_3025_0;
	reg [2:0] r_3026_0;
	reg [2:0] r_3027_0;
	reg [2:0] r_3028_0;
	reg [2:0] r_3029_0;
	reg [2:0] r_3030_0;
	reg [2:0] r_3031_0;
	reg [2:0] r_3032_0;
	reg [2:0] r_3033_0;
	reg [2:0] r_3034_0;
	reg [2:0] r_3035_0;
	reg [2:0] r_3036_0;
	reg [2:0] r_3037_0;
	reg [2:0] r_3038_0;
	reg [2:0] r_3039_0;
	reg [2:0] r_3040_0;
	reg [2:0] r_3041_0;
	reg [2:0] r_3042_0;
	reg [2:0] r_3043_0;
	reg [2:0] r_3044_0;
	reg [2:0] r_3045_0;
	reg [2:0] r_3046_0;
	reg [2:0] r_3047_0;
	reg [2:0] r_3048_0;
	reg [2:0] r_3049_0;
	reg [2:0] r_3050_0;
	reg [2:0] r_3051_0;
	reg [2:0] r_3052_0;
	reg [2:0] r_3053_0;
	reg [2:0] r_3054_0;
	reg [2:0] r_3055_0;
	reg [2:0] r_3056_0;
	reg [2:0] r_3057_0;
	reg [2:0] r_3058_0;
	reg [2:0] r_3059_0;
	reg [2:0] r_3060_0;
	reg [2:0] r_3061_0;
	reg [2:0] r_3062_0;
	reg [2:0] r_3063_0;
	reg [2:0] r_3064_0;
	reg [2:0] r_3065_0;
	reg [2:0] r_3066_0;
	reg [2:0] r_3067_0;
	reg [2:0] r_3068_0;
	reg [2:0] r_3069_0;
	reg [2:0] r_3070_0;
	reg [2:0] r_3071_0;
	reg r_3072_0;
	reg r_3073_0;
	reg r_3074_0;
	reg r_3075_0;
	reg r_3076_0;
	reg r_3077_0;
	reg r_3078_0;
	reg r_3079_0;
	reg r_3080_0;
	reg r_3081_0;
	reg r_3082_0;
	reg r_3083_0;
	reg r_3084_0;
	reg r_3085_0;
	reg r_3086_0;
	reg r_3087_0;
	reg r_3088_0;
	reg r_3089_0;
	reg r_3090_0;
	reg r_3091_0;
	reg r_3092_0;
	reg r_3093_0;
	reg r_3094_0;
	reg r_3095_0;
	reg r_3096_0;
	reg r_3097_0;
	reg r_3098_0;
	reg r_3099_0;
	reg r_3100_0;
	reg r_3101_0;
	reg r_3102_0;
	reg r_3103_0;
	reg r_3104_0;
	reg r_3105_0;
	reg r_3106_0;
	reg r_3107_0;
	reg r_3108_0;
	reg r_3109_0;
	reg r_3110_0;
	reg r_3111_0;
	reg r_3112_0;
	reg r_3113_0;
	reg r_3114_0;
	reg r_3115_0;
	reg r_3116_0;
	reg r_3117_0;
	reg r_3118_0;
	reg r_3119_0;
	reg r_3120_0;
	reg r_3121_0;
	reg r_3122_0;
	reg r_3123_0;
	reg r_3124_0;
	reg r_3125_0;
	reg r_3126_0;
	reg r_3127_0;
	reg r_3128_0;
	reg r_3129_0;
	reg r_3130_0;
	reg r_3131_0;
	reg r_3132_0;
	reg r_3133_0;
	reg r_3134_0;
	reg r_3135_0;
	reg r_3136_0;
	reg r_3137_0;
	reg r_3138_0;
	reg r_3139_0;
	reg r_3140_0;
	reg r_3141_0;
	reg r_3142_0;
	reg r_3143_0;
	reg r_3144_0;
	reg r_3145_0;
	reg r_3146_0;
	reg r_3147_0;
	reg r_3148_0;
	reg r_3149_0;
	reg r_3150_0;
	reg r_3151_0;
	reg r_3152_0;
	reg r_3153_0;
	reg r_3154_0;
	reg r_3155_0;
	reg r_3156_0;
	reg r_3157_0;
	reg r_3158_0;
	reg r_3159_0;
	reg r_3160_0;
	reg r_3161_0;
	reg r_3162_0;
	reg r_3163_0;
	reg r_3164_0;
	reg r_3165_0;
	reg r_3166_0;
	reg r_3167_0;
	reg r_3168_0;
	reg r_3169_0;
	reg r_3170_0;
	reg r_3171_0;
	reg r_3172_0;
	reg r_3173_0;
	reg r_3174_0;
	reg r_3175_0;
	reg r_3176_0;
	reg r_3177_0;
	reg r_3178_0;
	reg r_3179_0;
	reg r_3180_0;
	reg r_3181_0;
	reg r_3182_0;
	reg r_3183_0;
	reg r_3184_0;
	reg r_3185_0;
	reg r_3186_0;
	reg r_3187_0;
	reg r_3188_0;
	reg r_3189_0;
	reg r_3190_0;
	reg r_3191_0;
	reg r_3192_0;
	reg r_3193_0;
	reg r_3194_0;
	reg r_3195_0;
	reg r_3196_0;
	reg r_3197_0;
	reg r_3198_0;
	reg r_3199_0;
	reg r_3200_0;
	reg r_3201_0;
	reg r_3202_0;
	reg r_3203_0;
	reg r_3204_0;
	reg r_3205_0;
	reg r_3206_0;
	reg r_3207_0;
	reg r_3208_0;
	reg r_3209_0;
	reg r_3210_0;
	reg r_3211_0;
	reg r_3212_0;
	reg r_3213_0;
	reg r_3214_0;
	reg r_3215_0;
	reg r_3216_0;
	reg r_3217_0;
	reg r_3218_0;
	reg r_3219_0;
	reg r_3220_0;
	reg r_3221_0;
	reg r_3222_0;
	reg r_3223_0;
	reg r_3224_0;
	reg r_3225_0;
	reg r_3226_0;
	reg r_3227_0;
	reg r_3228_0;
	reg r_3229_0;
	reg r_3230_0;
	reg r_3231_0;
	reg r_3232_0;
	reg r_3233_0;
	reg r_3234_0;
	reg r_3235_0;
	reg r_3236_0;
	reg r_3237_0;
	reg r_3238_0;
	reg r_3239_0;
	reg r_3240_0;
	reg r_3241_0;
	reg r_3242_0;
	reg r_3243_0;
	reg r_3244_0;
	reg r_3245_0;
	reg r_3246_0;
	reg r_3247_0;
	reg r_3248_0;
	reg r_3249_0;
	reg r_3250_0;
	reg r_3251_0;
	reg r_3252_0;
	reg r_3253_0;
	reg r_3254_0;
	reg r_3255_0;
	reg r_3256_0;
	reg r_3257_0;
	reg r_3258_0;
	reg r_3259_0;
	reg r_3260_0;
	reg r_3261_0;
	reg r_3262_0;
	reg r_3263_0;
	reg r_3264_0;
	reg r_3265_0;
	reg r_3266_0;
	reg r_3267_0;
	reg r_3268_0;
	reg r_3269_0;
	reg r_3270_0;
	reg r_3271_0;
	reg r_3272_0;
	reg r_3273_0;
	reg r_3274_0;
	reg r_3275_0;
	reg r_3276_0;
	reg r_3277_0;
	reg r_3278_0;
	reg r_3279_0;
	reg r_3280_0;
	reg r_3281_0;
	reg r_3282_0;
	reg r_3283_0;
	reg r_3284_0;
	reg r_3285_0;
	reg r_3286_0;
	reg r_3287_0;
	reg r_3288_0;
	reg r_3289_0;
	reg r_3290_0;
	reg r_3291_0;
	reg r_3292_0;
	reg r_3293_0;
	reg r_3294_0;
	reg r_3295_0;
	reg r_3296_0;
	reg r_3297_0;
	reg r_3298_0;
	reg r_3299_0;
	reg r_3300_0;
	reg r_3301_0;
	reg r_3302_0;
	reg r_3303_0;
	reg r_3304_0;
	reg r_3305_0;
	reg r_3306_0;
	reg r_3307_0;
	reg r_3308_0;
	reg r_3309_0;
	reg r_3310_0;
	reg r_3311_0;
	reg r_3312_0;
	reg r_3313_0;
	reg r_3314_0;
	reg r_3315_0;
	reg r_3316_0;
	reg r_3317_0;
	reg r_3318_0;
	reg r_3319_0;
	reg r_3320_0;
	reg r_3321_0;
	reg r_3322_0;
	reg r_3323_0;
	reg r_3324_0;
	reg r_3325_0;
	reg r_3326_0;
	reg r_3327_0;
	reg r_3328_0;
	reg r_3329_0;
	reg r_3330_0;
	reg r_3331_0;
	reg r_3332_0;
	reg r_3333_0;
	reg r_3334_0;
	reg r_3335_0;
	reg r_3336_0;
	reg r_3337_0;
	reg r_3338_0;
	reg r_3339_0;
	reg r_3340_0;
	reg r_3341_0;
	reg r_3342_0;
	reg r_3343_0;
	reg r_3344_0;
	reg r_3345_0;
	reg r_3346_0;
	reg r_3347_0;
	reg r_3348_0;
	reg r_3349_0;
	reg r_3350_0;
	reg r_3351_0;
	reg r_3352_0;
	reg r_3353_0;
	reg r_3354_0;
	reg r_3355_0;
	reg r_3356_0;
	reg r_3357_0;
	reg r_3358_0;
	reg r_3359_0;
	reg r_3360_0;
	reg r_3361_0;
	reg r_3362_0;
	reg r_3363_0;
	reg r_3364_0;
	reg r_3365_0;
	reg r_3366_0;
	reg r_3367_0;
	reg r_3368_0;
	reg r_3369_0;
	reg r_3370_0;
	reg r_3371_0;
	reg r_3372_0;
	reg r_3373_0;
	reg r_3374_0;
	reg r_3375_0;
	reg r_3376_0;
	reg r_3377_0;
	reg r_3378_0;
	reg r_3379_0;
	reg r_3380_0;
	reg r_3381_0;
	reg r_3382_0;
	reg r_3383_0;
	reg r_3384_0;
	reg r_3385_0;
	reg r_3386_0;
	reg r_3387_0;
	reg r_3388_0;
	reg r_3389_0;
	reg r_3390_0;
	reg r_3391_0;
	reg r_3392_0;
	reg r_3393_0;
	reg r_3394_0;
	reg r_3395_0;
	reg r_3396_0;
	reg r_3397_0;
	reg r_3398_0;
	reg r_3399_0;
	reg r_3400_0;
	reg r_3401_0;
	reg r_3402_0;
	reg r_3403_0;
	reg r_3404_0;
	reg r_3405_0;
	reg r_3406_0;
	reg r_3407_0;
	reg r_3408_0;
	reg r_3409_0;
	reg r_3410_0;
	reg r_3411_0;
	reg r_3412_0;
	reg r_3413_0;
	reg r_3414_0;
	reg r_3415_0;
	reg r_3416_0;
	reg r_3417_0;
	reg r_3418_0;
	reg r_3419_0;
	reg r_3420_0;
	reg r_3421_0;
	reg r_3422_0;
	reg r_3423_0;
	reg r_3424_0;
	reg r_3425_0;
	reg r_3426_0;
	reg r_3427_0;
	reg r_3428_0;
	reg r_3429_0;
	reg r_3430_0;
	reg r_3431_0;
	reg r_3432_0;
	reg r_3433_0;
	reg r_3434_0;
	reg r_3435_0;
	reg r_3436_0;
	reg r_3437_0;
	reg r_3438_0;
	reg r_3439_0;
	reg r_3440_0;
	reg r_3441_0;
	reg r_3442_0;
	reg r_3443_0;
	reg r_3444_0;
	reg r_3445_0;
	reg r_3446_0;
	reg r_3447_0;
	reg r_3448_0;
	reg r_3449_0;
	reg r_3450_0;
	reg r_3451_0;
	reg r_3452_0;
	reg r_3453_0;
	reg r_3454_0;
	reg r_3455_0;
	reg r_3456_0;
	reg r_3457_0;
	reg r_3458_0;
	reg r_3459_0;
	reg r_3460_0;
	reg r_3461_0;
	reg r_3462_0;
	reg r_3463_0;
	reg r_3464_0;
	reg r_3465_0;
	reg r_3466_0;
	reg r_3467_0;
	reg r_3468_0;
	reg r_3469_0;
	reg r_3470_0;
	reg r_3471_0;
	reg r_3472_0;
	reg r_3473_0;
	reg r_3474_0;
	reg r_3475_0;
	reg r_3476_0;
	reg r_3477_0;
	reg r_3478_0;
	reg r_3479_0;
	reg r_3480_0;
	reg r_3481_0;
	reg r_3482_0;
	reg r_3483_0;
	reg r_3484_0;
	reg r_3485_0;
	reg r_3486_0;
	reg r_3487_0;
	reg r_3488_0;
	reg r_3489_0;
	reg r_3490_0;
	reg r_3491_0;
	reg r_3492_0;
	reg r_3493_0;
	reg r_3494_0;
	reg r_3495_0;
	reg r_3496_0;
	reg r_3497_0;
	reg r_3498_0;
	reg r_3499_0;
	reg r_3500_0;
	reg r_3501_0;
	reg r_3502_0;
	reg r_3503_0;
	reg r_3504_0;
	reg r_3505_0;
	reg r_3506_0;
	reg r_3507_0;
	reg r_3508_0;
	reg r_3509_0;
	reg r_3510_0;
	reg r_3511_0;
	reg r_3512_0;
	reg r_3513_0;
	reg r_3514_0;
	reg r_3515_0;
	reg r_3516_0;
	reg r_3517_0;
	reg r_3518_0;
	reg r_3519_0;
	reg r_3520_0;
	reg r_3521_0;
	reg r_3522_0;
	reg r_3523_0;
	reg r_3524_0;
	reg r_3525_0;
	reg r_3526_0;
	reg r_3527_0;
	reg r_3528_0;
	reg r_3529_0;
	reg r_3530_0;
	reg r_3531_0;
	reg r_3532_0;
	reg r_3533_0;
	reg r_3534_0;
	reg r_3535_0;
	reg r_3536_0;
	reg r_3537_0;
	reg r_3538_0;
	reg r_3539_0;
	reg r_3540_0;
	reg r_3541_0;
	reg r_3542_0;
	reg r_3543_0;
	reg r_3544_0;
	reg r_3545_0;
	reg r_3546_0;
	reg r_3547_0;
	reg r_3548_0;
	reg r_3549_0;
	reg r_3550_0;
	reg r_3551_0;
	reg r_3552_0;
	reg r_3553_0;
	reg r_3554_0;
	reg r_3555_0;
	reg r_3556_0;
	reg r_3557_0;
	reg r_3558_0;
	reg r_3559_0;
	reg r_3560_0;
	reg r_3561_0;
	reg r_3562_0;
	reg r_3563_0;
	reg r_3564_0;
	reg r_3565_0;
	reg r_3566_0;
	reg r_3567_0;
	reg r_3568_0;
	reg r_3569_0;
	reg r_3570_0;
	reg r_3571_0;
	reg r_3572_0;
	reg r_3573_0;
	reg r_3574_0;
	reg r_3575_0;
	reg r_3576_0;
	reg r_3577_0;
	reg r_3578_0;
	reg r_3579_0;
	reg r_3580_0;
	reg r_3581_0;
	reg r_3582_0;
	reg r_3583_0;
	reg r_3584_0;
	reg r_3585_0;
	reg r_3586_0;
	reg r_3587_0;
	reg r_3588_0;
	reg r_3589_0;
	reg r_3590_0;
	reg r_3591_0;
	reg r_3592_0;
	reg r_3593_0;
	reg r_3594_0;
	reg r_3595_0;
	reg r_3596_0;
	reg r_3597_0;
	reg r_3598_0;
	reg r_3599_0;
	reg r_3600_0;
	reg r_3601_0;
	reg r_3602_0;
	reg r_3603_0;
	reg r_3604_0;
	reg r_3605_0;
	reg r_3606_0;
	reg r_3607_0;
	reg r_3608_0;
	reg r_3609_0;
	reg r_3610_0;
	reg r_3611_0;
	reg r_3612_0;
	reg r_3613_0;
	reg r_3614_0;
	reg r_3615_0;
	reg r_3616_0;
	reg r_3617_0;
	reg r_3618_0;
	reg r_3619_0;
	reg r_3620_0;
	reg r_3621_0;
	reg r_3622_0;
	reg r_3623_0;
	reg r_3624_0;
	reg r_3625_0;
	reg r_3626_0;
	reg r_3627_0;
	reg r_3628_0;
	reg r_3629_0;
	reg r_3630_0;
	reg r_3631_0;
	reg r_3632_0;
	reg r_3633_0;
	reg r_3634_0;
	reg r_3635_0;
	reg r_3636_0;
	reg r_3637_0;
	reg r_3638_0;
	reg r_3639_0;
	reg r_3640_0;
	reg r_3641_0;
	reg r_3642_0;
	reg r_3643_0;
	reg r_3644_0;
	reg r_3645_0;
	reg r_3646_0;
	reg r_3647_0;
	reg r_3648_0;
	reg r_3649_0;
	reg r_3650_0;
	reg r_3651_0;
	reg r_3652_0;
	reg r_3653_0;
	reg r_3654_0;
	reg r_3655_0;
	reg r_3656_0;
	reg r_3657_0;
	reg r_3658_0;
	reg r_3659_0;
	reg r_3660_0;
	reg r_3661_0;
	reg r_3662_0;
	reg r_3663_0;
	reg r_3664_0;
	reg r_3665_0;
	reg r_3666_0;
	reg r_3667_0;
	reg r_3668_0;
	reg r_3669_0;
	reg r_3670_0;
	reg r_3671_0;
	reg r_3672_0;
	reg r_3673_0;
	reg r_3674_0;
	reg r_3675_0;
	reg r_3676_0;
	reg r_3677_0;
	reg r_3678_0;
	reg r_3679_0;
	reg r_3680_0;
	reg r_3681_0;
	reg r_3682_0;
	reg r_3683_0;
	reg r_3684_0;
	reg r_3685_0;
	reg r_3686_0;
	reg r_3687_0;
	reg r_3688_0;
	reg r_3689_0;
	reg r_3690_0;
	reg r_3691_0;
	reg r_3692_0;
	reg r_3693_0;
	reg r_3694_0;
	reg r_3695_0;
	reg r_3696_0;
	reg r_3697_0;
	reg r_3698_0;
	reg r_3699_0;
	reg r_3700_0;
	reg r_3701_0;
	reg r_3702_0;
	reg r_3703_0;
	reg r_3704_0;
	reg r_3705_0;
	reg r_3706_0;
	reg r_3707_0;
	reg r_3708_0;
	reg r_3709_0;
	reg r_3710_0;
	reg r_3711_0;
	reg r_3712_0;
	reg r_3713_0;
	reg r_3714_0;
	reg r_3715_0;
	reg r_3716_0;
	reg r_3717_0;
	reg r_3718_0;
	reg r_3719_0;
	reg r_3720_0;
	reg r_3721_0;
	reg r_3722_0;
	reg r_3723_0;
	reg r_3724_0;
	reg r_3725_0;
	reg r_3726_0;
	reg r_3727_0;
	reg r_3728_0;
	reg r_3729_0;
	reg r_3730_0;
	reg r_3731_0;
	reg r_3732_0;
	reg r_3733_0;
	reg r_3734_0;
	reg r_3735_0;
	reg r_3736_0;
	reg r_3737_0;
	reg r_3738_0;
	reg r_3739_0;
	reg r_3740_0;
	reg r_3741_0;
	reg r_3742_0;
	reg r_3743_0;
	reg r_3744_0;
	reg r_3745_0;
	reg r_3746_0;
	reg r_3747_0;
	reg r_3748_0;
	reg r_3749_0;
	reg r_3750_0;
	reg r_3751_0;
	reg r_3752_0;
	reg r_3753_0;
	reg r_3754_0;
	reg r_3755_0;
	reg r_3756_0;
	reg r_3757_0;
	reg r_3758_0;
	reg r_3759_0;
	reg r_3760_0;
	reg r_3761_0;
	reg r_3762_0;
	reg r_3763_0;
	reg r_3764_0;
	reg r_3765_0;
	reg r_3766_0;
	reg r_3767_0;
	reg r_3768_0;
	reg r_3769_0;
	reg r_3770_0;
	reg r_3771_0;
	reg r_3772_0;
	reg r_3773_0;
	reg r_3774_0;
	reg r_3775_0;
	reg r_3776_0;
	reg r_3777_0;
	reg r_3778_0;
	reg r_3779_0;
	reg r_3780_0;
	reg r_3781_0;
	reg r_3782_0;
	reg r_3783_0;
	reg r_3784_0;
	reg r_3785_0;
	reg r_3786_0;
	reg r_3787_0;
	reg r_3788_0;
	reg r_3789_0;
	reg r_3790_0;
	reg r_3791_0;
	reg r_3792_0;
	reg r_3793_0;
	reg r_3794_0;
	reg r_3795_0;
	reg r_3796_0;
	reg r_3797_0;
	reg r_3798_0;
	reg r_3799_0;
	reg r_3800_0;
	reg r_3801_0;
	reg r_3802_0;
	reg r_3803_0;
	reg r_3804_0;
	reg r_3805_0;
	reg r_3806_0;
	reg r_3807_0;
	reg r_3808_0;
	reg r_3809_0;
	reg r_3810_0;
	reg r_3811_0;
	reg r_3812_0;
	reg r_3813_0;
	reg r_3814_0;
	reg r_3815_0;
	reg r_3816_0;
	reg r_3817_0;
	reg r_3818_0;
	reg r_3819_0;
	reg r_3820_0;
	reg r_3821_0;
	reg r_3822_0;
	reg r_3823_0;
	reg r_3824_0;
	reg r_3825_0;
	reg r_3826_0;
	reg r_3827_0;
	reg r_3828_0;
	reg r_3829_0;
	reg r_3830_0;
	reg r_3831_0;
	reg r_3832_0;
	reg r_3833_0;
	reg r_3834_0;
	reg r_3835_0;
	reg r_3836_0;
	reg r_3837_0;
	reg r_3838_0;
	reg r_3839_0;
	reg r_3840_0;
	reg r_3841_0;
	reg r_3842_0;
	reg r_3843_0;
	reg r_3844_0;
	reg r_3845_0;
	reg r_3846_0;
	reg r_3847_0;
	reg r_3848_0;
	reg r_3849_0;
	reg r_3850_0;
	reg r_3851_0;
	reg r_3852_0;
	reg r_3853_0;
	reg r_3854_0;
	reg r_3855_0;
	reg r_3856_0;
	reg r_3857_0;
	reg r_3858_0;
	reg r_3859_0;
	reg r_3860_0;
	reg r_3861_0;
	reg r_3862_0;
	reg r_3863_0;
	reg r_3864_0;
	reg r_3865_0;
	reg r_3866_0;
	reg r_3867_0;
	reg r_3868_0;
	reg r_3869_0;
	reg r_3870_0;
	reg r_3871_0;
	reg r_3872_0;
	reg r_3873_0;
	reg r_3874_0;
	reg r_3875_0;
	reg r_3876_0;
	reg r_3877_0;
	reg r_3878_0;
	reg r_3879_0;
	reg r_3880_0;
	reg r_3881_0;
	reg r_3882_0;
	reg r_3883_0;
	reg r_3884_0;
	reg r_3885_0;
	reg r_3886_0;
	reg r_3887_0;
	reg r_3888_0;
	reg r_3889_0;
	reg r_3890_0;
	reg r_3891_0;
	reg r_3892_0;
	reg r_3893_0;
	reg r_3894_0;
	reg r_3895_0;
	reg r_3896_0;
	reg r_3897_0;
	reg r_3898_0;
	reg r_3899_0;
	reg r_3900_0;
	reg r_3901_0;
	reg r_3902_0;
	reg r_3903_0;
	reg r_3904_0;
	reg r_3905_0;
	reg r_3906_0;
	reg r_3907_0;
	reg r_3908_0;
	reg r_3909_0;
	reg r_3910_0;
	reg r_3911_0;
	reg r_3912_0;
	reg r_3913_0;
	reg r_3914_0;
	reg r_3915_0;
	reg r_3916_0;
	reg r_3917_0;
	reg r_3918_0;
	reg r_3919_0;
	reg r_3920_0;
	reg r_3921_0;
	reg r_3922_0;
	reg r_3923_0;
	reg r_3924_0;
	reg r_3925_0;
	reg r_3926_0;
	reg r_3927_0;
	reg r_3928_0;
	reg r_3929_0;
	reg r_3930_0;
	reg r_3931_0;
	reg r_3932_0;
	reg r_3933_0;
	reg r_3934_0;
	reg r_3935_0;
	reg r_3936_0;
	reg r_3937_0;
	reg r_3938_0;
	reg r_3939_0;
	reg r_3940_0;
	reg r_3941_0;
	reg r_3942_0;
	reg r_3943_0;
	reg r_3944_0;
	reg r_3945_0;
	reg r_3946_0;
	reg r_3947_0;
	reg r_3948_0;
	reg r_3949_0;
	reg r_3950_0;
	reg r_3951_0;
	reg r_3952_0;
	reg r_3953_0;
	reg r_3954_0;
	reg r_3955_0;
	reg r_3956_0;
	reg r_3957_0;
	reg r_3958_0;
	reg r_3959_0;
	reg r_3960_0;
	reg r_3961_0;
	reg r_3962_0;
	reg r_3963_0;
	reg r_3964_0;
	reg r_3965_0;
	reg r_3966_0;
	reg r_3967_0;
	reg r_3968_0;
	reg r_3969_0;
	reg r_3970_0;
	reg r_3971_0;
	reg r_3972_0;
	reg r_3973_0;
	reg r_3974_0;
	reg r_3975_0;
	reg r_3976_0;
	reg r_3977_0;
	reg r_3978_0;
	reg r_3979_0;
	reg r_3980_0;
	reg r_3981_0;
	reg r_3982_0;
	reg r_3983_0;
	reg r_3984_0;
	reg r_3985_0;
	reg r_3986_0;
	reg r_3987_0;
	reg r_3988_0;
	reg r_3989_0;
	reg r_3990_0;
	reg r_3991_0;
	reg r_3992_0;
	reg r_3993_0;
	reg r_3994_0;
	reg r_3995_0;
	reg r_3996_0;
	reg r_3997_0;
	reg r_3998_0;
	reg r_3999_0;
	reg r_4000_0;
	reg r_4001_0;
	reg r_4002_0;
	reg r_4003_0;
	reg r_4004_0;
	reg r_4005_0;
	reg r_4006_0;
	reg r_4007_0;
	reg r_4008_0;
	reg r_4009_0;
	reg r_4010_0;
	reg r_4011_0;
	reg r_4012_0;
	reg r_4013_0;
	reg r_4014_0;
	reg r_4015_0;
	reg r_4016_0;
	reg r_4017_0;
	reg r_4018_0;
	reg r_4019_0;
	reg r_4020_0;
	reg r_4021_0;
	reg r_4022_0;
	reg r_4023_0;
	reg r_4024_0;
	reg r_4025_0;
	reg r_4026_0;
	reg r_4027_0;
	reg r_4028_0;
	reg r_4029_0;
	reg r_4030_0;
	reg r_4031_0;
	reg r_4032_0;
	reg r_4033_0;
	reg r_4034_0;
	reg r_4035_0;
	reg r_4036_0;
	reg r_4037_0;
	reg r_4038_0;
	reg r_4039_0;
	reg r_4040_0;
	reg r_4041_0;
	reg r_4042_0;
	reg r_4043_0;
	reg r_4044_0;
	reg r_4045_0;
	reg r_4046_0;
	reg r_4047_0;
	reg r_4048_0;
	reg r_4049_0;
	reg r_4050_0;
	reg r_4051_0;
	reg r_4052_0;
	reg r_4053_0;
	reg r_4054_0;
	reg r_4055_0;
	reg r_4056_0;
	reg r_4057_0;
	reg r_4058_0;
	reg r_4059_0;
	reg r_4060_0;
	reg r_4061_0;
	reg r_4062_0;
	reg r_4063_0;
	reg r_4064_0;
	reg r_4065_0;
	reg r_4066_0;
	reg r_4067_0;
	reg r_4068_0;
	reg r_4069_0;
	reg r_4070_0;
	reg r_4071_0;
	reg r_4072_0;
	reg r_4073_0;
	reg r_4074_0;
	reg r_4075_0;
	reg r_4076_0;
	reg r_4077_0;
	reg r_4078_0;
	reg r_4079_0;
	reg r_4080_0;
	reg r_4081_0;
	reg r_4082_0;
	reg r_4083_0;
	reg r_4084_0;
	reg r_4085_0;
	reg r_4086_0;
	reg r_4087_0;
	reg r_4088_0;
	reg r_4089_0;
	reg r_4090_0;
	reg r_4091_0;
	reg r_4092_0;
	reg r_4093_0;
	reg r_4094_0;
	reg r_4095_0;
	reg [31:0] r_4096_0;
	reg [31:0] r_4097_0;
	reg r_4098_0;
	reg r_4099_0_dataflow;
	reg [2:0] r_4100_0;
	reg r_4101_0;
	reg [31:0] r_4102_0;
	reg [31:0] r_4103_0;
	reg [31:0] r_4108_0;
	reg [31:0] r_4109_0;
	reg [31:0] r_4114_0;
	reg [31:0] r_4115_0;
	reg [31:0] r_4120_0;
	reg [31:0] r_4121_0;
	reg [31:0] r_4126_0;
	reg [31:0] r_4127_0;
	reg [31:0] r_4132_0;
	reg [31:0] r_4133_0;
	reg [31:0] r_4138_0;
	reg [31:0] r_4139_0;
	reg [31:0] r_4144_0;
	reg [31:0] r_4145_0;
	reg [31:0] r_4150_0;
	reg [31:0] r_4151_0;
	reg [31:0] r_4156_0;
	reg [31:0] r_4157_0;
	reg [31:0] r_4162_0;
	reg [31:0] r_4163_0;
	reg [31:0] r_4168_0;
	reg [31:0] r_4169_0;
	reg [31:0] r_4174_0;
	reg [31:0] r_4175_0;
	reg [31:0] r_4180_0;
	reg [31:0] r_4181_0;
	reg [31:0] r_4186_0;
	reg [31:0] r_4187_0;
	reg [31:0] r_4192_0;
	reg [31:0] r_4193_0;
	reg [31:0] r_4198_0;
	reg [31:0] r_4199_0;
	reg [31:0] r_4204_0;
	reg [31:0] r_4205_0;
	reg [31:0] r_4210_0;
	reg [31:0] r_4211_0;
	reg [31:0] r_4216_0;
	reg [31:0] r_4217_0;
	reg [31:0] r_4222_0;
	reg [31:0] r_4223_0;
	reg [31:0] r_4228_0;
	reg [31:0] r_4229_0;
	reg [31:0] r_4234_0;
	reg [31:0] r_4235_0;
	reg [31:0] r_4240_0;
	reg [31:0] r_4241_0;
	reg [31:0] r_4246_0;
	reg [31:0] r_4247_0;
	reg [31:0] r_4252_0;
	reg [31:0] r_4253_0;
	reg [31:0] r_4258_0;
	reg [31:0] r_4259_0;
	reg [31:0] r_4264_0;
	reg [31:0] r_4265_0;
	reg [31:0] r_4270_0;
	reg [31:0] r_4271_0;
	reg [31:0] r_4276_0;
	reg [31:0] r_4277_0;
	reg [31:0] r_4282_0;
	reg [31:0] r_4283_0;
	always @(posedge clock) begin
		r_0 <=( io_in_a_0_0) ^ ((fiEnable && (17 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1_0 <=( _mesh_0_0_io_out_a_0) ^ ((fiEnable && (18 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_2_0 <=( _mesh_0_1_io_out_a_0) ^ ((fiEnable && (19 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_3_0 <=( _mesh_0_2_io_out_a_0) ^ ((fiEnable && (20 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4_0 <=( _mesh_0_3_io_out_a_0) ^ ((fiEnable && (21 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_5_0 <=( _mesh_0_4_io_out_a_0) ^ ((fiEnable && (22 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_6_0 <=( _mesh_0_5_io_out_a_0) ^ ((fiEnable && (23 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_7_0 <=( _mesh_0_6_io_out_a_0) ^ ((fiEnable && (24 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_8_0 <=( _mesh_0_7_io_out_a_0) ^ ((fiEnable && (25 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_9_0 <=( _mesh_0_8_io_out_a_0) ^ ((fiEnable && (26 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_10_0 <=( _mesh_0_9_io_out_a_0) ^ ((fiEnable && (27 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_11_0 <=( _mesh_0_10_io_out_a_0) ^ ((fiEnable && (28 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_12_0 <=( _mesh_0_11_io_out_a_0) ^ ((fiEnable && (29 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_13_0 <=( _mesh_0_12_io_out_a_0) ^ ((fiEnable && (30 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_14_0 <=( _mesh_0_13_io_out_a_0) ^ ((fiEnable && (31 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_15_0 <=( _mesh_0_14_io_out_a_0) ^ ((fiEnable && (32 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_16_0 <=( _mesh_0_15_io_out_a_0) ^ ((fiEnable && (33 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_17_0 <=( _mesh_0_16_io_out_a_0) ^ ((fiEnable && (34 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_18_0 <=( _mesh_0_17_io_out_a_0) ^ ((fiEnable && (35 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_19_0 <=( _mesh_0_18_io_out_a_0) ^ ((fiEnable && (36 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_20_0 <=( _mesh_0_19_io_out_a_0) ^ ((fiEnable && (37 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_21_0 <=( _mesh_0_20_io_out_a_0) ^ ((fiEnable && (38 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_22_0 <=( _mesh_0_21_io_out_a_0) ^ ((fiEnable && (39 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_23_0 <=( _mesh_0_22_io_out_a_0) ^ ((fiEnable && (40 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_24_0 <=( _mesh_0_23_io_out_a_0) ^ ((fiEnable && (41 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_25_0 <=( _mesh_0_24_io_out_a_0) ^ ((fiEnable && (42 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_26_0 <=( _mesh_0_25_io_out_a_0) ^ ((fiEnable && (43 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_27_0 <=( _mesh_0_26_io_out_a_0) ^ ((fiEnable && (44 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_28_0 <=( _mesh_0_27_io_out_a_0) ^ ((fiEnable && (45 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_29_0 <=( _mesh_0_28_io_out_a_0) ^ ((fiEnable && (46 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_30_0 <=( _mesh_0_29_io_out_a_0) ^ ((fiEnable && (47 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_31_0 <=( _mesh_0_30_io_out_a_0) ^ ((fiEnable && (48 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_32_0 <=( io_in_a_1_0) ^ ((fiEnable && (49 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_33_0 <=( _mesh_1_0_io_out_a_0) ^ ((fiEnable && (50 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_34_0 <=( _mesh_1_1_io_out_a_0) ^ ((fiEnable && (51 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_35_0 <=( _mesh_1_2_io_out_a_0) ^ ((fiEnable && (52 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_36_0 <=( _mesh_1_3_io_out_a_0) ^ ((fiEnable && (53 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_37_0 <=( _mesh_1_4_io_out_a_0) ^ ((fiEnable && (54 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_38_0 <=( _mesh_1_5_io_out_a_0) ^ ((fiEnable && (55 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_39_0 <=( _mesh_1_6_io_out_a_0) ^ ((fiEnable && (56 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_40_0 <=( _mesh_1_7_io_out_a_0) ^ ((fiEnable && (57 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_41_0 <=( _mesh_1_8_io_out_a_0) ^ ((fiEnable && (58 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_42_0 <=( _mesh_1_9_io_out_a_0) ^ ((fiEnable && (59 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_43_0 <=( _mesh_1_10_io_out_a_0) ^ ((fiEnable && (60 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_44_0 <=( _mesh_1_11_io_out_a_0) ^ ((fiEnable && (61 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_45_0 <=( _mesh_1_12_io_out_a_0) ^ ((fiEnable && (62 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_46_0 <=( _mesh_1_13_io_out_a_0) ^ ((fiEnable && (63 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_47_0 <=( _mesh_1_14_io_out_a_0) ^ ((fiEnable && (64 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_48_0 <=( _mesh_1_15_io_out_a_0) ^ ((fiEnable && (65 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_49_0 <=( _mesh_1_16_io_out_a_0) ^ ((fiEnable && (66 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_50_0 <=( _mesh_1_17_io_out_a_0) ^ ((fiEnable && (67 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_51_0 <=( _mesh_1_18_io_out_a_0) ^ ((fiEnable && (68 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_52_0 <=( _mesh_1_19_io_out_a_0) ^ ((fiEnable && (69 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_53_0 <=( _mesh_1_20_io_out_a_0) ^ ((fiEnable && (70 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_54_0 <=( _mesh_1_21_io_out_a_0) ^ ((fiEnable && (71 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_55_0 <=( _mesh_1_22_io_out_a_0) ^ ((fiEnable && (72 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_56_0 <=( _mesh_1_23_io_out_a_0) ^ ((fiEnable && (73 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_57_0 <=( _mesh_1_24_io_out_a_0) ^ ((fiEnable && (74 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_58_0 <=( _mesh_1_25_io_out_a_0) ^ ((fiEnable && (75 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_59_0 <=( _mesh_1_26_io_out_a_0) ^ ((fiEnable && (76 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_60_0 <=( _mesh_1_27_io_out_a_0) ^ ((fiEnable && (77 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_61_0 <=( _mesh_1_28_io_out_a_0) ^ ((fiEnable && (78 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_62_0 <=( _mesh_1_29_io_out_a_0) ^ ((fiEnable && (79 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_63_0 <=( _mesh_1_30_io_out_a_0) ^ ((fiEnable && (80 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_64_0 <=( io_in_a_2_0) ^ ((fiEnable && (81 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_65_0 <=( _mesh_2_0_io_out_a_0) ^ ((fiEnable && (82 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_66_0 <=( _mesh_2_1_io_out_a_0) ^ ((fiEnable && (83 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_67_0 <=( _mesh_2_2_io_out_a_0) ^ ((fiEnable && (84 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_68_0 <=( _mesh_2_3_io_out_a_0) ^ ((fiEnable && (85 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_69_0 <=( _mesh_2_4_io_out_a_0) ^ ((fiEnable && (86 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_70_0 <=( _mesh_2_5_io_out_a_0) ^ ((fiEnable && (87 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_71_0 <=( _mesh_2_6_io_out_a_0) ^ ((fiEnable && (88 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_72_0 <=( _mesh_2_7_io_out_a_0) ^ ((fiEnable && (89 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_73_0 <=( _mesh_2_8_io_out_a_0) ^ ((fiEnable && (90 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_74_0 <=( _mesh_2_9_io_out_a_0) ^ ((fiEnable && (91 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_75_0 <=( _mesh_2_10_io_out_a_0) ^ ((fiEnable && (92 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_76_0 <=( _mesh_2_11_io_out_a_0) ^ ((fiEnable && (93 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_77_0 <=( _mesh_2_12_io_out_a_0) ^ ((fiEnable && (94 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_78_0 <=( _mesh_2_13_io_out_a_0) ^ ((fiEnable && (95 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_79_0 <=( _mesh_2_14_io_out_a_0) ^ ((fiEnable && (96 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_80_0 <=( _mesh_2_15_io_out_a_0) ^ ((fiEnable && (97 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_81_0 <=( _mesh_2_16_io_out_a_0) ^ ((fiEnable && (98 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_82_0 <=( _mesh_2_17_io_out_a_0) ^ ((fiEnable && (99 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_83_0 <=( _mesh_2_18_io_out_a_0) ^ ((fiEnable && (100 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_84_0 <=( _mesh_2_19_io_out_a_0) ^ ((fiEnable && (101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_85_0 <=( _mesh_2_20_io_out_a_0) ^ ((fiEnable && (102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_86_0 <=( _mesh_2_21_io_out_a_0) ^ ((fiEnable && (103 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_87_0 <=( _mesh_2_22_io_out_a_0) ^ ((fiEnable && (104 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_88_0 <=( _mesh_2_23_io_out_a_0) ^ ((fiEnable && (105 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_89_0 <=( _mesh_2_24_io_out_a_0) ^ ((fiEnable && (106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_90_0 <=( _mesh_2_25_io_out_a_0) ^ ((fiEnable && (107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_91_0 <=( _mesh_2_26_io_out_a_0) ^ ((fiEnable && (108 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_92_0 <=( _mesh_2_27_io_out_a_0) ^ ((fiEnable && (109 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_93_0 <=( _mesh_2_28_io_out_a_0) ^ ((fiEnable && (110 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_94_0 <=( _mesh_2_29_io_out_a_0) ^ ((fiEnable && (111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_95_0 <=( _mesh_2_30_io_out_a_0) ^ ((fiEnable && (112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_96_0 <=( io_in_a_3_0) ^ ((fiEnable && (113 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_97_0 <=( _mesh_3_0_io_out_a_0) ^ ((fiEnable && (114 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_98_0 <=( _mesh_3_1_io_out_a_0) ^ ((fiEnable && (115 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_99_0 <=( _mesh_3_2_io_out_a_0) ^ ((fiEnable && (116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_100_0 <=( _mesh_3_3_io_out_a_0) ^ ((fiEnable && (117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_101_0 <=( _mesh_3_4_io_out_a_0) ^ ((fiEnable && (118 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_102_0 <=( _mesh_3_5_io_out_a_0) ^ ((fiEnable && (119 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_103_0 <=( _mesh_3_6_io_out_a_0) ^ ((fiEnable && (120 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_104_0 <=( _mesh_3_7_io_out_a_0) ^ ((fiEnable && (121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_105_0 <=( _mesh_3_8_io_out_a_0) ^ ((fiEnable && (122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_106_0 <=( _mesh_3_9_io_out_a_0) ^ ((fiEnable && (123 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_107_0 <=( _mesh_3_10_io_out_a_0) ^ ((fiEnable && (124 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_108_0 <=( _mesh_3_11_io_out_a_0) ^ ((fiEnable && (125 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_109_0 <=( _mesh_3_12_io_out_a_0) ^ ((fiEnable && (126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_110_0 <=( _mesh_3_13_io_out_a_0) ^ ((fiEnable && (127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_111_0 <=( _mesh_3_14_io_out_a_0) ^ ((fiEnable && (128 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_112_0 <=( _mesh_3_15_io_out_a_0) ^ ((fiEnable && (129 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_113_0 <=( _mesh_3_16_io_out_a_0) ^ ((fiEnable && (130 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_114_0 <=( _mesh_3_17_io_out_a_0) ^ ((fiEnable && (131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_115_0 <=( _mesh_3_18_io_out_a_0) ^ ((fiEnable && (132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_116_0 <=( _mesh_3_19_io_out_a_0) ^ ((fiEnable && (133 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_117_0 <=( _mesh_3_20_io_out_a_0) ^ ((fiEnable && (134 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_118_0 <=( _mesh_3_21_io_out_a_0) ^ ((fiEnable && (135 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_119_0 <=( _mesh_3_22_io_out_a_0) ^ ((fiEnable && (136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_120_0 <=( _mesh_3_23_io_out_a_0) ^ ((fiEnable && (137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_121_0 <=( _mesh_3_24_io_out_a_0) ^ ((fiEnable && (138 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_122_0 <=( _mesh_3_25_io_out_a_0) ^ ((fiEnable && (139 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_123_0 <=( _mesh_3_26_io_out_a_0) ^ ((fiEnable && (140 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_124_0 <=( _mesh_3_27_io_out_a_0) ^ ((fiEnable && (141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_125_0 <=( _mesh_3_28_io_out_a_0) ^ ((fiEnable && (142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_126_0 <=( _mesh_3_29_io_out_a_0) ^ ((fiEnable && (143 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_127_0 <=( _mesh_3_30_io_out_a_0) ^ ((fiEnable && (144 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_128_0 <=( io_in_a_4_0) ^ ((fiEnable && (145 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_129_0 <=( _mesh_4_0_io_out_a_0) ^ ((fiEnable && (146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_130_0 <=( _mesh_4_1_io_out_a_0) ^ ((fiEnable && (147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_131_0 <=( _mesh_4_2_io_out_a_0) ^ ((fiEnable && (148 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_132_0 <=( _mesh_4_3_io_out_a_0) ^ ((fiEnable && (149 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_133_0 <=( _mesh_4_4_io_out_a_0) ^ ((fiEnable && (150 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_134_0 <=( _mesh_4_5_io_out_a_0) ^ ((fiEnable && (151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_135_0 <=( _mesh_4_6_io_out_a_0) ^ ((fiEnable && (152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_136_0 <=( _mesh_4_7_io_out_a_0) ^ ((fiEnable && (153 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_137_0 <=( _mesh_4_8_io_out_a_0) ^ ((fiEnable && (154 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_138_0 <=( _mesh_4_9_io_out_a_0) ^ ((fiEnable && (155 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_139_0 <=( _mesh_4_10_io_out_a_0) ^ ((fiEnable && (156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_140_0 <=( _mesh_4_11_io_out_a_0) ^ ((fiEnable && (157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_141_0 <=( _mesh_4_12_io_out_a_0) ^ ((fiEnable && (158 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_142_0 <=( _mesh_4_13_io_out_a_0) ^ ((fiEnable && (159 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_143_0 <=( _mesh_4_14_io_out_a_0) ^ ((fiEnable && (160 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_144_0 <=( _mesh_4_15_io_out_a_0) ^ ((fiEnable && (161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_145_0 <=( _mesh_4_16_io_out_a_0) ^ ((fiEnable && (162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_146_0 <=( _mesh_4_17_io_out_a_0) ^ ((fiEnable && (163 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_147_0 <=( _mesh_4_18_io_out_a_0) ^ ((fiEnable && (164 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_148_0 <=( _mesh_4_19_io_out_a_0) ^ ((fiEnable && (165 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_149_0 <=( _mesh_4_20_io_out_a_0) ^ ((fiEnable && (166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_150_0 <=( _mesh_4_21_io_out_a_0) ^ ((fiEnable && (167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_151_0 <=( _mesh_4_22_io_out_a_0) ^ ((fiEnable && (168 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_152_0 <=( _mesh_4_23_io_out_a_0) ^ ((fiEnable && (169 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_153_0 <=( _mesh_4_24_io_out_a_0) ^ ((fiEnable && (170 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_154_0 <=( _mesh_4_25_io_out_a_0) ^ ((fiEnable && (171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_155_0 <=( _mesh_4_26_io_out_a_0) ^ ((fiEnable && (172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_156_0 <=( _mesh_4_27_io_out_a_0) ^ ((fiEnable && (173 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_157_0 <=( _mesh_4_28_io_out_a_0) ^ ((fiEnable && (174 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_158_0 <=( _mesh_4_29_io_out_a_0) ^ ((fiEnable && (175 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_159_0 <=( _mesh_4_30_io_out_a_0) ^ ((fiEnable && (176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_160_0 <=( io_in_a_5_0) ^ ((fiEnable && (177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_161_0 <=( _mesh_5_0_io_out_a_0) ^ ((fiEnable && (178 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_162_0 <=( _mesh_5_1_io_out_a_0) ^ ((fiEnable && (179 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_163_0 <=( _mesh_5_2_io_out_a_0) ^ ((fiEnable && (180 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_164_0 <=( _mesh_5_3_io_out_a_0) ^ ((fiEnable && (181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_165_0 <=( _mesh_5_4_io_out_a_0) ^ ((fiEnable && (182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_166_0 <=( _mesh_5_5_io_out_a_0) ^ ((fiEnable && (183 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_167_0 <=( _mesh_5_6_io_out_a_0) ^ ((fiEnable && (184 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_168_0 <=( _mesh_5_7_io_out_a_0) ^ ((fiEnable && (185 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_169_0 <=( _mesh_5_8_io_out_a_0) ^ ((fiEnable && (186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_170_0 <=( _mesh_5_9_io_out_a_0) ^ ((fiEnable && (187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_171_0 <=( _mesh_5_10_io_out_a_0) ^ ((fiEnable && (188 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_172_0 <=( _mesh_5_11_io_out_a_0) ^ ((fiEnable && (189 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_173_0 <=( _mesh_5_12_io_out_a_0) ^ ((fiEnable && (190 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_174_0 <=( _mesh_5_13_io_out_a_0) ^ ((fiEnable && (191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_175_0 <=( _mesh_5_14_io_out_a_0) ^ ((fiEnable && (192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_176_0 <=( _mesh_5_15_io_out_a_0) ^ ((fiEnable && (193 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_177_0 <=( _mesh_5_16_io_out_a_0) ^ ((fiEnable && (194 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_178_0 <=( _mesh_5_17_io_out_a_0) ^ ((fiEnable && (195 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_179_0 <=( _mesh_5_18_io_out_a_0) ^ ((fiEnable && (196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_180_0 <=( _mesh_5_19_io_out_a_0) ^ ((fiEnable && (197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_181_0 <=( _mesh_5_20_io_out_a_0) ^ ((fiEnable && (198 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_182_0 <=( _mesh_5_21_io_out_a_0) ^ ((fiEnable && (199 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_183_0 <=( _mesh_5_22_io_out_a_0) ^ ((fiEnable && (200 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_184_0 <=( _mesh_5_23_io_out_a_0) ^ ((fiEnable && (201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_185_0 <=( _mesh_5_24_io_out_a_0) ^ ((fiEnable && (202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_186_0 <=( _mesh_5_25_io_out_a_0) ^ ((fiEnable && (203 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_187_0 <=( _mesh_5_26_io_out_a_0) ^ ((fiEnable && (204 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_188_0 <=( _mesh_5_27_io_out_a_0) ^ ((fiEnable && (205 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_189_0 <=( _mesh_5_28_io_out_a_0) ^ ((fiEnable && (206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_190_0 <=( _mesh_5_29_io_out_a_0) ^ ((fiEnable && (207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_191_0 <=( _mesh_5_30_io_out_a_0) ^ ((fiEnable && (208 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_192_0 <=( io_in_a_6_0) ^ ((fiEnable && (209 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_193_0 <=( _mesh_6_0_io_out_a_0) ^ ((fiEnable && (210 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_194_0 <=( _mesh_6_1_io_out_a_0) ^ ((fiEnable && (211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_195_0 <=( _mesh_6_2_io_out_a_0) ^ ((fiEnable && (212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_196_0 <=( _mesh_6_3_io_out_a_0) ^ ((fiEnable && (213 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_197_0 <=( _mesh_6_4_io_out_a_0) ^ ((fiEnable && (214 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_198_0 <=( _mesh_6_5_io_out_a_0) ^ ((fiEnable && (215 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_199_0 <=( _mesh_6_6_io_out_a_0) ^ ((fiEnable && (216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_200_0 <=( _mesh_6_7_io_out_a_0) ^ ((fiEnable && (217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_201_0 <=( _mesh_6_8_io_out_a_0) ^ ((fiEnable && (218 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_202_0 <=( _mesh_6_9_io_out_a_0) ^ ((fiEnable && (219 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_203_0 <=( _mesh_6_10_io_out_a_0) ^ ((fiEnable && (220 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_204_0 <=( _mesh_6_11_io_out_a_0) ^ ((fiEnable && (221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_205_0 <=( _mesh_6_12_io_out_a_0) ^ ((fiEnable && (222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_206_0 <=( _mesh_6_13_io_out_a_0) ^ ((fiEnable && (223 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_207_0 <=( _mesh_6_14_io_out_a_0) ^ ((fiEnable && (224 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_208_0 <=( _mesh_6_15_io_out_a_0) ^ ((fiEnable && (225 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_209_0 <=( _mesh_6_16_io_out_a_0) ^ ((fiEnable && (226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_210_0 <=( _mesh_6_17_io_out_a_0) ^ ((fiEnable && (227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_211_0 <=( _mesh_6_18_io_out_a_0) ^ ((fiEnable && (228 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_212_0 <=( _mesh_6_19_io_out_a_0) ^ ((fiEnable && (229 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_213_0 <=( _mesh_6_20_io_out_a_0) ^ ((fiEnable && (230 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_214_0 <=( _mesh_6_21_io_out_a_0) ^ ((fiEnable && (231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_215_0 <=( _mesh_6_22_io_out_a_0) ^ ((fiEnable && (232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_216_0 <=( _mesh_6_23_io_out_a_0) ^ ((fiEnable && (233 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_217_0 <=( _mesh_6_24_io_out_a_0) ^ ((fiEnable && (234 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_218_0 <=( _mesh_6_25_io_out_a_0) ^ ((fiEnable && (235 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_219_0 <=( _mesh_6_26_io_out_a_0) ^ ((fiEnable && (236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_220_0 <=( _mesh_6_27_io_out_a_0) ^ ((fiEnable && (237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_221_0 <=( _mesh_6_28_io_out_a_0) ^ ((fiEnable && (238 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_222_0 <=( _mesh_6_29_io_out_a_0) ^ ((fiEnable && (239 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_223_0 <=( _mesh_6_30_io_out_a_0) ^ ((fiEnable && (240 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_224_0 <=( io_in_a_7_0) ^ ((fiEnable && (241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_225_0 <=( _mesh_7_0_io_out_a_0) ^ ((fiEnable && (242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_226_0 <=( _mesh_7_1_io_out_a_0) ^ ((fiEnable && (243 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_227_0 <=( _mesh_7_2_io_out_a_0) ^ ((fiEnable && (244 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_228_0 <=( _mesh_7_3_io_out_a_0) ^ ((fiEnable && (245 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_229_0 <=( _mesh_7_4_io_out_a_0) ^ ((fiEnable && (246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_230_0 <=( _mesh_7_5_io_out_a_0) ^ ((fiEnable && (247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_231_0 <=( _mesh_7_6_io_out_a_0) ^ ((fiEnable && (248 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_232_0 <=( _mesh_7_7_io_out_a_0) ^ ((fiEnable && (249 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_233_0 <=( _mesh_7_8_io_out_a_0) ^ ((fiEnable && (250 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_234_0 <=( _mesh_7_9_io_out_a_0) ^ ((fiEnable && (251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_235_0 <=( _mesh_7_10_io_out_a_0) ^ ((fiEnable && (252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_236_0 <=( _mesh_7_11_io_out_a_0) ^ ((fiEnable && (253 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_237_0 <=( _mesh_7_12_io_out_a_0) ^ ((fiEnable && (254 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_238_0 <=( _mesh_7_13_io_out_a_0) ^ ((fiEnable && (255 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_239_0 <=( _mesh_7_14_io_out_a_0) ^ ((fiEnable && (256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_240_0 <=( _mesh_7_15_io_out_a_0) ^ ((fiEnable && (257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_241_0 <=( _mesh_7_16_io_out_a_0) ^ ((fiEnable && (258 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_242_0 <=( _mesh_7_17_io_out_a_0) ^ ((fiEnable && (259 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_243_0 <=( _mesh_7_18_io_out_a_0) ^ ((fiEnable && (260 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_244_0 <=( _mesh_7_19_io_out_a_0) ^ ((fiEnable && (261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_245_0 <=( _mesh_7_20_io_out_a_0) ^ ((fiEnable && (262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_246_0 <=( _mesh_7_21_io_out_a_0) ^ ((fiEnable && (263 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_247_0 <=( _mesh_7_22_io_out_a_0) ^ ((fiEnable && (264 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_248_0 <=( _mesh_7_23_io_out_a_0) ^ ((fiEnable && (265 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_249_0 <=( _mesh_7_24_io_out_a_0) ^ ((fiEnable && (266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_250_0 <=( _mesh_7_25_io_out_a_0) ^ ((fiEnable && (267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_251_0 <=( _mesh_7_26_io_out_a_0) ^ ((fiEnable && (268 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_252_0 <=( _mesh_7_27_io_out_a_0) ^ ((fiEnable && (269 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_253_0 <=( _mesh_7_28_io_out_a_0) ^ ((fiEnable && (270 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_254_0 <=( _mesh_7_29_io_out_a_0) ^ ((fiEnable && (271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_255_0 <=( _mesh_7_30_io_out_a_0) ^ ((fiEnable && (272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_256_0 <=( io_in_a_8_0) ^ ((fiEnable && (273 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_257_0 <=( _mesh_8_0_io_out_a_0) ^ ((fiEnable && (274 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_258_0 <=( _mesh_8_1_io_out_a_0) ^ ((fiEnable && (275 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_259_0 <=( _mesh_8_2_io_out_a_0) ^ ((fiEnable && (276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_260_0 <=( _mesh_8_3_io_out_a_0) ^ ((fiEnable && (277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_261_0 <=( _mesh_8_4_io_out_a_0) ^ ((fiEnable && (278 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_262_0 <=( _mesh_8_5_io_out_a_0) ^ ((fiEnable && (279 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_263_0 <=( _mesh_8_6_io_out_a_0) ^ ((fiEnable && (280 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_264_0 <=( _mesh_8_7_io_out_a_0) ^ ((fiEnable && (281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_265_0 <=( _mesh_8_8_io_out_a_0) ^ ((fiEnable && (282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_266_0 <=( _mesh_8_9_io_out_a_0) ^ ((fiEnable && (283 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_267_0 <=( _mesh_8_10_io_out_a_0) ^ ((fiEnable && (284 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_268_0 <=( _mesh_8_11_io_out_a_0) ^ ((fiEnable && (285 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_269_0 <=( _mesh_8_12_io_out_a_0) ^ ((fiEnable && (286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_270_0 <=( _mesh_8_13_io_out_a_0) ^ ((fiEnable && (287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_271_0 <=( _mesh_8_14_io_out_a_0) ^ ((fiEnable && (288 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_272_0 <=( _mesh_8_15_io_out_a_0) ^ ((fiEnable && (289 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_273_0 <=( _mesh_8_16_io_out_a_0) ^ ((fiEnable && (290 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_274_0 <=( _mesh_8_17_io_out_a_0) ^ ((fiEnable && (291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_275_0 <=( _mesh_8_18_io_out_a_0) ^ ((fiEnable && (292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_276_0 <=( _mesh_8_19_io_out_a_0) ^ ((fiEnable && (293 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_277_0 <=( _mesh_8_20_io_out_a_0) ^ ((fiEnable && (294 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_278_0 <=( _mesh_8_21_io_out_a_0) ^ ((fiEnable && (295 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_279_0 <=( _mesh_8_22_io_out_a_0) ^ ((fiEnable && (296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_280_0 <=( _mesh_8_23_io_out_a_0) ^ ((fiEnable && (297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_281_0 <=( _mesh_8_24_io_out_a_0) ^ ((fiEnable && (298 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_282_0 <=( _mesh_8_25_io_out_a_0) ^ ((fiEnable && (299 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_283_0 <=( _mesh_8_26_io_out_a_0) ^ ((fiEnable && (300 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_284_0 <=( _mesh_8_27_io_out_a_0) ^ ((fiEnable && (301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_285_0 <=( _mesh_8_28_io_out_a_0) ^ ((fiEnable && (302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_286_0 <=( _mesh_8_29_io_out_a_0) ^ ((fiEnable && (303 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_287_0 <=( _mesh_8_30_io_out_a_0) ^ ((fiEnable && (304 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_288_0 <=( io_in_a_9_0) ^ ((fiEnable && (305 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_289_0 <=( _mesh_9_0_io_out_a_0) ^ ((fiEnable && (306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_290_0 <=( _mesh_9_1_io_out_a_0) ^ ((fiEnable && (307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_291_0 <=( _mesh_9_2_io_out_a_0) ^ ((fiEnable && (308 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_292_0 <=( _mesh_9_3_io_out_a_0) ^ ((fiEnable && (309 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_293_0 <=( _mesh_9_4_io_out_a_0) ^ ((fiEnable && (310 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_294_0 <=( _mesh_9_5_io_out_a_0) ^ ((fiEnable && (311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_295_0 <=( _mesh_9_6_io_out_a_0) ^ ((fiEnable && (312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_296_0 <=( _mesh_9_7_io_out_a_0) ^ ((fiEnable && (313 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_297_0 <=( _mesh_9_8_io_out_a_0) ^ ((fiEnable && (314 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_298_0 <=( _mesh_9_9_io_out_a_0) ^ ((fiEnable && (315 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_299_0 <=( _mesh_9_10_io_out_a_0) ^ ((fiEnable && (316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_300_0 <=( _mesh_9_11_io_out_a_0) ^ ((fiEnable && (317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_301_0 <=( _mesh_9_12_io_out_a_0) ^ ((fiEnable && (318 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_302_0 <=( _mesh_9_13_io_out_a_0) ^ ((fiEnable && (319 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_303_0 <=( _mesh_9_14_io_out_a_0) ^ ((fiEnable && (320 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_304_0 <=( _mesh_9_15_io_out_a_0) ^ ((fiEnable && (321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_305_0 <=( _mesh_9_16_io_out_a_0) ^ ((fiEnable && (322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_306_0 <=( _mesh_9_17_io_out_a_0) ^ ((fiEnable && (323 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_307_0 <=( _mesh_9_18_io_out_a_0) ^ ((fiEnable && (324 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_308_0 <=( _mesh_9_19_io_out_a_0) ^ ((fiEnable && (325 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_309_0 <=( _mesh_9_20_io_out_a_0) ^ ((fiEnable && (326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_310_0 <=( _mesh_9_21_io_out_a_0) ^ ((fiEnable && (327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_311_0 <=( _mesh_9_22_io_out_a_0) ^ ((fiEnable && (328 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_312_0 <=( _mesh_9_23_io_out_a_0) ^ ((fiEnable && (329 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_313_0 <=( _mesh_9_24_io_out_a_0) ^ ((fiEnable && (330 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_314_0 <=( _mesh_9_25_io_out_a_0) ^ ((fiEnable && (331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_315_0 <=( _mesh_9_26_io_out_a_0) ^ ((fiEnable && (332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_316_0 <=( _mesh_9_27_io_out_a_0) ^ ((fiEnable && (333 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_317_0 <=( _mesh_9_28_io_out_a_0) ^ ((fiEnable && (334 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_318_0 <=( _mesh_9_29_io_out_a_0) ^ ((fiEnable && (335 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_319_0 <=( _mesh_9_30_io_out_a_0) ^ ((fiEnable && (336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_320_0 <=( io_in_a_10_0) ^ ((fiEnable && (337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_321_0 <=( _mesh_10_0_io_out_a_0) ^ ((fiEnable && (338 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_322_0 <=( _mesh_10_1_io_out_a_0) ^ ((fiEnable && (339 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_323_0 <=( _mesh_10_2_io_out_a_0) ^ ((fiEnable && (340 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_324_0 <=( _mesh_10_3_io_out_a_0) ^ ((fiEnable && (341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_325_0 <=( _mesh_10_4_io_out_a_0) ^ ((fiEnable && (342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_326_0 <=( _mesh_10_5_io_out_a_0) ^ ((fiEnable && (343 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_327_0 <=( _mesh_10_6_io_out_a_0) ^ ((fiEnable && (344 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_328_0 <=( _mesh_10_7_io_out_a_0) ^ ((fiEnable && (345 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_329_0 <=( _mesh_10_8_io_out_a_0) ^ ((fiEnable && (346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_330_0 <=( _mesh_10_9_io_out_a_0) ^ ((fiEnable && (347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_331_0 <=( _mesh_10_10_io_out_a_0) ^ ((fiEnable && (348 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_332_0 <=( _mesh_10_11_io_out_a_0) ^ ((fiEnable && (349 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_333_0 <=( _mesh_10_12_io_out_a_0) ^ ((fiEnable && (350 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_334_0 <=( _mesh_10_13_io_out_a_0) ^ ((fiEnable && (351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_335_0 <=( _mesh_10_14_io_out_a_0) ^ ((fiEnable && (352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_336_0 <=( _mesh_10_15_io_out_a_0) ^ ((fiEnable && (353 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_337_0 <=( _mesh_10_16_io_out_a_0) ^ ((fiEnable && (354 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_338_0 <=( _mesh_10_17_io_out_a_0) ^ ((fiEnable && (355 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_339_0 <=( _mesh_10_18_io_out_a_0) ^ ((fiEnable && (356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_340_0 <=( _mesh_10_19_io_out_a_0) ^ ((fiEnable && (357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_341_0 <=( _mesh_10_20_io_out_a_0) ^ ((fiEnable && (358 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_342_0 <=( _mesh_10_21_io_out_a_0) ^ ((fiEnable && (359 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_343_0 <=( _mesh_10_22_io_out_a_0) ^ ((fiEnable && (360 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_344_0 <=( _mesh_10_23_io_out_a_0) ^ ((fiEnable && (361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_345_0 <=( _mesh_10_24_io_out_a_0) ^ ((fiEnable && (362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_346_0 <=( _mesh_10_25_io_out_a_0) ^ ((fiEnable && (363 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_347_0 <=( _mesh_10_26_io_out_a_0) ^ ((fiEnable && (364 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_348_0 <=( _mesh_10_27_io_out_a_0) ^ ((fiEnable && (365 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_349_0 <=( _mesh_10_28_io_out_a_0) ^ ((fiEnable && (366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_350_0 <=( _mesh_10_29_io_out_a_0) ^ ((fiEnable && (367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_351_0 <=( _mesh_10_30_io_out_a_0) ^ ((fiEnable && (368 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_352_0 <=( io_in_a_11_0) ^ ((fiEnable && (369 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_353_0 <=( _mesh_11_0_io_out_a_0) ^ ((fiEnable && (370 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_354_0 <=( _mesh_11_1_io_out_a_0) ^ ((fiEnable && (371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_355_0 <=( _mesh_11_2_io_out_a_0) ^ ((fiEnable && (372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_356_0 <=( _mesh_11_3_io_out_a_0) ^ ((fiEnable && (373 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_357_0 <=( _mesh_11_4_io_out_a_0) ^ ((fiEnable && (374 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_358_0 <=( _mesh_11_5_io_out_a_0) ^ ((fiEnable && (375 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_359_0 <=( _mesh_11_6_io_out_a_0) ^ ((fiEnable && (376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_360_0 <=( _mesh_11_7_io_out_a_0) ^ ((fiEnable && (377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_361_0 <=( _mesh_11_8_io_out_a_0) ^ ((fiEnable && (378 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_362_0 <=( _mesh_11_9_io_out_a_0) ^ ((fiEnable && (379 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_363_0 <=( _mesh_11_10_io_out_a_0) ^ ((fiEnable && (380 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_364_0 <=( _mesh_11_11_io_out_a_0) ^ ((fiEnable && (381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_365_0 <=( _mesh_11_12_io_out_a_0) ^ ((fiEnable && (382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_366_0 <=( _mesh_11_13_io_out_a_0) ^ ((fiEnable && (383 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_367_0 <=( _mesh_11_14_io_out_a_0) ^ ((fiEnable && (384 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_368_0 <=( _mesh_11_15_io_out_a_0) ^ ((fiEnable && (385 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_369_0 <=( _mesh_11_16_io_out_a_0) ^ ((fiEnable && (386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_370_0 <=( _mesh_11_17_io_out_a_0) ^ ((fiEnable && (387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_371_0 <=( _mesh_11_18_io_out_a_0) ^ ((fiEnable && (388 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_372_0 <=( _mesh_11_19_io_out_a_0) ^ ((fiEnable && (389 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_373_0 <=( _mesh_11_20_io_out_a_0) ^ ((fiEnable && (390 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_374_0 <=( _mesh_11_21_io_out_a_0) ^ ((fiEnable && (391 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_375_0 <=( _mesh_11_22_io_out_a_0) ^ ((fiEnable && (392 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_376_0 <=( _mesh_11_23_io_out_a_0) ^ ((fiEnable && (393 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_377_0 <=( _mesh_11_24_io_out_a_0) ^ ((fiEnable && (394 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_378_0 <=( _mesh_11_25_io_out_a_0) ^ ((fiEnable && (395 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_379_0 <=( _mesh_11_26_io_out_a_0) ^ ((fiEnable && (396 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_380_0 <=( _mesh_11_27_io_out_a_0) ^ ((fiEnable && (397 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_381_0 <=( _mesh_11_28_io_out_a_0) ^ ((fiEnable && (398 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_382_0 <=( _mesh_11_29_io_out_a_0) ^ ((fiEnable && (399 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_383_0 <=( _mesh_11_30_io_out_a_0) ^ ((fiEnable && (400 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_384_0 <=( io_in_a_12_0) ^ ((fiEnable && (401 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_385_0 <=( _mesh_12_0_io_out_a_0) ^ ((fiEnable && (402 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_386_0 <=( _mesh_12_1_io_out_a_0) ^ ((fiEnable && (403 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_387_0 <=( _mesh_12_2_io_out_a_0) ^ ((fiEnable && (404 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_388_0 <=( _mesh_12_3_io_out_a_0) ^ ((fiEnable && (405 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_389_0 <=( _mesh_12_4_io_out_a_0) ^ ((fiEnable && (406 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_390_0 <=( _mesh_12_5_io_out_a_0) ^ ((fiEnable && (407 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_391_0 <=( _mesh_12_6_io_out_a_0) ^ ((fiEnable && (408 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_392_0 <=( _mesh_12_7_io_out_a_0) ^ ((fiEnable && (409 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_393_0 <=( _mesh_12_8_io_out_a_0) ^ ((fiEnable && (410 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_394_0 <=( _mesh_12_9_io_out_a_0) ^ ((fiEnable && (411 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_395_0 <=( _mesh_12_10_io_out_a_0) ^ ((fiEnable && (412 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_396_0 <=( _mesh_12_11_io_out_a_0) ^ ((fiEnable && (413 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_397_0 <=( _mesh_12_12_io_out_a_0) ^ ((fiEnable && (414 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_398_0 <=( _mesh_12_13_io_out_a_0) ^ ((fiEnable && (415 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_399_0 <=( _mesh_12_14_io_out_a_0) ^ ((fiEnable && (416 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_400_0 <=( _mesh_12_15_io_out_a_0) ^ ((fiEnable && (417 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_401_0 <=( _mesh_12_16_io_out_a_0) ^ ((fiEnable && (418 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_402_0 <=( _mesh_12_17_io_out_a_0) ^ ((fiEnable && (419 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_403_0 <=( _mesh_12_18_io_out_a_0) ^ ((fiEnable && (420 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_404_0 <=( _mesh_12_19_io_out_a_0) ^ ((fiEnable && (421 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_405_0 <=( _mesh_12_20_io_out_a_0) ^ ((fiEnable && (422 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_406_0 <=( _mesh_12_21_io_out_a_0) ^ ((fiEnable && (423 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_407_0 <=( _mesh_12_22_io_out_a_0) ^ ((fiEnable && (424 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_408_0 <=( _mesh_12_23_io_out_a_0) ^ ((fiEnable && (425 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_409_0 <=( _mesh_12_24_io_out_a_0) ^ ((fiEnable && (426 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_410_0 <=( _mesh_12_25_io_out_a_0) ^ ((fiEnable && (427 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_411_0 <=( _mesh_12_26_io_out_a_0) ^ ((fiEnable && (428 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_412_0 <=( _mesh_12_27_io_out_a_0) ^ ((fiEnable && (429 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_413_0 <=( _mesh_12_28_io_out_a_0) ^ ((fiEnable && (430 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_414_0 <=( _mesh_12_29_io_out_a_0) ^ ((fiEnable && (431 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_415_0 <=( _mesh_12_30_io_out_a_0) ^ ((fiEnable && (432 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_416_0 <=( io_in_a_13_0) ^ ((fiEnable && (433 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_417_0 <=( _mesh_13_0_io_out_a_0) ^ ((fiEnable && (434 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_418_0 <=( _mesh_13_1_io_out_a_0) ^ ((fiEnable && (435 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_419_0 <=( _mesh_13_2_io_out_a_0) ^ ((fiEnable && (436 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_420_0 <=( _mesh_13_3_io_out_a_0) ^ ((fiEnable && (437 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_421_0 <=( _mesh_13_4_io_out_a_0) ^ ((fiEnable && (438 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_422_0 <=( _mesh_13_5_io_out_a_0) ^ ((fiEnable && (439 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_423_0 <=( _mesh_13_6_io_out_a_0) ^ ((fiEnable && (440 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_424_0 <=( _mesh_13_7_io_out_a_0) ^ ((fiEnable && (441 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_425_0 <=( _mesh_13_8_io_out_a_0) ^ ((fiEnable && (442 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_426_0 <=( _mesh_13_9_io_out_a_0) ^ ((fiEnable && (443 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_427_0 <=( _mesh_13_10_io_out_a_0) ^ ((fiEnable && (444 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_428_0 <=( _mesh_13_11_io_out_a_0) ^ ((fiEnable && (445 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_429_0 <=( _mesh_13_12_io_out_a_0) ^ ((fiEnable && (446 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_430_0 <=( _mesh_13_13_io_out_a_0) ^ ((fiEnable && (447 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_431_0 <=( _mesh_13_14_io_out_a_0) ^ ((fiEnable && (448 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_432_0 <=( _mesh_13_15_io_out_a_0) ^ ((fiEnable && (449 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_433_0 <=( _mesh_13_16_io_out_a_0) ^ ((fiEnable && (450 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_434_0 <=( _mesh_13_17_io_out_a_0) ^ ((fiEnable && (451 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_435_0 <=( _mesh_13_18_io_out_a_0) ^ ((fiEnable && (452 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_436_0 <=( _mesh_13_19_io_out_a_0) ^ ((fiEnable && (453 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_437_0 <=( _mesh_13_20_io_out_a_0) ^ ((fiEnable && (454 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_438_0 <=( _mesh_13_21_io_out_a_0) ^ ((fiEnable && (455 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_439_0 <=( _mesh_13_22_io_out_a_0) ^ ((fiEnable && (456 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_440_0 <=( _mesh_13_23_io_out_a_0) ^ ((fiEnable && (457 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_441_0 <=( _mesh_13_24_io_out_a_0) ^ ((fiEnable && (458 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_442_0 <=( _mesh_13_25_io_out_a_0) ^ ((fiEnable && (459 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_443_0 <=( _mesh_13_26_io_out_a_0) ^ ((fiEnable && (460 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_444_0 <=( _mesh_13_27_io_out_a_0) ^ ((fiEnable && (461 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_445_0 <=( _mesh_13_28_io_out_a_0) ^ ((fiEnable && (462 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_446_0 <=( _mesh_13_29_io_out_a_0) ^ ((fiEnable && (463 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_447_0 <=( _mesh_13_30_io_out_a_0) ^ ((fiEnable && (464 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_448_0 <=( io_in_a_14_0) ^ ((fiEnable && (465 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_449_0 <=( _mesh_14_0_io_out_a_0) ^ ((fiEnable && (466 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_450_0 <=( _mesh_14_1_io_out_a_0) ^ ((fiEnable && (467 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_451_0 <=( _mesh_14_2_io_out_a_0) ^ ((fiEnable && (468 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_452_0 <=( _mesh_14_3_io_out_a_0) ^ ((fiEnable && (469 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_453_0 <=( _mesh_14_4_io_out_a_0) ^ ((fiEnable && (470 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_454_0 <=( _mesh_14_5_io_out_a_0) ^ ((fiEnable && (471 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_455_0 <=( _mesh_14_6_io_out_a_0) ^ ((fiEnable && (472 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_456_0 <=( _mesh_14_7_io_out_a_0) ^ ((fiEnable && (473 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_457_0 <=( _mesh_14_8_io_out_a_0) ^ ((fiEnable && (474 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_458_0 <=( _mesh_14_9_io_out_a_0) ^ ((fiEnable && (475 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_459_0 <=( _mesh_14_10_io_out_a_0) ^ ((fiEnable && (476 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_460_0 <=( _mesh_14_11_io_out_a_0) ^ ((fiEnable && (477 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_461_0 <=( _mesh_14_12_io_out_a_0) ^ ((fiEnable && (478 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_462_0 <=( _mesh_14_13_io_out_a_0) ^ ((fiEnable && (479 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_463_0 <=( _mesh_14_14_io_out_a_0) ^ ((fiEnable && (480 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_464_0 <=( _mesh_14_15_io_out_a_0) ^ ((fiEnable && (481 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_465_0 <=( _mesh_14_16_io_out_a_0) ^ ((fiEnable && (482 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_466_0 <=( _mesh_14_17_io_out_a_0) ^ ((fiEnable && (483 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_467_0 <=( _mesh_14_18_io_out_a_0) ^ ((fiEnable && (484 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_468_0 <=( _mesh_14_19_io_out_a_0) ^ ((fiEnable && (485 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_469_0 <=( _mesh_14_20_io_out_a_0) ^ ((fiEnable && (486 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_470_0 <=( _mesh_14_21_io_out_a_0) ^ ((fiEnable && (487 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_471_0 <=( _mesh_14_22_io_out_a_0) ^ ((fiEnable && (488 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_472_0 <=( _mesh_14_23_io_out_a_0) ^ ((fiEnable && (489 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_473_0 <=( _mesh_14_24_io_out_a_0) ^ ((fiEnable && (490 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_474_0 <=( _mesh_14_25_io_out_a_0) ^ ((fiEnable && (491 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_475_0 <=( _mesh_14_26_io_out_a_0) ^ ((fiEnable && (492 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_476_0 <=( _mesh_14_27_io_out_a_0) ^ ((fiEnable && (493 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_477_0 <=( _mesh_14_28_io_out_a_0) ^ ((fiEnable && (494 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_478_0 <=( _mesh_14_29_io_out_a_0) ^ ((fiEnable && (495 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_479_0 <=( _mesh_14_30_io_out_a_0) ^ ((fiEnable && (496 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_480_0 <=( io_in_a_15_0) ^ ((fiEnable && (497 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_481_0 <=( _mesh_15_0_io_out_a_0) ^ ((fiEnable && (498 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_482_0 <=( _mesh_15_1_io_out_a_0) ^ ((fiEnable && (499 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_483_0 <=( _mesh_15_2_io_out_a_0) ^ ((fiEnable && (500 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_484_0 <=( _mesh_15_3_io_out_a_0) ^ ((fiEnable && (501 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_485_0 <=( _mesh_15_4_io_out_a_0) ^ ((fiEnable && (502 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_486_0 <=( _mesh_15_5_io_out_a_0) ^ ((fiEnable && (503 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_487_0 <=( _mesh_15_6_io_out_a_0) ^ ((fiEnable && (504 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_488_0 <=( _mesh_15_7_io_out_a_0) ^ ((fiEnable && (505 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_489_0 <=( _mesh_15_8_io_out_a_0) ^ ((fiEnable && (506 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_490_0 <=( _mesh_15_9_io_out_a_0) ^ ((fiEnable && (507 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_491_0 <=( _mesh_15_10_io_out_a_0) ^ ((fiEnable && (508 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_492_0 <=( _mesh_15_11_io_out_a_0) ^ ((fiEnable && (509 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_493_0 <=( _mesh_15_12_io_out_a_0) ^ ((fiEnable && (510 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_494_0 <=( _mesh_15_13_io_out_a_0) ^ ((fiEnable && (511 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_495_0 <=( _mesh_15_14_io_out_a_0) ^ ((fiEnable && (512 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_496_0 <=( _mesh_15_15_io_out_a_0) ^ ((fiEnable && (513 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_497_0 <=( _mesh_15_16_io_out_a_0) ^ ((fiEnable && (514 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_498_0 <=( _mesh_15_17_io_out_a_0) ^ ((fiEnable && (515 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_499_0 <=( _mesh_15_18_io_out_a_0) ^ ((fiEnable && (516 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_500_0 <=( _mesh_15_19_io_out_a_0) ^ ((fiEnable && (517 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_501_0 <=( _mesh_15_20_io_out_a_0) ^ ((fiEnable && (518 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_502_0 <=( _mesh_15_21_io_out_a_0) ^ ((fiEnable && (519 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_503_0 <=( _mesh_15_22_io_out_a_0) ^ ((fiEnable && (520 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_504_0 <=( _mesh_15_23_io_out_a_0) ^ ((fiEnable && (521 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_505_0 <=( _mesh_15_24_io_out_a_0) ^ ((fiEnable && (522 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_506_0 <=( _mesh_15_25_io_out_a_0) ^ ((fiEnable && (523 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_507_0 <=( _mesh_15_26_io_out_a_0) ^ ((fiEnable && (524 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_508_0 <=( _mesh_15_27_io_out_a_0) ^ ((fiEnable && (525 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_509_0 <=( _mesh_15_28_io_out_a_0) ^ ((fiEnable && (526 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_510_0 <=( _mesh_15_29_io_out_a_0) ^ ((fiEnable && (527 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_511_0 <=( _mesh_15_30_io_out_a_0) ^ ((fiEnable && (528 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_512_0 <=( io_in_a_16_0) ^ ((fiEnable && (529 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_513_0 <=( _mesh_16_0_io_out_a_0) ^ ((fiEnable && (530 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_514_0 <=( _mesh_16_1_io_out_a_0) ^ ((fiEnable && (531 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_515_0 <=( _mesh_16_2_io_out_a_0) ^ ((fiEnable && (532 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_516_0 <=( _mesh_16_3_io_out_a_0) ^ ((fiEnable && (533 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_517_0 <=( _mesh_16_4_io_out_a_0) ^ ((fiEnable && (534 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_518_0 <=( _mesh_16_5_io_out_a_0) ^ ((fiEnable && (535 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_519_0 <=( _mesh_16_6_io_out_a_0) ^ ((fiEnable && (536 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_520_0 <=( _mesh_16_7_io_out_a_0) ^ ((fiEnable && (537 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_521_0 <=( _mesh_16_8_io_out_a_0) ^ ((fiEnable && (538 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_522_0 <=( _mesh_16_9_io_out_a_0) ^ ((fiEnable && (539 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_523_0 <=( _mesh_16_10_io_out_a_0) ^ ((fiEnable && (540 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_524_0 <=( _mesh_16_11_io_out_a_0) ^ ((fiEnable && (541 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_525_0 <=( _mesh_16_12_io_out_a_0) ^ ((fiEnable && (542 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_526_0 <=( _mesh_16_13_io_out_a_0) ^ ((fiEnable && (543 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_527_0 <=( _mesh_16_14_io_out_a_0) ^ ((fiEnable && (544 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_528_0 <=( _mesh_16_15_io_out_a_0) ^ ((fiEnable && (545 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_529_0 <=( _mesh_16_16_io_out_a_0) ^ ((fiEnable && (546 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_530_0 <=( _mesh_16_17_io_out_a_0) ^ ((fiEnable && (547 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_531_0 <=( _mesh_16_18_io_out_a_0) ^ ((fiEnable && (548 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_532_0 <=( _mesh_16_19_io_out_a_0) ^ ((fiEnable && (549 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_533_0 <=( _mesh_16_20_io_out_a_0) ^ ((fiEnable && (550 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_534_0 <=( _mesh_16_21_io_out_a_0) ^ ((fiEnable && (551 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_535_0 <=( _mesh_16_22_io_out_a_0) ^ ((fiEnable && (552 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_536_0 <=( _mesh_16_23_io_out_a_0) ^ ((fiEnable && (553 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_537_0 <=( _mesh_16_24_io_out_a_0) ^ ((fiEnable && (554 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_538_0 <=( _mesh_16_25_io_out_a_0) ^ ((fiEnable && (555 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_539_0 <=( _mesh_16_26_io_out_a_0) ^ ((fiEnable && (556 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_540_0 <=( _mesh_16_27_io_out_a_0) ^ ((fiEnable && (557 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_541_0 <=( _mesh_16_28_io_out_a_0) ^ ((fiEnable && (558 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_542_0 <=( _mesh_16_29_io_out_a_0) ^ ((fiEnable && (559 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_543_0 <=( _mesh_16_30_io_out_a_0) ^ ((fiEnable && (560 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_544_0 <=( io_in_a_17_0) ^ ((fiEnable && (561 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_545_0 <=( _mesh_17_0_io_out_a_0) ^ ((fiEnable && (562 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_546_0 <=( _mesh_17_1_io_out_a_0) ^ ((fiEnable && (563 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_547_0 <=( _mesh_17_2_io_out_a_0) ^ ((fiEnable && (564 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_548_0 <=( _mesh_17_3_io_out_a_0) ^ ((fiEnable && (565 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_549_0 <=( _mesh_17_4_io_out_a_0) ^ ((fiEnable && (566 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_550_0 <=( _mesh_17_5_io_out_a_0) ^ ((fiEnable && (567 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_551_0 <=( _mesh_17_6_io_out_a_0) ^ ((fiEnable && (568 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_552_0 <=( _mesh_17_7_io_out_a_0) ^ ((fiEnable && (569 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_553_0 <=( _mesh_17_8_io_out_a_0) ^ ((fiEnable && (570 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_554_0 <=( _mesh_17_9_io_out_a_0) ^ ((fiEnable && (571 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_555_0 <=( _mesh_17_10_io_out_a_0) ^ ((fiEnable && (572 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_556_0 <=( _mesh_17_11_io_out_a_0) ^ ((fiEnable && (573 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_557_0 <=( _mesh_17_12_io_out_a_0) ^ ((fiEnable && (574 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_558_0 <=( _mesh_17_13_io_out_a_0) ^ ((fiEnable && (575 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_559_0 <=( _mesh_17_14_io_out_a_0) ^ ((fiEnable && (576 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_560_0 <=( _mesh_17_15_io_out_a_0) ^ ((fiEnable && (577 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_561_0 <=( _mesh_17_16_io_out_a_0) ^ ((fiEnable && (578 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_562_0 <=( _mesh_17_17_io_out_a_0) ^ ((fiEnable && (579 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_563_0 <=( _mesh_17_18_io_out_a_0) ^ ((fiEnable && (580 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_564_0 <=( _mesh_17_19_io_out_a_0) ^ ((fiEnable && (581 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_565_0 <=( _mesh_17_20_io_out_a_0) ^ ((fiEnable && (582 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_566_0 <=( _mesh_17_21_io_out_a_0) ^ ((fiEnable && (583 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_567_0 <=( _mesh_17_22_io_out_a_0) ^ ((fiEnable && (584 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_568_0 <=( _mesh_17_23_io_out_a_0) ^ ((fiEnable && (585 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_569_0 <=( _mesh_17_24_io_out_a_0) ^ ((fiEnable && (586 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_570_0 <=( _mesh_17_25_io_out_a_0) ^ ((fiEnable && (587 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_571_0 <=( _mesh_17_26_io_out_a_0) ^ ((fiEnable && (588 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_572_0 <=( _mesh_17_27_io_out_a_0) ^ ((fiEnable && (589 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_573_0 <=( _mesh_17_28_io_out_a_0) ^ ((fiEnable && (590 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_574_0 <=( _mesh_17_29_io_out_a_0) ^ ((fiEnable && (591 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_575_0 <=( _mesh_17_30_io_out_a_0) ^ ((fiEnable && (592 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_576_0 <=( io_in_a_18_0) ^ ((fiEnable && (593 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_577_0 <=( _mesh_18_0_io_out_a_0) ^ ((fiEnable && (594 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_578_0 <=( _mesh_18_1_io_out_a_0) ^ ((fiEnable && (595 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_579_0 <=( _mesh_18_2_io_out_a_0) ^ ((fiEnable && (596 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_580_0 <=( _mesh_18_3_io_out_a_0) ^ ((fiEnable && (597 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_581_0 <=( _mesh_18_4_io_out_a_0) ^ ((fiEnable && (598 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_582_0 <=( _mesh_18_5_io_out_a_0) ^ ((fiEnable && (599 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_583_0 <=( _mesh_18_6_io_out_a_0) ^ ((fiEnable && (600 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_584_0 <=( _mesh_18_7_io_out_a_0) ^ ((fiEnable && (601 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_585_0 <=( _mesh_18_8_io_out_a_0) ^ ((fiEnable && (602 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_586_0 <=( _mesh_18_9_io_out_a_0) ^ ((fiEnable && (603 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_587_0 <=( _mesh_18_10_io_out_a_0) ^ ((fiEnable && (604 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_588_0 <=( _mesh_18_11_io_out_a_0) ^ ((fiEnable && (605 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_589_0 <=( _mesh_18_12_io_out_a_0) ^ ((fiEnable && (606 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_590_0 <=( _mesh_18_13_io_out_a_0) ^ ((fiEnable && (607 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_591_0 <=( _mesh_18_14_io_out_a_0) ^ ((fiEnable && (608 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_592_0 <=( _mesh_18_15_io_out_a_0) ^ ((fiEnable && (609 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_593_0 <=( _mesh_18_16_io_out_a_0) ^ ((fiEnable && (610 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_594_0 <=( _mesh_18_17_io_out_a_0) ^ ((fiEnable && (611 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_595_0 <=( _mesh_18_18_io_out_a_0) ^ ((fiEnable && (612 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_596_0 <=( _mesh_18_19_io_out_a_0) ^ ((fiEnable && (613 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_597_0 <=( _mesh_18_20_io_out_a_0) ^ ((fiEnable && (614 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_598_0 <=( _mesh_18_21_io_out_a_0) ^ ((fiEnable && (615 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_599_0 <=( _mesh_18_22_io_out_a_0) ^ ((fiEnable && (616 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_600_0 <=( _mesh_18_23_io_out_a_0) ^ ((fiEnable && (617 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_601_0 <=( _mesh_18_24_io_out_a_0) ^ ((fiEnable && (618 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_602_0 <=( _mesh_18_25_io_out_a_0) ^ ((fiEnable && (619 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_603_0 <=( _mesh_18_26_io_out_a_0) ^ ((fiEnable && (620 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_604_0 <=( _mesh_18_27_io_out_a_0) ^ ((fiEnable && (621 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_605_0 <=( _mesh_18_28_io_out_a_0) ^ ((fiEnable && (622 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_606_0 <=( _mesh_18_29_io_out_a_0) ^ ((fiEnable && (623 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_607_0 <=( _mesh_18_30_io_out_a_0) ^ ((fiEnable && (624 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_608_0 <=( io_in_a_19_0) ^ ((fiEnable && (625 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_609_0 <=( _mesh_19_0_io_out_a_0) ^ ((fiEnable && (626 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_610_0 <=( _mesh_19_1_io_out_a_0) ^ ((fiEnable && (627 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_611_0 <=( _mesh_19_2_io_out_a_0) ^ ((fiEnable && (628 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_612_0 <=( _mesh_19_3_io_out_a_0) ^ ((fiEnable && (629 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_613_0 <=( _mesh_19_4_io_out_a_0) ^ ((fiEnable && (630 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_614_0 <=( _mesh_19_5_io_out_a_0) ^ ((fiEnable && (631 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_615_0 <=( _mesh_19_6_io_out_a_0) ^ ((fiEnable && (632 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_616_0 <=( _mesh_19_7_io_out_a_0) ^ ((fiEnable && (633 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_617_0 <=( _mesh_19_8_io_out_a_0) ^ ((fiEnable && (634 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_618_0 <=( _mesh_19_9_io_out_a_0) ^ ((fiEnable && (635 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_619_0 <=( _mesh_19_10_io_out_a_0) ^ ((fiEnable && (636 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_620_0 <=( _mesh_19_11_io_out_a_0) ^ ((fiEnable && (637 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_621_0 <=( _mesh_19_12_io_out_a_0) ^ ((fiEnable && (638 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_622_0 <=( _mesh_19_13_io_out_a_0) ^ ((fiEnable && (639 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_623_0 <=( _mesh_19_14_io_out_a_0) ^ ((fiEnable && (640 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_624_0 <=( _mesh_19_15_io_out_a_0) ^ ((fiEnable && (641 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_625_0 <=( _mesh_19_16_io_out_a_0) ^ ((fiEnable && (642 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_626_0 <=( _mesh_19_17_io_out_a_0) ^ ((fiEnable && (643 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_627_0 <=( _mesh_19_18_io_out_a_0) ^ ((fiEnable && (644 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_628_0 <=( _mesh_19_19_io_out_a_0) ^ ((fiEnable && (645 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_629_0 <=( _mesh_19_20_io_out_a_0) ^ ((fiEnable && (646 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_630_0 <=( _mesh_19_21_io_out_a_0) ^ ((fiEnable && (647 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_631_0 <=( _mesh_19_22_io_out_a_0) ^ ((fiEnable && (648 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_632_0 <=( _mesh_19_23_io_out_a_0) ^ ((fiEnable && (649 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_633_0 <=( _mesh_19_24_io_out_a_0) ^ ((fiEnable && (650 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_634_0 <=( _mesh_19_25_io_out_a_0) ^ ((fiEnable && (651 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_635_0 <=( _mesh_19_26_io_out_a_0) ^ ((fiEnable && (652 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_636_0 <=( _mesh_19_27_io_out_a_0) ^ ((fiEnable && (653 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_637_0 <=( _mesh_19_28_io_out_a_0) ^ ((fiEnable && (654 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_638_0 <=( _mesh_19_29_io_out_a_0) ^ ((fiEnable && (655 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_639_0 <=( _mesh_19_30_io_out_a_0) ^ ((fiEnable && (656 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_640_0 <=( io_in_a_20_0) ^ ((fiEnable && (657 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_641_0 <=( _mesh_20_0_io_out_a_0) ^ ((fiEnable && (658 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_642_0 <=( _mesh_20_1_io_out_a_0) ^ ((fiEnable && (659 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_643_0 <=( _mesh_20_2_io_out_a_0) ^ ((fiEnable && (660 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_644_0 <=( _mesh_20_3_io_out_a_0) ^ ((fiEnable && (661 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_645_0 <=( _mesh_20_4_io_out_a_0) ^ ((fiEnable && (662 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_646_0 <=( _mesh_20_5_io_out_a_0) ^ ((fiEnable && (663 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_647_0 <=( _mesh_20_6_io_out_a_0) ^ ((fiEnable && (664 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_648_0 <=( _mesh_20_7_io_out_a_0) ^ ((fiEnable && (665 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_649_0 <=( _mesh_20_8_io_out_a_0) ^ ((fiEnable && (666 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_650_0 <=( _mesh_20_9_io_out_a_0) ^ ((fiEnable && (667 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_651_0 <=( _mesh_20_10_io_out_a_0) ^ ((fiEnable && (668 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_652_0 <=( _mesh_20_11_io_out_a_0) ^ ((fiEnable && (669 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_653_0 <=( _mesh_20_12_io_out_a_0) ^ ((fiEnable && (670 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_654_0 <=( _mesh_20_13_io_out_a_0) ^ ((fiEnable && (671 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_655_0 <=( _mesh_20_14_io_out_a_0) ^ ((fiEnable && (672 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_656_0 <=( _mesh_20_15_io_out_a_0) ^ ((fiEnable && (673 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_657_0 <=( _mesh_20_16_io_out_a_0) ^ ((fiEnable && (674 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_658_0 <=( _mesh_20_17_io_out_a_0) ^ ((fiEnable && (675 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_659_0 <=( _mesh_20_18_io_out_a_0) ^ ((fiEnable && (676 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_660_0 <=( _mesh_20_19_io_out_a_0) ^ ((fiEnable && (677 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_661_0 <=( _mesh_20_20_io_out_a_0) ^ ((fiEnable && (678 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_662_0 <=( _mesh_20_21_io_out_a_0) ^ ((fiEnable && (679 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_663_0 <=( _mesh_20_22_io_out_a_0) ^ ((fiEnable && (680 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_664_0 <=( _mesh_20_23_io_out_a_0) ^ ((fiEnable && (681 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_665_0 <=( _mesh_20_24_io_out_a_0) ^ ((fiEnable && (682 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_666_0 <=( _mesh_20_25_io_out_a_0) ^ ((fiEnable && (683 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_667_0 <=( _mesh_20_26_io_out_a_0) ^ ((fiEnable && (684 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_668_0 <=( _mesh_20_27_io_out_a_0) ^ ((fiEnable && (685 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_669_0 <=( _mesh_20_28_io_out_a_0) ^ ((fiEnable && (686 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_670_0 <=( _mesh_20_29_io_out_a_0) ^ ((fiEnable && (687 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_671_0 <=( _mesh_20_30_io_out_a_0) ^ ((fiEnable && (688 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_672_0 <=( io_in_a_21_0) ^ ((fiEnable && (689 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_673_0 <=( _mesh_21_0_io_out_a_0) ^ ((fiEnable && (690 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_674_0 <=( _mesh_21_1_io_out_a_0) ^ ((fiEnable && (691 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_675_0 <=( _mesh_21_2_io_out_a_0) ^ ((fiEnable && (692 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_676_0 <=( _mesh_21_3_io_out_a_0) ^ ((fiEnable && (693 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_677_0 <=( _mesh_21_4_io_out_a_0) ^ ((fiEnable && (694 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_678_0 <=( _mesh_21_5_io_out_a_0) ^ ((fiEnable && (695 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_679_0 <=( _mesh_21_6_io_out_a_0) ^ ((fiEnable && (696 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_680_0 <=( _mesh_21_7_io_out_a_0) ^ ((fiEnable && (697 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_681_0 <=( _mesh_21_8_io_out_a_0) ^ ((fiEnable && (698 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_682_0 <=( _mesh_21_9_io_out_a_0) ^ ((fiEnable && (699 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_683_0 <=( _mesh_21_10_io_out_a_0) ^ ((fiEnable && (700 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_684_0 <=( _mesh_21_11_io_out_a_0) ^ ((fiEnable && (701 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_685_0 <=( _mesh_21_12_io_out_a_0) ^ ((fiEnable && (702 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_686_0 <=( _mesh_21_13_io_out_a_0) ^ ((fiEnable && (703 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_687_0 <=( _mesh_21_14_io_out_a_0) ^ ((fiEnable && (704 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_688_0 <=( _mesh_21_15_io_out_a_0) ^ ((fiEnable && (705 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_689_0 <=( _mesh_21_16_io_out_a_0) ^ ((fiEnable && (706 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_690_0 <=( _mesh_21_17_io_out_a_0) ^ ((fiEnable && (707 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_691_0 <=( _mesh_21_18_io_out_a_0) ^ ((fiEnable && (708 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_692_0 <=( _mesh_21_19_io_out_a_0) ^ ((fiEnable && (709 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_693_0 <=( _mesh_21_20_io_out_a_0) ^ ((fiEnable && (710 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_694_0 <=( _mesh_21_21_io_out_a_0) ^ ((fiEnable && (711 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_695_0 <=( _mesh_21_22_io_out_a_0) ^ ((fiEnable && (712 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_696_0 <=( _mesh_21_23_io_out_a_0) ^ ((fiEnable && (713 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_697_0 <=( _mesh_21_24_io_out_a_0) ^ ((fiEnable && (714 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_698_0 <=( _mesh_21_25_io_out_a_0) ^ ((fiEnable && (715 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_699_0 <=( _mesh_21_26_io_out_a_0) ^ ((fiEnable && (716 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_700_0 <=( _mesh_21_27_io_out_a_0) ^ ((fiEnable && (717 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_701_0 <=( _mesh_21_28_io_out_a_0) ^ ((fiEnable && (718 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_702_0 <=( _mesh_21_29_io_out_a_0) ^ ((fiEnable && (719 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_703_0 <=( _mesh_21_30_io_out_a_0) ^ ((fiEnable && (720 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_704_0 <=( io_in_a_22_0) ^ ((fiEnable && (721 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_705_0 <=( _mesh_22_0_io_out_a_0) ^ ((fiEnable && (722 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_706_0 <=( _mesh_22_1_io_out_a_0) ^ ((fiEnable && (723 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_707_0 <=( _mesh_22_2_io_out_a_0) ^ ((fiEnable && (724 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_708_0 <=( _mesh_22_3_io_out_a_0) ^ ((fiEnable && (725 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_709_0 <=( _mesh_22_4_io_out_a_0) ^ ((fiEnable && (726 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_710_0 <=( _mesh_22_5_io_out_a_0) ^ ((fiEnable && (727 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_711_0 <=( _mesh_22_6_io_out_a_0) ^ ((fiEnable && (728 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_712_0 <=( _mesh_22_7_io_out_a_0) ^ ((fiEnable && (729 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_713_0 <=( _mesh_22_8_io_out_a_0) ^ ((fiEnable && (730 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_714_0 <=( _mesh_22_9_io_out_a_0) ^ ((fiEnable && (731 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_715_0 <=( _mesh_22_10_io_out_a_0) ^ ((fiEnable && (732 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_716_0 <=( _mesh_22_11_io_out_a_0) ^ ((fiEnable && (733 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_717_0 <=( _mesh_22_12_io_out_a_0) ^ ((fiEnable && (734 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_718_0 <=( _mesh_22_13_io_out_a_0) ^ ((fiEnable && (735 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_719_0 <=( _mesh_22_14_io_out_a_0) ^ ((fiEnable && (736 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_720_0 <=( _mesh_22_15_io_out_a_0) ^ ((fiEnable && (737 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_721_0 <=( _mesh_22_16_io_out_a_0) ^ ((fiEnable && (738 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_722_0 <=( _mesh_22_17_io_out_a_0) ^ ((fiEnable && (739 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_723_0 <=( _mesh_22_18_io_out_a_0) ^ ((fiEnable && (740 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_724_0 <=( _mesh_22_19_io_out_a_0) ^ ((fiEnable && (741 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_725_0 <=( _mesh_22_20_io_out_a_0) ^ ((fiEnable && (742 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_726_0 <=( _mesh_22_21_io_out_a_0) ^ ((fiEnable && (743 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_727_0 <=( _mesh_22_22_io_out_a_0) ^ ((fiEnable && (744 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_728_0 <=( _mesh_22_23_io_out_a_0) ^ ((fiEnable && (745 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_729_0 <=( _mesh_22_24_io_out_a_0) ^ ((fiEnable && (746 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_730_0 <=( _mesh_22_25_io_out_a_0) ^ ((fiEnable && (747 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_731_0 <=( _mesh_22_26_io_out_a_0) ^ ((fiEnable && (748 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_732_0 <=( _mesh_22_27_io_out_a_0) ^ ((fiEnable && (749 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_733_0 <=( _mesh_22_28_io_out_a_0) ^ ((fiEnable && (750 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_734_0 <=( _mesh_22_29_io_out_a_0) ^ ((fiEnable && (751 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_735_0 <=( _mesh_22_30_io_out_a_0) ^ ((fiEnable && (752 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_736_0 <=( io_in_a_23_0) ^ ((fiEnable && (753 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_737_0 <=( _mesh_23_0_io_out_a_0) ^ ((fiEnable && (754 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_738_0 <=( _mesh_23_1_io_out_a_0) ^ ((fiEnable && (755 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_739_0 <=( _mesh_23_2_io_out_a_0) ^ ((fiEnable && (756 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_740_0 <=( _mesh_23_3_io_out_a_0) ^ ((fiEnable && (757 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_741_0 <=( _mesh_23_4_io_out_a_0) ^ ((fiEnable && (758 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_742_0 <=( _mesh_23_5_io_out_a_0) ^ ((fiEnable && (759 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_743_0 <=( _mesh_23_6_io_out_a_0) ^ ((fiEnable && (760 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_744_0 <=( _mesh_23_7_io_out_a_0) ^ ((fiEnable && (761 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_745_0 <=( _mesh_23_8_io_out_a_0) ^ ((fiEnable && (762 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_746_0 <=( _mesh_23_9_io_out_a_0) ^ ((fiEnable && (763 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_747_0 <=( _mesh_23_10_io_out_a_0) ^ ((fiEnable && (764 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_748_0 <=( _mesh_23_11_io_out_a_0) ^ ((fiEnable && (765 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_749_0 <=( _mesh_23_12_io_out_a_0) ^ ((fiEnable && (766 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_750_0 <=( _mesh_23_13_io_out_a_0) ^ ((fiEnable && (767 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_751_0 <=( _mesh_23_14_io_out_a_0) ^ ((fiEnable && (768 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_752_0 <=( _mesh_23_15_io_out_a_0) ^ ((fiEnable && (769 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_753_0 <=( _mesh_23_16_io_out_a_0) ^ ((fiEnable && (770 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_754_0 <=( _mesh_23_17_io_out_a_0) ^ ((fiEnable && (771 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_755_0 <=( _mesh_23_18_io_out_a_0) ^ ((fiEnable && (772 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_756_0 <=( _mesh_23_19_io_out_a_0) ^ ((fiEnable && (773 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_757_0 <=( _mesh_23_20_io_out_a_0) ^ ((fiEnable && (774 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_758_0 <=( _mesh_23_21_io_out_a_0) ^ ((fiEnable && (775 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_759_0 <=( _mesh_23_22_io_out_a_0) ^ ((fiEnable && (776 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_760_0 <=( _mesh_23_23_io_out_a_0) ^ ((fiEnable && (777 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_761_0 <=( _mesh_23_24_io_out_a_0) ^ ((fiEnable && (778 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_762_0 <=( _mesh_23_25_io_out_a_0) ^ ((fiEnable && (779 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_763_0 <=( _mesh_23_26_io_out_a_0) ^ ((fiEnable && (780 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_764_0 <=( _mesh_23_27_io_out_a_0) ^ ((fiEnable && (781 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_765_0 <=( _mesh_23_28_io_out_a_0) ^ ((fiEnable && (782 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_766_0 <=( _mesh_23_29_io_out_a_0) ^ ((fiEnable && (783 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_767_0 <=( _mesh_23_30_io_out_a_0) ^ ((fiEnable && (784 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_768_0 <=( io_in_a_24_0) ^ ((fiEnable && (785 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_769_0 <=( _mesh_24_0_io_out_a_0) ^ ((fiEnable && (786 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_770_0 <=( _mesh_24_1_io_out_a_0) ^ ((fiEnable && (787 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_771_0 <=( _mesh_24_2_io_out_a_0) ^ ((fiEnable && (788 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_772_0 <=( _mesh_24_3_io_out_a_0) ^ ((fiEnable && (789 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_773_0 <=( _mesh_24_4_io_out_a_0) ^ ((fiEnable && (790 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_774_0 <=( _mesh_24_5_io_out_a_0) ^ ((fiEnable && (791 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_775_0 <=( _mesh_24_6_io_out_a_0) ^ ((fiEnable && (792 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_776_0 <=( _mesh_24_7_io_out_a_0) ^ ((fiEnable && (793 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_777_0 <=( _mesh_24_8_io_out_a_0) ^ ((fiEnable && (794 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_778_0 <=( _mesh_24_9_io_out_a_0) ^ ((fiEnable && (795 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_779_0 <=( _mesh_24_10_io_out_a_0) ^ ((fiEnable && (796 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_780_0 <=( _mesh_24_11_io_out_a_0) ^ ((fiEnable && (797 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_781_0 <=( _mesh_24_12_io_out_a_0) ^ ((fiEnable && (798 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_782_0 <=( _mesh_24_13_io_out_a_0) ^ ((fiEnable && (799 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_783_0 <=( _mesh_24_14_io_out_a_0) ^ ((fiEnable && (800 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_784_0 <=( _mesh_24_15_io_out_a_0) ^ ((fiEnable && (801 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_785_0 <=( _mesh_24_16_io_out_a_0) ^ ((fiEnable && (802 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_786_0 <=( _mesh_24_17_io_out_a_0) ^ ((fiEnable && (803 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_787_0 <=( _mesh_24_18_io_out_a_0) ^ ((fiEnable && (804 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_788_0 <=( _mesh_24_19_io_out_a_0) ^ ((fiEnable && (805 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_789_0 <=( _mesh_24_20_io_out_a_0) ^ ((fiEnable && (806 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_790_0 <=( _mesh_24_21_io_out_a_0) ^ ((fiEnable && (807 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_791_0 <=( _mesh_24_22_io_out_a_0) ^ ((fiEnable && (808 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_792_0 <=( _mesh_24_23_io_out_a_0) ^ ((fiEnable && (809 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_793_0 <=( _mesh_24_24_io_out_a_0) ^ ((fiEnable && (810 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_794_0 <=( _mesh_24_25_io_out_a_0) ^ ((fiEnable && (811 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_795_0 <=( _mesh_24_26_io_out_a_0) ^ ((fiEnable && (812 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_796_0 <=( _mesh_24_27_io_out_a_0) ^ ((fiEnable && (813 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_797_0 <=( _mesh_24_28_io_out_a_0) ^ ((fiEnable && (814 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_798_0 <=( _mesh_24_29_io_out_a_0) ^ ((fiEnable && (815 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_799_0 <=( _mesh_24_30_io_out_a_0) ^ ((fiEnable && (816 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_800_0 <=( io_in_a_25_0) ^ ((fiEnable && (817 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_801_0 <=( _mesh_25_0_io_out_a_0) ^ ((fiEnable && (818 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_802_0 <=( _mesh_25_1_io_out_a_0) ^ ((fiEnable && (819 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_803_0 <=( _mesh_25_2_io_out_a_0) ^ ((fiEnable && (820 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_804_0 <=( _mesh_25_3_io_out_a_0) ^ ((fiEnable && (821 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_805_0 <=( _mesh_25_4_io_out_a_0) ^ ((fiEnable && (822 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_806_0 <=( _mesh_25_5_io_out_a_0) ^ ((fiEnable && (823 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_807_0 <=( _mesh_25_6_io_out_a_0) ^ ((fiEnable && (824 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_808_0 <=( _mesh_25_7_io_out_a_0) ^ ((fiEnable && (825 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_809_0 <=( _mesh_25_8_io_out_a_0) ^ ((fiEnable && (826 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_810_0 <=( _mesh_25_9_io_out_a_0) ^ ((fiEnable && (827 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_811_0 <=( _mesh_25_10_io_out_a_0) ^ ((fiEnable && (828 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_812_0 <=( _mesh_25_11_io_out_a_0) ^ ((fiEnable && (829 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_813_0 <=( _mesh_25_12_io_out_a_0) ^ ((fiEnable && (830 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_814_0 <=( _mesh_25_13_io_out_a_0) ^ ((fiEnable && (831 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_815_0 <=( _mesh_25_14_io_out_a_0) ^ ((fiEnable && (832 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_816_0 <=( _mesh_25_15_io_out_a_0) ^ ((fiEnable && (833 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_817_0 <=( _mesh_25_16_io_out_a_0) ^ ((fiEnable && (834 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_818_0 <=( _mesh_25_17_io_out_a_0) ^ ((fiEnable && (835 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_819_0 <=( _mesh_25_18_io_out_a_0) ^ ((fiEnable && (836 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_820_0 <=( _mesh_25_19_io_out_a_0) ^ ((fiEnable && (837 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_821_0 <=( _mesh_25_20_io_out_a_0) ^ ((fiEnable && (838 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_822_0 <=( _mesh_25_21_io_out_a_0) ^ ((fiEnable && (839 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_823_0 <=( _mesh_25_22_io_out_a_0) ^ ((fiEnable && (840 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_824_0 <=( _mesh_25_23_io_out_a_0) ^ ((fiEnable && (841 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_825_0 <=( _mesh_25_24_io_out_a_0) ^ ((fiEnable && (842 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_826_0 <=( _mesh_25_25_io_out_a_0) ^ ((fiEnable && (843 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_827_0 <=( _mesh_25_26_io_out_a_0) ^ ((fiEnable && (844 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_828_0 <=( _mesh_25_27_io_out_a_0) ^ ((fiEnable && (845 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_829_0 <=( _mesh_25_28_io_out_a_0) ^ ((fiEnable && (846 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_830_0 <=( _mesh_25_29_io_out_a_0) ^ ((fiEnable && (847 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_831_0 <=( _mesh_25_30_io_out_a_0) ^ ((fiEnable && (848 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_832_0 <=( io_in_a_26_0) ^ ((fiEnable && (849 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_833_0 <=( _mesh_26_0_io_out_a_0) ^ ((fiEnable && (850 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_834_0 <=( _mesh_26_1_io_out_a_0) ^ ((fiEnable && (851 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_835_0 <=( _mesh_26_2_io_out_a_0) ^ ((fiEnable && (852 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_836_0 <=( _mesh_26_3_io_out_a_0) ^ ((fiEnable && (853 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_837_0 <=( _mesh_26_4_io_out_a_0) ^ ((fiEnable && (854 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_838_0 <=( _mesh_26_5_io_out_a_0) ^ ((fiEnable && (855 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_839_0 <=( _mesh_26_6_io_out_a_0) ^ ((fiEnable && (856 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_840_0 <=( _mesh_26_7_io_out_a_0) ^ ((fiEnable && (857 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_841_0 <=( _mesh_26_8_io_out_a_0) ^ ((fiEnable && (858 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_842_0 <=( _mesh_26_9_io_out_a_0) ^ ((fiEnable && (859 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_843_0 <=( _mesh_26_10_io_out_a_0) ^ ((fiEnable && (860 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_844_0 <=( _mesh_26_11_io_out_a_0) ^ ((fiEnable && (861 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_845_0 <=( _mesh_26_12_io_out_a_0) ^ ((fiEnable && (862 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_846_0 <=( _mesh_26_13_io_out_a_0) ^ ((fiEnable && (863 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_847_0 <=( _mesh_26_14_io_out_a_0) ^ ((fiEnable && (864 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_848_0 <=( _mesh_26_15_io_out_a_0) ^ ((fiEnable && (865 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_849_0 <=( _mesh_26_16_io_out_a_0) ^ ((fiEnable && (866 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_850_0 <=( _mesh_26_17_io_out_a_0) ^ ((fiEnable && (867 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_851_0 <=( _mesh_26_18_io_out_a_0) ^ ((fiEnable && (868 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_852_0 <=( _mesh_26_19_io_out_a_0) ^ ((fiEnable && (869 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_853_0 <=( _mesh_26_20_io_out_a_0) ^ ((fiEnable && (870 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_854_0 <=( _mesh_26_21_io_out_a_0) ^ ((fiEnable && (871 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_855_0 <=( _mesh_26_22_io_out_a_0) ^ ((fiEnable && (872 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_856_0 <=( _mesh_26_23_io_out_a_0) ^ ((fiEnable && (873 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_857_0 <=( _mesh_26_24_io_out_a_0) ^ ((fiEnable && (874 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_858_0 <=( _mesh_26_25_io_out_a_0) ^ ((fiEnable && (875 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_859_0 <=( _mesh_26_26_io_out_a_0) ^ ((fiEnable && (876 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_860_0 <=( _mesh_26_27_io_out_a_0) ^ ((fiEnable && (877 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_861_0 <=( _mesh_26_28_io_out_a_0) ^ ((fiEnable && (878 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_862_0 <=( _mesh_26_29_io_out_a_0) ^ ((fiEnable && (879 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_863_0 <=( _mesh_26_30_io_out_a_0) ^ ((fiEnable && (880 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_864_0 <=( io_in_a_27_0) ^ ((fiEnable && (881 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_865_0 <=( _mesh_27_0_io_out_a_0) ^ ((fiEnable && (882 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_866_0 <=( _mesh_27_1_io_out_a_0) ^ ((fiEnable && (883 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_867_0 <=( _mesh_27_2_io_out_a_0) ^ ((fiEnable && (884 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_868_0 <=( _mesh_27_3_io_out_a_0) ^ ((fiEnable && (885 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_869_0 <=( _mesh_27_4_io_out_a_0) ^ ((fiEnable && (886 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_870_0 <=( _mesh_27_5_io_out_a_0) ^ ((fiEnable && (887 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_871_0 <=( _mesh_27_6_io_out_a_0) ^ ((fiEnable && (888 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_872_0 <=( _mesh_27_7_io_out_a_0) ^ ((fiEnable && (889 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_873_0 <=( _mesh_27_8_io_out_a_0) ^ ((fiEnable && (890 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_874_0 <=( _mesh_27_9_io_out_a_0) ^ ((fiEnable && (891 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_875_0 <=( _mesh_27_10_io_out_a_0) ^ ((fiEnable && (892 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_876_0 <=( _mesh_27_11_io_out_a_0) ^ ((fiEnable && (893 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_877_0 <=( _mesh_27_12_io_out_a_0) ^ ((fiEnable && (894 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_878_0 <=( _mesh_27_13_io_out_a_0) ^ ((fiEnable && (895 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_879_0 <=( _mesh_27_14_io_out_a_0) ^ ((fiEnable && (896 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_880_0 <=( _mesh_27_15_io_out_a_0) ^ ((fiEnable && (897 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_881_0 <=( _mesh_27_16_io_out_a_0) ^ ((fiEnable && (898 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_882_0 <=( _mesh_27_17_io_out_a_0) ^ ((fiEnable && (899 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_883_0 <=( _mesh_27_18_io_out_a_0) ^ ((fiEnable && (900 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_884_0 <=( _mesh_27_19_io_out_a_0) ^ ((fiEnable && (901 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_885_0 <=( _mesh_27_20_io_out_a_0) ^ ((fiEnable && (902 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_886_0 <=( _mesh_27_21_io_out_a_0) ^ ((fiEnable && (903 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_887_0 <=( _mesh_27_22_io_out_a_0) ^ ((fiEnable && (904 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_888_0 <=( _mesh_27_23_io_out_a_0) ^ ((fiEnable && (905 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_889_0 <=( _mesh_27_24_io_out_a_0) ^ ((fiEnable && (906 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_890_0 <=( _mesh_27_25_io_out_a_0) ^ ((fiEnable && (907 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_891_0 <=( _mesh_27_26_io_out_a_0) ^ ((fiEnable && (908 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_892_0 <=( _mesh_27_27_io_out_a_0) ^ ((fiEnable && (909 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_893_0 <=( _mesh_27_28_io_out_a_0) ^ ((fiEnable && (910 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_894_0 <=( _mesh_27_29_io_out_a_0) ^ ((fiEnable && (911 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_895_0 <=( _mesh_27_30_io_out_a_0) ^ ((fiEnable && (912 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_896_0 <=( io_in_a_28_0) ^ ((fiEnable && (913 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_897_0 <=( _mesh_28_0_io_out_a_0) ^ ((fiEnable && (914 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_898_0 <=( _mesh_28_1_io_out_a_0) ^ ((fiEnable && (915 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_899_0 <=( _mesh_28_2_io_out_a_0) ^ ((fiEnable && (916 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_900_0 <=( _mesh_28_3_io_out_a_0) ^ ((fiEnable && (917 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_901_0 <=( _mesh_28_4_io_out_a_0) ^ ((fiEnable && (918 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_902_0 <=( _mesh_28_5_io_out_a_0) ^ ((fiEnable && (919 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_903_0 <=( _mesh_28_6_io_out_a_0) ^ ((fiEnable && (920 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_904_0 <=( _mesh_28_7_io_out_a_0) ^ ((fiEnable && (921 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_905_0 <=( _mesh_28_8_io_out_a_0) ^ ((fiEnable && (922 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_906_0 <=( _mesh_28_9_io_out_a_0) ^ ((fiEnable && (923 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_907_0 <=( _mesh_28_10_io_out_a_0) ^ ((fiEnable && (924 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_908_0 <=( _mesh_28_11_io_out_a_0) ^ ((fiEnable && (925 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_909_0 <=( _mesh_28_12_io_out_a_0) ^ ((fiEnable && (926 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_910_0 <=( _mesh_28_13_io_out_a_0) ^ ((fiEnable && (927 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_911_0 <=( _mesh_28_14_io_out_a_0) ^ ((fiEnable && (928 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_912_0 <=( _mesh_28_15_io_out_a_0) ^ ((fiEnable && (929 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_913_0 <=( _mesh_28_16_io_out_a_0) ^ ((fiEnable && (930 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_914_0 <=( _mesh_28_17_io_out_a_0) ^ ((fiEnable && (931 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_915_0 <=( _mesh_28_18_io_out_a_0) ^ ((fiEnable && (932 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_916_0 <=( _mesh_28_19_io_out_a_0) ^ ((fiEnable && (933 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_917_0 <=( _mesh_28_20_io_out_a_0) ^ ((fiEnable && (934 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_918_0 <=( _mesh_28_21_io_out_a_0) ^ ((fiEnable && (935 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_919_0 <=( _mesh_28_22_io_out_a_0) ^ ((fiEnable && (936 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_920_0 <=( _mesh_28_23_io_out_a_0) ^ ((fiEnable && (937 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_921_0 <=( _mesh_28_24_io_out_a_0) ^ ((fiEnable && (938 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_922_0 <=( _mesh_28_25_io_out_a_0) ^ ((fiEnable && (939 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_923_0 <=( _mesh_28_26_io_out_a_0) ^ ((fiEnable && (940 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_924_0 <=( _mesh_28_27_io_out_a_0) ^ ((fiEnable && (941 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_925_0 <=( _mesh_28_28_io_out_a_0) ^ ((fiEnable && (942 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_926_0 <=( _mesh_28_29_io_out_a_0) ^ ((fiEnable && (943 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_927_0 <=( _mesh_28_30_io_out_a_0) ^ ((fiEnable && (944 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_928_0 <=( io_in_a_29_0) ^ ((fiEnable && (945 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_929_0 <=( _mesh_29_0_io_out_a_0) ^ ((fiEnable && (946 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_930_0 <=( _mesh_29_1_io_out_a_0) ^ ((fiEnable && (947 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_931_0 <=( _mesh_29_2_io_out_a_0) ^ ((fiEnable && (948 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_932_0 <=( _mesh_29_3_io_out_a_0) ^ ((fiEnable && (949 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_933_0 <=( _mesh_29_4_io_out_a_0) ^ ((fiEnable && (950 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_934_0 <=( _mesh_29_5_io_out_a_0) ^ ((fiEnable && (951 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_935_0 <=( _mesh_29_6_io_out_a_0) ^ ((fiEnable && (952 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_936_0 <=( _mesh_29_7_io_out_a_0) ^ ((fiEnable && (953 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_937_0 <=( _mesh_29_8_io_out_a_0) ^ ((fiEnable && (954 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_938_0 <=( _mesh_29_9_io_out_a_0) ^ ((fiEnable && (955 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_939_0 <=( _mesh_29_10_io_out_a_0) ^ ((fiEnable && (956 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_940_0 <=( _mesh_29_11_io_out_a_0) ^ ((fiEnable && (957 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_941_0 <=( _mesh_29_12_io_out_a_0) ^ ((fiEnable && (958 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_942_0 <=( _mesh_29_13_io_out_a_0) ^ ((fiEnable && (959 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_943_0 <=( _mesh_29_14_io_out_a_0) ^ ((fiEnable && (960 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_944_0 <=( _mesh_29_15_io_out_a_0) ^ ((fiEnable && (961 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_945_0 <=( _mesh_29_16_io_out_a_0) ^ ((fiEnable && (962 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_946_0 <=( _mesh_29_17_io_out_a_0) ^ ((fiEnable && (963 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_947_0 <=( _mesh_29_18_io_out_a_0) ^ ((fiEnable && (964 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_948_0 <=( _mesh_29_19_io_out_a_0) ^ ((fiEnable && (965 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_949_0 <=( _mesh_29_20_io_out_a_0) ^ ((fiEnable && (966 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_950_0 <=( _mesh_29_21_io_out_a_0) ^ ((fiEnable && (967 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_951_0 <=( _mesh_29_22_io_out_a_0) ^ ((fiEnable && (968 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_952_0 <=( _mesh_29_23_io_out_a_0) ^ ((fiEnable && (969 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_953_0 <=( _mesh_29_24_io_out_a_0) ^ ((fiEnable && (970 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_954_0 <=( _mesh_29_25_io_out_a_0) ^ ((fiEnable && (971 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_955_0 <=( _mesh_29_26_io_out_a_0) ^ ((fiEnable && (972 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_956_0 <=( _mesh_29_27_io_out_a_0) ^ ((fiEnable && (973 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_957_0 <=( _mesh_29_28_io_out_a_0) ^ ((fiEnable && (974 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_958_0 <=( _mesh_29_29_io_out_a_0) ^ ((fiEnable && (975 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_959_0 <=( _mesh_29_30_io_out_a_0) ^ ((fiEnable && (976 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_960_0 <=( io_in_a_30_0) ^ ((fiEnable && (977 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_961_0 <=( _mesh_30_0_io_out_a_0) ^ ((fiEnable && (978 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_962_0 <=( _mesh_30_1_io_out_a_0) ^ ((fiEnable && (979 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_963_0 <=( _mesh_30_2_io_out_a_0) ^ ((fiEnable && (980 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_964_0 <=( _mesh_30_3_io_out_a_0) ^ ((fiEnable && (981 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_965_0 <=( _mesh_30_4_io_out_a_0) ^ ((fiEnable && (982 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_966_0 <=( _mesh_30_5_io_out_a_0) ^ ((fiEnable && (983 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_967_0 <=( _mesh_30_6_io_out_a_0) ^ ((fiEnable && (984 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_968_0 <=( _mesh_30_7_io_out_a_0) ^ ((fiEnable && (985 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_969_0 <=( _mesh_30_8_io_out_a_0) ^ ((fiEnable && (986 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_970_0 <=( _mesh_30_9_io_out_a_0) ^ ((fiEnable && (987 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_971_0 <=( _mesh_30_10_io_out_a_0) ^ ((fiEnable && (988 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_972_0 <=( _mesh_30_11_io_out_a_0) ^ ((fiEnable && (989 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_973_0 <=( _mesh_30_12_io_out_a_0) ^ ((fiEnable && (990 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_974_0 <=( _mesh_30_13_io_out_a_0) ^ ((fiEnable && (991 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_975_0 <=( _mesh_30_14_io_out_a_0) ^ ((fiEnable && (992 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_976_0 <=( _mesh_30_15_io_out_a_0) ^ ((fiEnable && (993 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_977_0 <=( _mesh_30_16_io_out_a_0) ^ ((fiEnable && (994 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_978_0 <=( _mesh_30_17_io_out_a_0) ^ ((fiEnable && (995 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_979_0 <=( _mesh_30_18_io_out_a_0) ^ ((fiEnable && (996 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_980_0 <=( _mesh_30_19_io_out_a_0) ^ ((fiEnable && (997 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_981_0 <=( _mesh_30_20_io_out_a_0) ^ ((fiEnable && (998 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_982_0 <=( _mesh_30_21_io_out_a_0) ^ ((fiEnable && (999 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_983_0 <=( _mesh_30_22_io_out_a_0) ^ ((fiEnable && (1000 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_984_0 <=( _mesh_30_23_io_out_a_0) ^ ((fiEnable && (1001 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_985_0 <=( _mesh_30_24_io_out_a_0) ^ ((fiEnable && (1002 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_986_0 <=( _mesh_30_25_io_out_a_0) ^ ((fiEnable && (1003 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_987_0 <=( _mesh_30_26_io_out_a_0) ^ ((fiEnable && (1004 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_988_0 <=( _mesh_30_27_io_out_a_0) ^ ((fiEnable && (1005 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_989_0 <=( _mesh_30_28_io_out_a_0) ^ ((fiEnable && (1006 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_990_0 <=( _mesh_30_29_io_out_a_0) ^ ((fiEnable && (1007 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_991_0 <=( _mesh_30_30_io_out_a_0) ^ ((fiEnable && (1008 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_992_0 <=( io_in_a_31_0) ^ ((fiEnable && (1009 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_993_0 <=( _mesh_31_0_io_out_a_0) ^ ((fiEnable && (1010 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_994_0 <=( _mesh_31_1_io_out_a_0) ^ ((fiEnable && (1011 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_995_0 <=( _mesh_31_2_io_out_a_0) ^ ((fiEnable && (1012 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_996_0 <=( _mesh_31_3_io_out_a_0) ^ ((fiEnable && (1013 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_997_0 <=( _mesh_31_4_io_out_a_0) ^ ((fiEnable && (1014 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_998_0 <=( _mesh_31_5_io_out_a_0) ^ ((fiEnable && (1015 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_999_0 <=( _mesh_31_6_io_out_a_0) ^ ((fiEnable && (1016 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1000_0 <=( _mesh_31_7_io_out_a_0) ^ ((fiEnable && (1017 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1001_0 <=( _mesh_31_8_io_out_a_0) ^ ((fiEnable && (1018 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1002_0 <=( _mesh_31_9_io_out_a_0) ^ ((fiEnable && (1019 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1003_0 <=( _mesh_31_10_io_out_a_0) ^ ((fiEnable && (1020 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1004_0 <=( _mesh_31_11_io_out_a_0) ^ ((fiEnable && (1021 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1005_0 <=( _mesh_31_12_io_out_a_0) ^ ((fiEnable && (1022 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1006_0 <=( _mesh_31_13_io_out_a_0) ^ ((fiEnable && (1023 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1007_0 <=( _mesh_31_14_io_out_a_0) ^ ((fiEnable && (1024 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1008_0 <=( _mesh_31_15_io_out_a_0) ^ ((fiEnable && (1025 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1009_0 <=( _mesh_31_16_io_out_a_0) ^ ((fiEnable && (1026 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1010_0 <=( _mesh_31_17_io_out_a_0) ^ ((fiEnable && (1027 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1011_0 <=( _mesh_31_18_io_out_a_0) ^ ((fiEnable && (1028 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1012_0 <=( _mesh_31_19_io_out_a_0) ^ ((fiEnable && (1029 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1013_0 <=( _mesh_31_20_io_out_a_0) ^ ((fiEnable && (1030 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1014_0 <=( _mesh_31_21_io_out_a_0) ^ ((fiEnable && (1031 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1015_0 <=( _mesh_31_22_io_out_a_0) ^ ((fiEnable && (1032 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1016_0 <=( _mesh_31_23_io_out_a_0) ^ ((fiEnable && (1033 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1017_0 <=( _mesh_31_24_io_out_a_0) ^ ((fiEnable && (1034 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1018_0 <=( _mesh_31_25_io_out_a_0) ^ ((fiEnable && (1035 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1019_0 <=( _mesh_31_26_io_out_a_0) ^ ((fiEnable && (1036 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1020_0 <=( _mesh_31_27_io_out_a_0) ^ ((fiEnable && (1037 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1021_0 <=( _mesh_31_28_io_out_a_0) ^ ((fiEnable && (1038 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1022_0 <=( _mesh_31_29_io_out_a_0) ^ ((fiEnable && (1039 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1023_0 <=( _mesh_31_30_io_out_a_0) ^ ((fiEnable && (1040 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		if (io_in_valid_0_0) begin
			b_0 <=( io_in_b_0_0) ^ ((fiEnable && (1041 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1024_0 <=( io_in_d_0_0) ^ ((fiEnable && (1042 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_0_io_in_control_0_shift_b <=( io_in_control_0_0_shift) ^ ((fiEnable && (1043 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_0_io_in_control_0_dataflow_b <=( io_in_control_0_0_dataflow) ^ ((fiEnable && (1044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_0_io_in_control_0_propagate_b <=( io_in_control_0_0_propagate) ^ ((fiEnable && (1045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_0_io_out_valid_0) begin
			b_1_0 <=( _mesh_0_0_io_out_b_0) ^ ((fiEnable && (1046 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1025_0 <=( _mesh_0_0_io_out_c_0) ^ ((fiEnable && (1047 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_0_io_in_control_0_shift_b <=( _mesh_0_0_io_out_control_0_shift) ^ ((fiEnable && (1048 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_0_io_in_control_0_dataflow_b <=( _mesh_0_0_io_out_control_0_dataflow) ^ ((fiEnable && (1049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_0_io_in_control_0_propagate_b <=( _mesh_0_0_io_out_control_0_propagate) ^ ((fiEnable && (1050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_0_io_out_valid_0) begin
			b_2_0 <=( _mesh_1_0_io_out_b_0) ^ ((fiEnable && (1051 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1026_0 <=( _mesh_1_0_io_out_c_0) ^ ((fiEnable && (1052 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_0_io_in_control_0_shift_b <=( _mesh_1_0_io_out_control_0_shift) ^ ((fiEnable && (1053 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_0_io_in_control_0_dataflow_b <=( _mesh_1_0_io_out_control_0_dataflow) ^ ((fiEnable && (1054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_0_io_in_control_0_propagate_b <=( _mesh_1_0_io_out_control_0_propagate) ^ ((fiEnable && (1055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_0_io_out_valid_0) begin
			b_3_0 <=( _mesh_2_0_io_out_b_0) ^ ((fiEnable && (1056 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1027_0 <=( _mesh_2_0_io_out_c_0) ^ ((fiEnable && (1057 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_0_io_in_control_0_shift_b <=( _mesh_2_0_io_out_control_0_shift) ^ ((fiEnable && (1058 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_0_io_in_control_0_dataflow_b <=( _mesh_2_0_io_out_control_0_dataflow) ^ ((fiEnable && (1059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_0_io_in_control_0_propagate_b <=( _mesh_2_0_io_out_control_0_propagate) ^ ((fiEnable && (1060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_0_io_out_valid_0) begin
			b_4_0 <=( _mesh_3_0_io_out_b_0) ^ ((fiEnable && (1061 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1028_0 <=( _mesh_3_0_io_out_c_0) ^ ((fiEnable && (1062 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_0_io_in_control_0_shift_b <=( _mesh_3_0_io_out_control_0_shift) ^ ((fiEnable && (1063 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_0_io_in_control_0_dataflow_b <=( _mesh_3_0_io_out_control_0_dataflow) ^ ((fiEnable && (1064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_0_io_in_control_0_propagate_b <=( _mesh_3_0_io_out_control_0_propagate) ^ ((fiEnable && (1065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_0_io_out_valid_0) begin
			b_5_0 <=( _mesh_4_0_io_out_b_0) ^ ((fiEnable && (1066 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1029_0 <=( _mesh_4_0_io_out_c_0) ^ ((fiEnable && (1067 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_0_io_in_control_0_shift_b <=( _mesh_4_0_io_out_control_0_shift) ^ ((fiEnable && (1068 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_0_io_in_control_0_dataflow_b <=( _mesh_4_0_io_out_control_0_dataflow) ^ ((fiEnable && (1069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_0_io_in_control_0_propagate_b <=( _mesh_4_0_io_out_control_0_propagate) ^ ((fiEnable && (1070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_0_io_out_valid_0) begin
			b_6_0 <=( _mesh_5_0_io_out_b_0) ^ ((fiEnable && (1071 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1030_0 <=( _mesh_5_0_io_out_c_0) ^ ((fiEnable && (1072 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_0_io_in_control_0_shift_b <=( _mesh_5_0_io_out_control_0_shift) ^ ((fiEnable && (1073 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_0_io_in_control_0_dataflow_b <=( _mesh_5_0_io_out_control_0_dataflow) ^ ((fiEnable && (1074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_0_io_in_control_0_propagate_b <=( _mesh_5_0_io_out_control_0_propagate) ^ ((fiEnable && (1075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_0_io_out_valid_0) begin
			b_7_0 <=( _mesh_6_0_io_out_b_0) ^ ((fiEnable && (1076 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1031_0 <=( _mesh_6_0_io_out_c_0) ^ ((fiEnable && (1077 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_0_io_in_control_0_shift_b <=( _mesh_6_0_io_out_control_0_shift) ^ ((fiEnable && (1078 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_0_io_in_control_0_dataflow_b <=( _mesh_6_0_io_out_control_0_dataflow) ^ ((fiEnable && (1079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_0_io_in_control_0_propagate_b <=( _mesh_6_0_io_out_control_0_propagate) ^ ((fiEnable && (1080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_0_io_out_valid_0) begin
			b_8_0 <=( _mesh_7_0_io_out_b_0) ^ ((fiEnable && (1081 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1032_0 <=( _mesh_7_0_io_out_c_0) ^ ((fiEnable && (1082 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_0_io_in_control_0_shift_b <=( _mesh_7_0_io_out_control_0_shift) ^ ((fiEnable && (1083 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_0_io_in_control_0_dataflow_b <=( _mesh_7_0_io_out_control_0_dataflow) ^ ((fiEnable && (1084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_0_io_in_control_0_propagate_b <=( _mesh_7_0_io_out_control_0_propagate) ^ ((fiEnable && (1085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_0_io_out_valid_0) begin
			b_9_0 <=( _mesh_8_0_io_out_b_0) ^ ((fiEnable && (1086 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1033_0 <=( _mesh_8_0_io_out_c_0) ^ ((fiEnable && (1087 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_0_io_in_control_0_shift_b <=( _mesh_8_0_io_out_control_0_shift) ^ ((fiEnable && (1088 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_0_io_in_control_0_dataflow_b <=( _mesh_8_0_io_out_control_0_dataflow) ^ ((fiEnable && (1089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_0_io_in_control_0_propagate_b <=( _mesh_8_0_io_out_control_0_propagate) ^ ((fiEnable && (1090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_0_io_out_valid_0) begin
			b_10_0 <=( _mesh_9_0_io_out_b_0) ^ ((fiEnable && (1091 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1034_0 <=( _mesh_9_0_io_out_c_0) ^ ((fiEnable && (1092 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_0_io_in_control_0_shift_b <=( _mesh_9_0_io_out_control_0_shift) ^ ((fiEnable && (1093 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_0_io_in_control_0_dataflow_b <=( _mesh_9_0_io_out_control_0_dataflow) ^ ((fiEnable && (1094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_0_io_in_control_0_propagate_b <=( _mesh_9_0_io_out_control_0_propagate) ^ ((fiEnable && (1095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_0_io_out_valid_0) begin
			b_11_0 <=( _mesh_10_0_io_out_b_0) ^ ((fiEnable && (1096 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1035_0 <=( _mesh_10_0_io_out_c_0) ^ ((fiEnable && (1097 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_0_io_in_control_0_shift_b <=( _mesh_10_0_io_out_control_0_shift) ^ ((fiEnable && (1098 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_0_io_in_control_0_dataflow_b <=( _mesh_10_0_io_out_control_0_dataflow) ^ ((fiEnable && (1099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_0_io_in_control_0_propagate_b <=( _mesh_10_0_io_out_control_0_propagate) ^ ((fiEnable && (1100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_0_io_out_valid_0) begin
			b_12_0 <=( _mesh_11_0_io_out_b_0) ^ ((fiEnable && (1101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1036_0 <=( _mesh_11_0_io_out_c_0) ^ ((fiEnable && (1102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_0_io_in_control_0_shift_b <=( _mesh_11_0_io_out_control_0_shift) ^ ((fiEnable && (1103 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_0_io_in_control_0_dataflow_b <=( _mesh_11_0_io_out_control_0_dataflow) ^ ((fiEnable && (1104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_0_io_in_control_0_propagate_b <=( _mesh_11_0_io_out_control_0_propagate) ^ ((fiEnable && (1105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_0_io_out_valid_0) begin
			b_13_0 <=( _mesh_12_0_io_out_b_0) ^ ((fiEnable && (1106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1037_0 <=( _mesh_12_0_io_out_c_0) ^ ((fiEnable && (1107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_0_io_in_control_0_shift_b <=( _mesh_12_0_io_out_control_0_shift) ^ ((fiEnable && (1108 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_0_io_in_control_0_dataflow_b <=( _mesh_12_0_io_out_control_0_dataflow) ^ ((fiEnable && (1109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_0_io_in_control_0_propagate_b <=( _mesh_12_0_io_out_control_0_propagate) ^ ((fiEnable && (1110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_0_io_out_valid_0) begin
			b_14_0 <=( _mesh_13_0_io_out_b_0) ^ ((fiEnable && (1111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1038_0 <=( _mesh_13_0_io_out_c_0) ^ ((fiEnable && (1112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_0_io_in_control_0_shift_b <=( _mesh_13_0_io_out_control_0_shift) ^ ((fiEnable && (1113 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_0_io_in_control_0_dataflow_b <=( _mesh_13_0_io_out_control_0_dataflow) ^ ((fiEnable && (1114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_0_io_in_control_0_propagate_b <=( _mesh_13_0_io_out_control_0_propagate) ^ ((fiEnable && (1115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_0_io_out_valid_0) begin
			b_15_0 <=( _mesh_14_0_io_out_b_0) ^ ((fiEnable && (1116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1039_0 <=( _mesh_14_0_io_out_c_0) ^ ((fiEnable && (1117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_0_io_in_control_0_shift_b <=( _mesh_14_0_io_out_control_0_shift) ^ ((fiEnable && (1118 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_0_io_in_control_0_dataflow_b <=( _mesh_14_0_io_out_control_0_dataflow) ^ ((fiEnable && (1119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_0_io_in_control_0_propagate_b <=( _mesh_14_0_io_out_control_0_propagate) ^ ((fiEnable && (1120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_0_io_out_valid_0) begin
			b_16_0 <=( _mesh_15_0_io_out_b_0) ^ ((fiEnable && (1121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1040_0 <=( _mesh_15_0_io_out_c_0) ^ ((fiEnable && (1122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_0_io_in_control_0_shift_b <=( _mesh_15_0_io_out_control_0_shift) ^ ((fiEnable && (1123 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_0_io_in_control_0_dataflow_b <=( _mesh_15_0_io_out_control_0_dataflow) ^ ((fiEnable && (1124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_0_io_in_control_0_propagate_b <=( _mesh_15_0_io_out_control_0_propagate) ^ ((fiEnable && (1125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_0_io_out_valid_0) begin
			b_17_0 <=( _mesh_16_0_io_out_b_0) ^ ((fiEnable && (1126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1041_0 <=( _mesh_16_0_io_out_c_0) ^ ((fiEnable && (1127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_0_io_in_control_0_shift_b <=( _mesh_16_0_io_out_control_0_shift) ^ ((fiEnable && (1128 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_0_io_in_control_0_dataflow_b <=( _mesh_16_0_io_out_control_0_dataflow) ^ ((fiEnable && (1129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_0_io_in_control_0_propagate_b <=( _mesh_16_0_io_out_control_0_propagate) ^ ((fiEnable && (1130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_0_io_out_valid_0) begin
			b_18_0 <=( _mesh_17_0_io_out_b_0) ^ ((fiEnable && (1131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1042_0 <=( _mesh_17_0_io_out_c_0) ^ ((fiEnable && (1132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_0_io_in_control_0_shift_b <=( _mesh_17_0_io_out_control_0_shift) ^ ((fiEnable && (1133 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_0_io_in_control_0_dataflow_b <=( _mesh_17_0_io_out_control_0_dataflow) ^ ((fiEnable && (1134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_0_io_in_control_0_propagate_b <=( _mesh_17_0_io_out_control_0_propagate) ^ ((fiEnable && (1135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_0_io_out_valid_0) begin
			b_19_0 <=( _mesh_18_0_io_out_b_0) ^ ((fiEnable && (1136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1043_0 <=( _mesh_18_0_io_out_c_0) ^ ((fiEnable && (1137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_0_io_in_control_0_shift_b <=( _mesh_18_0_io_out_control_0_shift) ^ ((fiEnable && (1138 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_0_io_in_control_0_dataflow_b <=( _mesh_18_0_io_out_control_0_dataflow) ^ ((fiEnable && (1139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_0_io_in_control_0_propagate_b <=( _mesh_18_0_io_out_control_0_propagate) ^ ((fiEnable && (1140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_0_io_out_valid_0) begin
			b_20_0 <=( _mesh_19_0_io_out_b_0) ^ ((fiEnable && (1141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1044_0 <=( _mesh_19_0_io_out_c_0) ^ ((fiEnable && (1142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_0_io_in_control_0_shift_b <=( _mesh_19_0_io_out_control_0_shift) ^ ((fiEnable && (1143 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_0_io_in_control_0_dataflow_b <=( _mesh_19_0_io_out_control_0_dataflow) ^ ((fiEnable && (1144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_0_io_in_control_0_propagate_b <=( _mesh_19_0_io_out_control_0_propagate) ^ ((fiEnable && (1145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_0_io_out_valid_0) begin
			b_21_0 <=( _mesh_20_0_io_out_b_0) ^ ((fiEnable && (1146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1045_0 <=( _mesh_20_0_io_out_c_0) ^ ((fiEnable && (1147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_0_io_in_control_0_shift_b <=( _mesh_20_0_io_out_control_0_shift) ^ ((fiEnable && (1148 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_0_io_in_control_0_dataflow_b <=( _mesh_20_0_io_out_control_0_dataflow) ^ ((fiEnable && (1149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_0_io_in_control_0_propagate_b <=( _mesh_20_0_io_out_control_0_propagate) ^ ((fiEnable && (1150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_0_io_out_valid_0) begin
			b_22_0 <=( _mesh_21_0_io_out_b_0) ^ ((fiEnable && (1151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1046_0 <=( _mesh_21_0_io_out_c_0) ^ ((fiEnable && (1152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_0_io_in_control_0_shift_b <=( _mesh_21_0_io_out_control_0_shift) ^ ((fiEnable && (1153 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_0_io_in_control_0_dataflow_b <=( _mesh_21_0_io_out_control_0_dataflow) ^ ((fiEnable && (1154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_0_io_in_control_0_propagate_b <=( _mesh_21_0_io_out_control_0_propagate) ^ ((fiEnable && (1155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_0_io_out_valid_0) begin
			b_23_0 <=( _mesh_22_0_io_out_b_0) ^ ((fiEnable && (1156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1047_0 <=( _mesh_22_0_io_out_c_0) ^ ((fiEnable && (1157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_0_io_in_control_0_shift_b <=( _mesh_22_0_io_out_control_0_shift) ^ ((fiEnable && (1158 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_0_io_in_control_0_dataflow_b <=( _mesh_22_0_io_out_control_0_dataflow) ^ ((fiEnable && (1159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_0_io_in_control_0_propagate_b <=( _mesh_22_0_io_out_control_0_propagate) ^ ((fiEnable && (1160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_0_io_out_valid_0) begin
			b_24_0 <=( _mesh_23_0_io_out_b_0) ^ ((fiEnable && (1161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1048_0 <=( _mesh_23_0_io_out_c_0) ^ ((fiEnable && (1162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_0_io_in_control_0_shift_b <=( _mesh_23_0_io_out_control_0_shift) ^ ((fiEnable && (1163 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_0_io_in_control_0_dataflow_b <=( _mesh_23_0_io_out_control_0_dataflow) ^ ((fiEnable && (1164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_0_io_in_control_0_propagate_b <=( _mesh_23_0_io_out_control_0_propagate) ^ ((fiEnable && (1165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_0_io_out_valid_0) begin
			b_25_0 <=( _mesh_24_0_io_out_b_0) ^ ((fiEnable && (1166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1049_0 <=( _mesh_24_0_io_out_c_0) ^ ((fiEnable && (1167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_0_io_in_control_0_shift_b <=( _mesh_24_0_io_out_control_0_shift) ^ ((fiEnable && (1168 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_0_io_in_control_0_dataflow_b <=( _mesh_24_0_io_out_control_0_dataflow) ^ ((fiEnable && (1169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_0_io_in_control_0_propagate_b <=( _mesh_24_0_io_out_control_0_propagate) ^ ((fiEnable && (1170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_0_io_out_valid_0) begin
			b_26_0 <=( _mesh_25_0_io_out_b_0) ^ ((fiEnable && (1171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1050_0 <=( _mesh_25_0_io_out_c_0) ^ ((fiEnable && (1172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_0_io_in_control_0_shift_b <=( _mesh_25_0_io_out_control_0_shift) ^ ((fiEnable && (1173 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_0_io_in_control_0_dataflow_b <=( _mesh_25_0_io_out_control_0_dataflow) ^ ((fiEnable && (1174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_0_io_in_control_0_propagate_b <=( _mesh_25_0_io_out_control_0_propagate) ^ ((fiEnable && (1175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_0_io_out_valid_0) begin
			b_27_0 <=( _mesh_26_0_io_out_b_0) ^ ((fiEnable && (1176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1051_0 <=( _mesh_26_0_io_out_c_0) ^ ((fiEnable && (1177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_0_io_in_control_0_shift_b <=( _mesh_26_0_io_out_control_0_shift) ^ ((fiEnable && (1178 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_0_io_in_control_0_dataflow_b <=( _mesh_26_0_io_out_control_0_dataflow) ^ ((fiEnable && (1179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_0_io_in_control_0_propagate_b <=( _mesh_26_0_io_out_control_0_propagate) ^ ((fiEnable && (1180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_0_io_out_valid_0) begin
			b_28_0 <=( _mesh_27_0_io_out_b_0) ^ ((fiEnable && (1181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1052_0 <=( _mesh_27_0_io_out_c_0) ^ ((fiEnable && (1182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_0_io_in_control_0_shift_b <=( _mesh_27_0_io_out_control_0_shift) ^ ((fiEnable && (1183 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_0_io_in_control_0_dataflow_b <=( _mesh_27_0_io_out_control_0_dataflow) ^ ((fiEnable && (1184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_0_io_in_control_0_propagate_b <=( _mesh_27_0_io_out_control_0_propagate) ^ ((fiEnable && (1185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_0_io_out_valid_0) begin
			b_29_0 <=( _mesh_28_0_io_out_b_0) ^ ((fiEnable && (1186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1053_0 <=( _mesh_28_0_io_out_c_0) ^ ((fiEnable && (1187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_0_io_in_control_0_shift_b <=( _mesh_28_0_io_out_control_0_shift) ^ ((fiEnable && (1188 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_0_io_in_control_0_dataflow_b <=( _mesh_28_0_io_out_control_0_dataflow) ^ ((fiEnable && (1189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_0_io_in_control_0_propagate_b <=( _mesh_28_0_io_out_control_0_propagate) ^ ((fiEnable && (1190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_0_io_out_valid_0) begin
			b_30_0 <=( _mesh_29_0_io_out_b_0) ^ ((fiEnable && (1191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1054_0 <=( _mesh_29_0_io_out_c_0) ^ ((fiEnable && (1192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_0_io_in_control_0_shift_b <=( _mesh_29_0_io_out_control_0_shift) ^ ((fiEnable && (1193 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_0_io_in_control_0_dataflow_b <=( _mesh_29_0_io_out_control_0_dataflow) ^ ((fiEnable && (1194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_0_io_in_control_0_propagate_b <=( _mesh_29_0_io_out_control_0_propagate) ^ ((fiEnable && (1195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_0_io_out_valid_0) begin
			b_31_0 <=( _mesh_30_0_io_out_b_0) ^ ((fiEnable && (1196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1055_0 <=( _mesh_30_0_io_out_c_0) ^ ((fiEnable && (1197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_0_io_in_control_0_shift_b <=( _mesh_30_0_io_out_control_0_shift) ^ ((fiEnable && (1198 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_0_io_in_control_0_dataflow_b <=( _mesh_30_0_io_out_control_0_dataflow) ^ ((fiEnable && (1199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_0_io_in_control_0_propagate_b <=( _mesh_30_0_io_out_control_0_propagate) ^ ((fiEnable && (1200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_1_0) begin
			b_32_0 <=( io_in_b_1_0) ^ ((fiEnable && (1201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1056_0 <=( io_in_d_1_0) ^ ((fiEnable && (1202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_1_io_in_control_0_shift_b <=( io_in_control_1_0_shift) ^ ((fiEnable && (1203 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_1_io_in_control_0_dataflow_b <=( io_in_control_1_0_dataflow) ^ ((fiEnable && (1204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_1_io_in_control_0_propagate_b <=( io_in_control_1_0_propagate) ^ ((fiEnable && (1205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_1_io_out_valid_0) begin
			b_33_0 <=( _mesh_0_1_io_out_b_0) ^ ((fiEnable && (1206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1057_0 <=( _mesh_0_1_io_out_c_0) ^ ((fiEnable && (1207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_1_io_in_control_0_shift_b <=( _mesh_0_1_io_out_control_0_shift) ^ ((fiEnable && (1208 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_1_io_in_control_0_dataflow_b <=( _mesh_0_1_io_out_control_0_dataflow) ^ ((fiEnable && (1209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_1_io_in_control_0_propagate_b <=( _mesh_0_1_io_out_control_0_propagate) ^ ((fiEnable && (1210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_1_io_out_valid_0) begin
			b_34_0 <=( _mesh_1_1_io_out_b_0) ^ ((fiEnable && (1211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1058_0 <=( _mesh_1_1_io_out_c_0) ^ ((fiEnable && (1212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_1_io_in_control_0_shift_b <=( _mesh_1_1_io_out_control_0_shift) ^ ((fiEnable && (1213 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_1_io_in_control_0_dataflow_b <=( _mesh_1_1_io_out_control_0_dataflow) ^ ((fiEnable && (1214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_1_io_in_control_0_propagate_b <=( _mesh_1_1_io_out_control_0_propagate) ^ ((fiEnable && (1215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_1_io_out_valid_0) begin
			b_35_0 <=( _mesh_2_1_io_out_b_0) ^ ((fiEnable && (1216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1059_0 <=( _mesh_2_1_io_out_c_0) ^ ((fiEnable && (1217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_1_io_in_control_0_shift_b <=( _mesh_2_1_io_out_control_0_shift) ^ ((fiEnable && (1218 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_1_io_in_control_0_dataflow_b <=( _mesh_2_1_io_out_control_0_dataflow) ^ ((fiEnable && (1219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_1_io_in_control_0_propagate_b <=( _mesh_2_1_io_out_control_0_propagate) ^ ((fiEnable && (1220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_1_io_out_valid_0) begin
			b_36_0 <=( _mesh_3_1_io_out_b_0) ^ ((fiEnable && (1221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1060_0 <=( _mesh_3_1_io_out_c_0) ^ ((fiEnable && (1222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_1_io_in_control_0_shift_b <=( _mesh_3_1_io_out_control_0_shift) ^ ((fiEnable && (1223 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_1_io_in_control_0_dataflow_b <=( _mesh_3_1_io_out_control_0_dataflow) ^ ((fiEnable && (1224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_1_io_in_control_0_propagate_b <=( _mesh_3_1_io_out_control_0_propagate) ^ ((fiEnable && (1225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_1_io_out_valid_0) begin
			b_37_0 <=( _mesh_4_1_io_out_b_0) ^ ((fiEnable && (1226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1061_0 <=( _mesh_4_1_io_out_c_0) ^ ((fiEnable && (1227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_1_io_in_control_0_shift_b <=( _mesh_4_1_io_out_control_0_shift) ^ ((fiEnable && (1228 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_1_io_in_control_0_dataflow_b <=( _mesh_4_1_io_out_control_0_dataflow) ^ ((fiEnable && (1229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_1_io_in_control_0_propagate_b <=( _mesh_4_1_io_out_control_0_propagate) ^ ((fiEnable && (1230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_1_io_out_valid_0) begin
			b_38_0 <=( _mesh_5_1_io_out_b_0) ^ ((fiEnable && (1231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1062_0 <=( _mesh_5_1_io_out_c_0) ^ ((fiEnable && (1232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_1_io_in_control_0_shift_b <=( _mesh_5_1_io_out_control_0_shift) ^ ((fiEnable && (1233 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_1_io_in_control_0_dataflow_b <=( _mesh_5_1_io_out_control_0_dataflow) ^ ((fiEnable && (1234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_1_io_in_control_0_propagate_b <=( _mesh_5_1_io_out_control_0_propagate) ^ ((fiEnable && (1235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_1_io_out_valid_0) begin
			b_39_0 <=( _mesh_6_1_io_out_b_0) ^ ((fiEnable && (1236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1063_0 <=( _mesh_6_1_io_out_c_0) ^ ((fiEnable && (1237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_1_io_in_control_0_shift_b <=( _mesh_6_1_io_out_control_0_shift) ^ ((fiEnable && (1238 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_1_io_in_control_0_dataflow_b <=( _mesh_6_1_io_out_control_0_dataflow) ^ ((fiEnable && (1239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_1_io_in_control_0_propagate_b <=( _mesh_6_1_io_out_control_0_propagate) ^ ((fiEnable && (1240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_1_io_out_valid_0) begin
			b_40_0 <=( _mesh_7_1_io_out_b_0) ^ ((fiEnable && (1241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1064_0 <=( _mesh_7_1_io_out_c_0) ^ ((fiEnable && (1242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_1_io_in_control_0_shift_b <=( _mesh_7_1_io_out_control_0_shift) ^ ((fiEnable && (1243 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_1_io_in_control_0_dataflow_b <=( _mesh_7_1_io_out_control_0_dataflow) ^ ((fiEnable && (1244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_1_io_in_control_0_propagate_b <=( _mesh_7_1_io_out_control_0_propagate) ^ ((fiEnable && (1245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_1_io_out_valid_0) begin
			b_41_0 <=( _mesh_8_1_io_out_b_0) ^ ((fiEnable && (1246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1065_0 <=( _mesh_8_1_io_out_c_0) ^ ((fiEnable && (1247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_1_io_in_control_0_shift_b <=( _mesh_8_1_io_out_control_0_shift) ^ ((fiEnable && (1248 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_1_io_in_control_0_dataflow_b <=( _mesh_8_1_io_out_control_0_dataflow) ^ ((fiEnable && (1249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_1_io_in_control_0_propagate_b <=( _mesh_8_1_io_out_control_0_propagate) ^ ((fiEnable && (1250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_1_io_out_valid_0) begin
			b_42_0 <=( _mesh_9_1_io_out_b_0) ^ ((fiEnable && (1251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1066_0 <=( _mesh_9_1_io_out_c_0) ^ ((fiEnable && (1252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_1_io_in_control_0_shift_b <=( _mesh_9_1_io_out_control_0_shift) ^ ((fiEnable && (1253 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_1_io_in_control_0_dataflow_b <=( _mesh_9_1_io_out_control_0_dataflow) ^ ((fiEnable && (1254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_1_io_in_control_0_propagate_b <=( _mesh_9_1_io_out_control_0_propagate) ^ ((fiEnable && (1255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_1_io_out_valid_0) begin
			b_43_0 <=( _mesh_10_1_io_out_b_0) ^ ((fiEnable && (1256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1067_0 <=( _mesh_10_1_io_out_c_0) ^ ((fiEnable && (1257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_1_io_in_control_0_shift_b <=( _mesh_10_1_io_out_control_0_shift) ^ ((fiEnable && (1258 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_1_io_in_control_0_dataflow_b <=( _mesh_10_1_io_out_control_0_dataflow) ^ ((fiEnable && (1259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_1_io_in_control_0_propagate_b <=( _mesh_10_1_io_out_control_0_propagate) ^ ((fiEnable && (1260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_1_io_out_valid_0) begin
			b_44_0 <=( _mesh_11_1_io_out_b_0) ^ ((fiEnable && (1261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1068_0 <=( _mesh_11_1_io_out_c_0) ^ ((fiEnable && (1262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_1_io_in_control_0_shift_b <=( _mesh_11_1_io_out_control_0_shift) ^ ((fiEnable && (1263 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_1_io_in_control_0_dataflow_b <=( _mesh_11_1_io_out_control_0_dataflow) ^ ((fiEnable && (1264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_1_io_in_control_0_propagate_b <=( _mesh_11_1_io_out_control_0_propagate) ^ ((fiEnable && (1265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_1_io_out_valid_0) begin
			b_45_0 <=( _mesh_12_1_io_out_b_0) ^ ((fiEnable && (1266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1069_0 <=( _mesh_12_1_io_out_c_0) ^ ((fiEnable && (1267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_1_io_in_control_0_shift_b <=( _mesh_12_1_io_out_control_0_shift) ^ ((fiEnable && (1268 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_1_io_in_control_0_dataflow_b <=( _mesh_12_1_io_out_control_0_dataflow) ^ ((fiEnable && (1269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_1_io_in_control_0_propagate_b <=( _mesh_12_1_io_out_control_0_propagate) ^ ((fiEnable && (1270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_1_io_out_valid_0) begin
			b_46_0 <=( _mesh_13_1_io_out_b_0) ^ ((fiEnable && (1271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1070_0 <=( _mesh_13_1_io_out_c_0) ^ ((fiEnable && (1272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_1_io_in_control_0_shift_b <=( _mesh_13_1_io_out_control_0_shift) ^ ((fiEnable && (1273 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_1_io_in_control_0_dataflow_b <=( _mesh_13_1_io_out_control_0_dataflow) ^ ((fiEnable && (1274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_1_io_in_control_0_propagate_b <=( _mesh_13_1_io_out_control_0_propagate) ^ ((fiEnable && (1275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_1_io_out_valid_0) begin
			b_47_0 <=( _mesh_14_1_io_out_b_0) ^ ((fiEnable && (1276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1071_0 <=( _mesh_14_1_io_out_c_0) ^ ((fiEnable && (1277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_1_io_in_control_0_shift_b <=( _mesh_14_1_io_out_control_0_shift) ^ ((fiEnable && (1278 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_1_io_in_control_0_dataflow_b <=( _mesh_14_1_io_out_control_0_dataflow) ^ ((fiEnable && (1279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_1_io_in_control_0_propagate_b <=( _mesh_14_1_io_out_control_0_propagate) ^ ((fiEnable && (1280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_1_io_out_valid_0) begin
			b_48_0 <=( _mesh_15_1_io_out_b_0) ^ ((fiEnable && (1281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1072_0 <=( _mesh_15_1_io_out_c_0) ^ ((fiEnable && (1282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_1_io_in_control_0_shift_b <=( _mesh_15_1_io_out_control_0_shift) ^ ((fiEnable && (1283 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_1_io_in_control_0_dataflow_b <=( _mesh_15_1_io_out_control_0_dataflow) ^ ((fiEnable && (1284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_1_io_in_control_0_propagate_b <=( _mesh_15_1_io_out_control_0_propagate) ^ ((fiEnable && (1285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_1_io_out_valid_0) begin
			b_49_0 <=( _mesh_16_1_io_out_b_0) ^ ((fiEnable && (1286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1073_0 <=( _mesh_16_1_io_out_c_0) ^ ((fiEnable && (1287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_1_io_in_control_0_shift_b <=( _mesh_16_1_io_out_control_0_shift) ^ ((fiEnable && (1288 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_1_io_in_control_0_dataflow_b <=( _mesh_16_1_io_out_control_0_dataflow) ^ ((fiEnable && (1289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_1_io_in_control_0_propagate_b <=( _mesh_16_1_io_out_control_0_propagate) ^ ((fiEnable && (1290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_1_io_out_valid_0) begin
			b_50_0 <=( _mesh_17_1_io_out_b_0) ^ ((fiEnable && (1291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1074_0 <=( _mesh_17_1_io_out_c_0) ^ ((fiEnable && (1292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_1_io_in_control_0_shift_b <=( _mesh_17_1_io_out_control_0_shift) ^ ((fiEnable && (1293 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_1_io_in_control_0_dataflow_b <=( _mesh_17_1_io_out_control_0_dataflow) ^ ((fiEnable && (1294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_1_io_in_control_0_propagate_b <=( _mesh_17_1_io_out_control_0_propagate) ^ ((fiEnable && (1295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_1_io_out_valid_0) begin
			b_51_0 <=( _mesh_18_1_io_out_b_0) ^ ((fiEnable && (1296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1075_0 <=( _mesh_18_1_io_out_c_0) ^ ((fiEnable && (1297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_1_io_in_control_0_shift_b <=( _mesh_18_1_io_out_control_0_shift) ^ ((fiEnable && (1298 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_1_io_in_control_0_dataflow_b <=( _mesh_18_1_io_out_control_0_dataflow) ^ ((fiEnable && (1299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_1_io_in_control_0_propagate_b <=( _mesh_18_1_io_out_control_0_propagate) ^ ((fiEnable && (1300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_1_io_out_valid_0) begin
			b_52_0 <=( _mesh_19_1_io_out_b_0) ^ ((fiEnable && (1301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1076_0 <=( _mesh_19_1_io_out_c_0) ^ ((fiEnable && (1302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_1_io_in_control_0_shift_b <=( _mesh_19_1_io_out_control_0_shift) ^ ((fiEnable && (1303 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_1_io_in_control_0_dataflow_b <=( _mesh_19_1_io_out_control_0_dataflow) ^ ((fiEnable && (1304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_1_io_in_control_0_propagate_b <=( _mesh_19_1_io_out_control_0_propagate) ^ ((fiEnable && (1305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_1_io_out_valid_0) begin
			b_53_0 <=( _mesh_20_1_io_out_b_0) ^ ((fiEnable && (1306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1077_0 <=( _mesh_20_1_io_out_c_0) ^ ((fiEnable && (1307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_1_io_in_control_0_shift_b <=( _mesh_20_1_io_out_control_0_shift) ^ ((fiEnable && (1308 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_1_io_in_control_0_dataflow_b <=( _mesh_20_1_io_out_control_0_dataflow) ^ ((fiEnable && (1309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_1_io_in_control_0_propagate_b <=( _mesh_20_1_io_out_control_0_propagate) ^ ((fiEnable && (1310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_1_io_out_valid_0) begin
			b_54_0 <=( _mesh_21_1_io_out_b_0) ^ ((fiEnable && (1311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1078_0 <=( _mesh_21_1_io_out_c_0) ^ ((fiEnable && (1312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_1_io_in_control_0_shift_b <=( _mesh_21_1_io_out_control_0_shift) ^ ((fiEnable && (1313 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_1_io_in_control_0_dataflow_b <=( _mesh_21_1_io_out_control_0_dataflow) ^ ((fiEnable && (1314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_1_io_in_control_0_propagate_b <=( _mesh_21_1_io_out_control_0_propagate) ^ ((fiEnable && (1315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_1_io_out_valid_0) begin
			b_55_0 <=( _mesh_22_1_io_out_b_0) ^ ((fiEnable && (1316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1079_0 <=( _mesh_22_1_io_out_c_0) ^ ((fiEnable && (1317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_1_io_in_control_0_shift_b <=( _mesh_22_1_io_out_control_0_shift) ^ ((fiEnable && (1318 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_1_io_in_control_0_dataflow_b <=( _mesh_22_1_io_out_control_0_dataflow) ^ ((fiEnable && (1319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_1_io_in_control_0_propagate_b <=( _mesh_22_1_io_out_control_0_propagate) ^ ((fiEnable && (1320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_1_io_out_valid_0) begin
			b_56_0 <=( _mesh_23_1_io_out_b_0) ^ ((fiEnable && (1321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1080_0 <=( _mesh_23_1_io_out_c_0) ^ ((fiEnable && (1322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_1_io_in_control_0_shift_b <=( _mesh_23_1_io_out_control_0_shift) ^ ((fiEnable && (1323 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_1_io_in_control_0_dataflow_b <=( _mesh_23_1_io_out_control_0_dataflow) ^ ((fiEnable && (1324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_1_io_in_control_0_propagate_b <=( _mesh_23_1_io_out_control_0_propagate) ^ ((fiEnable && (1325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_1_io_out_valid_0) begin
			b_57_0 <=( _mesh_24_1_io_out_b_0) ^ ((fiEnable && (1326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1081_0 <=( _mesh_24_1_io_out_c_0) ^ ((fiEnable && (1327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_1_io_in_control_0_shift_b <=( _mesh_24_1_io_out_control_0_shift) ^ ((fiEnable && (1328 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_1_io_in_control_0_dataflow_b <=( _mesh_24_1_io_out_control_0_dataflow) ^ ((fiEnable && (1329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_1_io_in_control_0_propagate_b <=( _mesh_24_1_io_out_control_0_propagate) ^ ((fiEnable && (1330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_1_io_out_valid_0) begin
			b_58_0 <=( _mesh_25_1_io_out_b_0) ^ ((fiEnable && (1331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1082_0 <=( _mesh_25_1_io_out_c_0) ^ ((fiEnable && (1332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_1_io_in_control_0_shift_b <=( _mesh_25_1_io_out_control_0_shift) ^ ((fiEnable && (1333 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_1_io_in_control_0_dataflow_b <=( _mesh_25_1_io_out_control_0_dataflow) ^ ((fiEnable && (1334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_1_io_in_control_0_propagate_b <=( _mesh_25_1_io_out_control_0_propagate) ^ ((fiEnable && (1335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_1_io_out_valid_0) begin
			b_59_0 <=( _mesh_26_1_io_out_b_0) ^ ((fiEnable && (1336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1083_0 <=( _mesh_26_1_io_out_c_0) ^ ((fiEnable && (1337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_1_io_in_control_0_shift_b <=( _mesh_26_1_io_out_control_0_shift) ^ ((fiEnable && (1338 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_1_io_in_control_0_dataflow_b <=( _mesh_26_1_io_out_control_0_dataflow) ^ ((fiEnable && (1339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_1_io_in_control_0_propagate_b <=( _mesh_26_1_io_out_control_0_propagate) ^ ((fiEnable && (1340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_1_io_out_valid_0) begin
			b_60_0 <=( _mesh_27_1_io_out_b_0) ^ ((fiEnable && (1341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1084_0 <=( _mesh_27_1_io_out_c_0) ^ ((fiEnable && (1342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_1_io_in_control_0_shift_b <=( _mesh_27_1_io_out_control_0_shift) ^ ((fiEnable && (1343 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_1_io_in_control_0_dataflow_b <=( _mesh_27_1_io_out_control_0_dataflow) ^ ((fiEnable && (1344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_1_io_in_control_0_propagate_b <=( _mesh_27_1_io_out_control_0_propagate) ^ ((fiEnable && (1345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_1_io_out_valid_0) begin
			b_61_0 <=( _mesh_28_1_io_out_b_0) ^ ((fiEnable && (1346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1085_0 <=( _mesh_28_1_io_out_c_0) ^ ((fiEnable && (1347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_1_io_in_control_0_shift_b <=( _mesh_28_1_io_out_control_0_shift) ^ ((fiEnable && (1348 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_1_io_in_control_0_dataflow_b <=( _mesh_28_1_io_out_control_0_dataflow) ^ ((fiEnable && (1349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_1_io_in_control_0_propagate_b <=( _mesh_28_1_io_out_control_0_propagate) ^ ((fiEnable && (1350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_1_io_out_valid_0) begin
			b_62_0 <=( _mesh_29_1_io_out_b_0) ^ ((fiEnable && (1351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1086_0 <=( _mesh_29_1_io_out_c_0) ^ ((fiEnable && (1352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_1_io_in_control_0_shift_b <=( _mesh_29_1_io_out_control_0_shift) ^ ((fiEnable && (1353 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_1_io_in_control_0_dataflow_b <=( _mesh_29_1_io_out_control_0_dataflow) ^ ((fiEnable && (1354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_1_io_in_control_0_propagate_b <=( _mesh_29_1_io_out_control_0_propagate) ^ ((fiEnable && (1355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_1_io_out_valid_0) begin
			b_63_0 <=( _mesh_30_1_io_out_b_0) ^ ((fiEnable && (1356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1087_0 <=( _mesh_30_1_io_out_c_0) ^ ((fiEnable && (1357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_1_io_in_control_0_shift_b <=( _mesh_30_1_io_out_control_0_shift) ^ ((fiEnable && (1358 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_1_io_in_control_0_dataflow_b <=( _mesh_30_1_io_out_control_0_dataflow) ^ ((fiEnable && (1359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_1_io_in_control_0_propagate_b <=( _mesh_30_1_io_out_control_0_propagate) ^ ((fiEnable && (1360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_2_0) begin
			b_64_0 <=( io_in_b_2_0) ^ ((fiEnable && (1361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1088_0 <=( io_in_d_2_0) ^ ((fiEnable && (1362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_2_io_in_control_0_shift_b <=( io_in_control_2_0_shift) ^ ((fiEnable && (1363 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_2_io_in_control_0_dataflow_b <=( io_in_control_2_0_dataflow) ^ ((fiEnable && (1364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_2_io_in_control_0_propagate_b <=( io_in_control_2_0_propagate) ^ ((fiEnable && (1365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_2_io_out_valid_0) begin
			b_65_0 <=( _mesh_0_2_io_out_b_0) ^ ((fiEnable && (1366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1089_0 <=( _mesh_0_2_io_out_c_0) ^ ((fiEnable && (1367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_2_io_in_control_0_shift_b <=( _mesh_0_2_io_out_control_0_shift) ^ ((fiEnable && (1368 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_2_io_in_control_0_dataflow_b <=( _mesh_0_2_io_out_control_0_dataflow) ^ ((fiEnable && (1369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_2_io_in_control_0_propagate_b <=( _mesh_0_2_io_out_control_0_propagate) ^ ((fiEnable && (1370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_2_io_out_valid_0) begin
			b_66_0 <=( _mesh_1_2_io_out_b_0) ^ ((fiEnable && (1371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1090_0 <=( _mesh_1_2_io_out_c_0) ^ ((fiEnable && (1372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_2_io_in_control_0_shift_b <=( _mesh_1_2_io_out_control_0_shift) ^ ((fiEnable && (1373 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_2_io_in_control_0_dataflow_b <=( _mesh_1_2_io_out_control_0_dataflow) ^ ((fiEnable && (1374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_2_io_in_control_0_propagate_b <=( _mesh_1_2_io_out_control_0_propagate) ^ ((fiEnable && (1375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_2_io_out_valid_0) begin
			b_67_0 <=( _mesh_2_2_io_out_b_0) ^ ((fiEnable && (1376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1091_0 <=( _mesh_2_2_io_out_c_0) ^ ((fiEnable && (1377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_2_io_in_control_0_shift_b <=( _mesh_2_2_io_out_control_0_shift) ^ ((fiEnable && (1378 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_2_io_in_control_0_dataflow_b <=( _mesh_2_2_io_out_control_0_dataflow) ^ ((fiEnable && (1379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_2_io_in_control_0_propagate_b <=( _mesh_2_2_io_out_control_0_propagate) ^ ((fiEnable && (1380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_2_io_out_valid_0) begin
			b_68_0 <=( _mesh_3_2_io_out_b_0) ^ ((fiEnable && (1381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1092_0 <=( _mesh_3_2_io_out_c_0) ^ ((fiEnable && (1382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_2_io_in_control_0_shift_b <=( _mesh_3_2_io_out_control_0_shift) ^ ((fiEnable && (1383 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_2_io_in_control_0_dataflow_b <=( _mesh_3_2_io_out_control_0_dataflow) ^ ((fiEnable && (1384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_2_io_in_control_0_propagate_b <=( _mesh_3_2_io_out_control_0_propagate) ^ ((fiEnable && (1385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_2_io_out_valid_0) begin
			b_69_0 <=( _mesh_4_2_io_out_b_0) ^ ((fiEnable && (1386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1093_0 <=( _mesh_4_2_io_out_c_0) ^ ((fiEnable && (1387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_2_io_in_control_0_shift_b <=( _mesh_4_2_io_out_control_0_shift) ^ ((fiEnable && (1388 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_2_io_in_control_0_dataflow_b <=( _mesh_4_2_io_out_control_0_dataflow) ^ ((fiEnable && (1389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_2_io_in_control_0_propagate_b <=( _mesh_4_2_io_out_control_0_propagate) ^ ((fiEnable && (1390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_2_io_out_valid_0) begin
			b_70_0 <=( _mesh_5_2_io_out_b_0) ^ ((fiEnable && (1391 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1094_0 <=( _mesh_5_2_io_out_c_0) ^ ((fiEnable && (1392 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_2_io_in_control_0_shift_b <=( _mesh_5_2_io_out_control_0_shift) ^ ((fiEnable && (1393 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_2_io_in_control_0_dataflow_b <=( _mesh_5_2_io_out_control_0_dataflow) ^ ((fiEnable && (1394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_2_io_in_control_0_propagate_b <=( _mesh_5_2_io_out_control_0_propagate) ^ ((fiEnable && (1395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_2_io_out_valid_0) begin
			b_71_0 <=( _mesh_6_2_io_out_b_0) ^ ((fiEnable && (1396 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1095_0 <=( _mesh_6_2_io_out_c_0) ^ ((fiEnable && (1397 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_2_io_in_control_0_shift_b <=( _mesh_6_2_io_out_control_0_shift) ^ ((fiEnable && (1398 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_2_io_in_control_0_dataflow_b <=( _mesh_6_2_io_out_control_0_dataflow) ^ ((fiEnable && (1399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_2_io_in_control_0_propagate_b <=( _mesh_6_2_io_out_control_0_propagate) ^ ((fiEnable && (1400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_2_io_out_valid_0) begin
			b_72_0 <=( _mesh_7_2_io_out_b_0) ^ ((fiEnable && (1401 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1096_0 <=( _mesh_7_2_io_out_c_0) ^ ((fiEnable && (1402 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_2_io_in_control_0_shift_b <=( _mesh_7_2_io_out_control_0_shift) ^ ((fiEnable && (1403 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_2_io_in_control_0_dataflow_b <=( _mesh_7_2_io_out_control_0_dataflow) ^ ((fiEnable && (1404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_2_io_in_control_0_propagate_b <=( _mesh_7_2_io_out_control_0_propagate) ^ ((fiEnable && (1405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_2_io_out_valid_0) begin
			b_73_0 <=( _mesh_8_2_io_out_b_0) ^ ((fiEnable && (1406 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1097_0 <=( _mesh_8_2_io_out_c_0) ^ ((fiEnable && (1407 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_2_io_in_control_0_shift_b <=( _mesh_8_2_io_out_control_0_shift) ^ ((fiEnable && (1408 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_2_io_in_control_0_dataflow_b <=( _mesh_8_2_io_out_control_0_dataflow) ^ ((fiEnable && (1409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_2_io_in_control_0_propagate_b <=( _mesh_8_2_io_out_control_0_propagate) ^ ((fiEnable && (1410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_2_io_out_valid_0) begin
			b_74_0 <=( _mesh_9_2_io_out_b_0) ^ ((fiEnable && (1411 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1098_0 <=( _mesh_9_2_io_out_c_0) ^ ((fiEnable && (1412 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_2_io_in_control_0_shift_b <=( _mesh_9_2_io_out_control_0_shift) ^ ((fiEnable && (1413 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_2_io_in_control_0_dataflow_b <=( _mesh_9_2_io_out_control_0_dataflow) ^ ((fiEnable && (1414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_2_io_in_control_0_propagate_b <=( _mesh_9_2_io_out_control_0_propagate) ^ ((fiEnable && (1415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_2_io_out_valid_0) begin
			b_75_0 <=( _mesh_10_2_io_out_b_0) ^ ((fiEnable && (1416 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1099_0 <=( _mesh_10_2_io_out_c_0) ^ ((fiEnable && (1417 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_2_io_in_control_0_shift_b <=( _mesh_10_2_io_out_control_0_shift) ^ ((fiEnable && (1418 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_2_io_in_control_0_dataflow_b <=( _mesh_10_2_io_out_control_0_dataflow) ^ ((fiEnable && (1419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_2_io_in_control_0_propagate_b <=( _mesh_10_2_io_out_control_0_propagate) ^ ((fiEnable && (1420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_2_io_out_valid_0) begin
			b_76_0 <=( _mesh_11_2_io_out_b_0) ^ ((fiEnable && (1421 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1100_0 <=( _mesh_11_2_io_out_c_0) ^ ((fiEnable && (1422 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_2_io_in_control_0_shift_b <=( _mesh_11_2_io_out_control_0_shift) ^ ((fiEnable && (1423 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_2_io_in_control_0_dataflow_b <=( _mesh_11_2_io_out_control_0_dataflow) ^ ((fiEnable && (1424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_2_io_in_control_0_propagate_b <=( _mesh_11_2_io_out_control_0_propagate) ^ ((fiEnable && (1425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_2_io_out_valid_0) begin
			b_77_0 <=( _mesh_12_2_io_out_b_0) ^ ((fiEnable && (1426 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1101_0 <=( _mesh_12_2_io_out_c_0) ^ ((fiEnable && (1427 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_2_io_in_control_0_shift_b <=( _mesh_12_2_io_out_control_0_shift) ^ ((fiEnable && (1428 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_2_io_in_control_0_dataflow_b <=( _mesh_12_2_io_out_control_0_dataflow) ^ ((fiEnable && (1429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_2_io_in_control_0_propagate_b <=( _mesh_12_2_io_out_control_0_propagate) ^ ((fiEnable && (1430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_2_io_out_valid_0) begin
			b_78_0 <=( _mesh_13_2_io_out_b_0) ^ ((fiEnable && (1431 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1102_0 <=( _mesh_13_2_io_out_c_0) ^ ((fiEnable && (1432 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_2_io_in_control_0_shift_b <=( _mesh_13_2_io_out_control_0_shift) ^ ((fiEnable && (1433 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_2_io_in_control_0_dataflow_b <=( _mesh_13_2_io_out_control_0_dataflow) ^ ((fiEnable && (1434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_2_io_in_control_0_propagate_b <=( _mesh_13_2_io_out_control_0_propagate) ^ ((fiEnable && (1435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_2_io_out_valid_0) begin
			b_79_0 <=( _mesh_14_2_io_out_b_0) ^ ((fiEnable && (1436 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1103_0 <=( _mesh_14_2_io_out_c_0) ^ ((fiEnable && (1437 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_2_io_in_control_0_shift_b <=( _mesh_14_2_io_out_control_0_shift) ^ ((fiEnable && (1438 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_2_io_in_control_0_dataflow_b <=( _mesh_14_2_io_out_control_0_dataflow) ^ ((fiEnable && (1439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_2_io_in_control_0_propagate_b <=( _mesh_14_2_io_out_control_0_propagate) ^ ((fiEnable && (1440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_2_io_out_valid_0) begin
			b_80_0 <=( _mesh_15_2_io_out_b_0) ^ ((fiEnable && (1441 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1104_0 <=( _mesh_15_2_io_out_c_0) ^ ((fiEnable && (1442 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_2_io_in_control_0_shift_b <=( _mesh_15_2_io_out_control_0_shift) ^ ((fiEnable && (1443 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_2_io_in_control_0_dataflow_b <=( _mesh_15_2_io_out_control_0_dataflow) ^ ((fiEnable && (1444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_2_io_in_control_0_propagate_b <=( _mesh_15_2_io_out_control_0_propagate) ^ ((fiEnable && (1445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_2_io_out_valid_0) begin
			b_81_0 <=( _mesh_16_2_io_out_b_0) ^ ((fiEnable && (1446 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1105_0 <=( _mesh_16_2_io_out_c_0) ^ ((fiEnable && (1447 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_2_io_in_control_0_shift_b <=( _mesh_16_2_io_out_control_0_shift) ^ ((fiEnable && (1448 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_2_io_in_control_0_dataflow_b <=( _mesh_16_2_io_out_control_0_dataflow) ^ ((fiEnable && (1449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_2_io_in_control_0_propagate_b <=( _mesh_16_2_io_out_control_0_propagate) ^ ((fiEnable && (1450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_2_io_out_valid_0) begin
			b_82_0 <=( _mesh_17_2_io_out_b_0) ^ ((fiEnable && (1451 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1106_0 <=( _mesh_17_2_io_out_c_0) ^ ((fiEnable && (1452 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_2_io_in_control_0_shift_b <=( _mesh_17_2_io_out_control_0_shift) ^ ((fiEnable && (1453 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_2_io_in_control_0_dataflow_b <=( _mesh_17_2_io_out_control_0_dataflow) ^ ((fiEnable && (1454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_2_io_in_control_0_propagate_b <=( _mesh_17_2_io_out_control_0_propagate) ^ ((fiEnable && (1455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_2_io_out_valid_0) begin
			b_83_0 <=( _mesh_18_2_io_out_b_0) ^ ((fiEnable && (1456 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1107_0 <=( _mesh_18_2_io_out_c_0) ^ ((fiEnable && (1457 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_2_io_in_control_0_shift_b <=( _mesh_18_2_io_out_control_0_shift) ^ ((fiEnable && (1458 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_2_io_in_control_0_dataflow_b <=( _mesh_18_2_io_out_control_0_dataflow) ^ ((fiEnable && (1459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_2_io_in_control_0_propagate_b <=( _mesh_18_2_io_out_control_0_propagate) ^ ((fiEnable && (1460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_2_io_out_valid_0) begin
			b_84_0 <=( _mesh_19_2_io_out_b_0) ^ ((fiEnable && (1461 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1108_0 <=( _mesh_19_2_io_out_c_0) ^ ((fiEnable && (1462 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_2_io_in_control_0_shift_b <=( _mesh_19_2_io_out_control_0_shift) ^ ((fiEnable && (1463 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_2_io_in_control_0_dataflow_b <=( _mesh_19_2_io_out_control_0_dataflow) ^ ((fiEnable && (1464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_2_io_in_control_0_propagate_b <=( _mesh_19_2_io_out_control_0_propagate) ^ ((fiEnable && (1465 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_2_io_out_valid_0) begin
			b_85_0 <=( _mesh_20_2_io_out_b_0) ^ ((fiEnable && (1466 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1109_0 <=( _mesh_20_2_io_out_c_0) ^ ((fiEnable && (1467 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_2_io_in_control_0_shift_b <=( _mesh_20_2_io_out_control_0_shift) ^ ((fiEnable && (1468 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_2_io_in_control_0_dataflow_b <=( _mesh_20_2_io_out_control_0_dataflow) ^ ((fiEnable && (1469 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_2_io_in_control_0_propagate_b <=( _mesh_20_2_io_out_control_0_propagate) ^ ((fiEnable && (1470 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_2_io_out_valid_0) begin
			b_86_0 <=( _mesh_21_2_io_out_b_0) ^ ((fiEnable && (1471 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1110_0 <=( _mesh_21_2_io_out_c_0) ^ ((fiEnable && (1472 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_2_io_in_control_0_shift_b <=( _mesh_21_2_io_out_control_0_shift) ^ ((fiEnable && (1473 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_2_io_in_control_0_dataflow_b <=( _mesh_21_2_io_out_control_0_dataflow) ^ ((fiEnable && (1474 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_2_io_in_control_0_propagate_b <=( _mesh_21_2_io_out_control_0_propagate) ^ ((fiEnable && (1475 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_2_io_out_valid_0) begin
			b_87_0 <=( _mesh_22_2_io_out_b_0) ^ ((fiEnable && (1476 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1111_0 <=( _mesh_22_2_io_out_c_0) ^ ((fiEnable && (1477 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_2_io_in_control_0_shift_b <=( _mesh_22_2_io_out_control_0_shift) ^ ((fiEnable && (1478 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_2_io_in_control_0_dataflow_b <=( _mesh_22_2_io_out_control_0_dataflow) ^ ((fiEnable && (1479 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_2_io_in_control_0_propagate_b <=( _mesh_22_2_io_out_control_0_propagate) ^ ((fiEnable && (1480 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_2_io_out_valid_0) begin
			b_88_0 <=( _mesh_23_2_io_out_b_0) ^ ((fiEnable && (1481 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1112_0 <=( _mesh_23_2_io_out_c_0) ^ ((fiEnable && (1482 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_2_io_in_control_0_shift_b <=( _mesh_23_2_io_out_control_0_shift) ^ ((fiEnable && (1483 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_2_io_in_control_0_dataflow_b <=( _mesh_23_2_io_out_control_0_dataflow) ^ ((fiEnable && (1484 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_2_io_in_control_0_propagate_b <=( _mesh_23_2_io_out_control_0_propagate) ^ ((fiEnable && (1485 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_2_io_out_valid_0) begin
			b_89_0 <=( _mesh_24_2_io_out_b_0) ^ ((fiEnable && (1486 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1113_0 <=( _mesh_24_2_io_out_c_0) ^ ((fiEnable && (1487 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_2_io_in_control_0_shift_b <=( _mesh_24_2_io_out_control_0_shift) ^ ((fiEnable && (1488 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_2_io_in_control_0_dataflow_b <=( _mesh_24_2_io_out_control_0_dataflow) ^ ((fiEnable && (1489 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_2_io_in_control_0_propagate_b <=( _mesh_24_2_io_out_control_0_propagate) ^ ((fiEnable && (1490 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_2_io_out_valid_0) begin
			b_90_0 <=( _mesh_25_2_io_out_b_0) ^ ((fiEnable && (1491 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1114_0 <=( _mesh_25_2_io_out_c_0) ^ ((fiEnable && (1492 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_2_io_in_control_0_shift_b <=( _mesh_25_2_io_out_control_0_shift) ^ ((fiEnable && (1493 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_2_io_in_control_0_dataflow_b <=( _mesh_25_2_io_out_control_0_dataflow) ^ ((fiEnable && (1494 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_2_io_in_control_0_propagate_b <=( _mesh_25_2_io_out_control_0_propagate) ^ ((fiEnable && (1495 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_2_io_out_valid_0) begin
			b_91_0 <=( _mesh_26_2_io_out_b_0) ^ ((fiEnable && (1496 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1115_0 <=( _mesh_26_2_io_out_c_0) ^ ((fiEnable && (1497 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_2_io_in_control_0_shift_b <=( _mesh_26_2_io_out_control_0_shift) ^ ((fiEnable && (1498 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_2_io_in_control_0_dataflow_b <=( _mesh_26_2_io_out_control_0_dataflow) ^ ((fiEnable && (1499 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_2_io_in_control_0_propagate_b <=( _mesh_26_2_io_out_control_0_propagate) ^ ((fiEnable && (1500 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_2_io_out_valid_0) begin
			b_92_0 <=( _mesh_27_2_io_out_b_0) ^ ((fiEnable && (1501 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1116_0 <=( _mesh_27_2_io_out_c_0) ^ ((fiEnable && (1502 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_2_io_in_control_0_shift_b <=( _mesh_27_2_io_out_control_0_shift) ^ ((fiEnable && (1503 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_2_io_in_control_0_dataflow_b <=( _mesh_27_2_io_out_control_0_dataflow) ^ ((fiEnable && (1504 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_2_io_in_control_0_propagate_b <=( _mesh_27_2_io_out_control_0_propagate) ^ ((fiEnable && (1505 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_2_io_out_valid_0) begin
			b_93_0 <=( _mesh_28_2_io_out_b_0) ^ ((fiEnable && (1506 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1117_0 <=( _mesh_28_2_io_out_c_0) ^ ((fiEnable && (1507 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_2_io_in_control_0_shift_b <=( _mesh_28_2_io_out_control_0_shift) ^ ((fiEnable && (1508 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_2_io_in_control_0_dataflow_b <=( _mesh_28_2_io_out_control_0_dataflow) ^ ((fiEnable && (1509 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_2_io_in_control_0_propagate_b <=( _mesh_28_2_io_out_control_0_propagate) ^ ((fiEnable && (1510 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_2_io_out_valid_0) begin
			b_94_0 <=( _mesh_29_2_io_out_b_0) ^ ((fiEnable && (1511 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1118_0 <=( _mesh_29_2_io_out_c_0) ^ ((fiEnable && (1512 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_2_io_in_control_0_shift_b <=( _mesh_29_2_io_out_control_0_shift) ^ ((fiEnable && (1513 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_2_io_in_control_0_dataflow_b <=( _mesh_29_2_io_out_control_0_dataflow) ^ ((fiEnable && (1514 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_2_io_in_control_0_propagate_b <=( _mesh_29_2_io_out_control_0_propagate) ^ ((fiEnable && (1515 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_2_io_out_valid_0) begin
			b_95_0 <=( _mesh_30_2_io_out_b_0) ^ ((fiEnable && (1516 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1119_0 <=( _mesh_30_2_io_out_c_0) ^ ((fiEnable && (1517 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_2_io_in_control_0_shift_b <=( _mesh_30_2_io_out_control_0_shift) ^ ((fiEnable && (1518 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_2_io_in_control_0_dataflow_b <=( _mesh_30_2_io_out_control_0_dataflow) ^ ((fiEnable && (1519 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_2_io_in_control_0_propagate_b <=( _mesh_30_2_io_out_control_0_propagate) ^ ((fiEnable && (1520 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_3_0) begin
			b_96_0 <=( io_in_b_3_0) ^ ((fiEnable && (1521 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1120_0 <=( io_in_d_3_0) ^ ((fiEnable && (1522 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_3_io_in_control_0_shift_b <=( io_in_control_3_0_shift) ^ ((fiEnable && (1523 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_3_io_in_control_0_dataflow_b <=( io_in_control_3_0_dataflow) ^ ((fiEnable && (1524 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_3_io_in_control_0_propagate_b <=( io_in_control_3_0_propagate) ^ ((fiEnable && (1525 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_3_io_out_valid_0) begin
			b_97_0 <=( _mesh_0_3_io_out_b_0) ^ ((fiEnable && (1526 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1121_0 <=( _mesh_0_3_io_out_c_0) ^ ((fiEnable && (1527 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_3_io_in_control_0_shift_b <=( _mesh_0_3_io_out_control_0_shift) ^ ((fiEnable && (1528 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_3_io_in_control_0_dataflow_b <=( _mesh_0_3_io_out_control_0_dataflow) ^ ((fiEnable && (1529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_3_io_in_control_0_propagate_b <=( _mesh_0_3_io_out_control_0_propagate) ^ ((fiEnable && (1530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_3_io_out_valid_0) begin
			b_98_0 <=( _mesh_1_3_io_out_b_0) ^ ((fiEnable && (1531 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1122_0 <=( _mesh_1_3_io_out_c_0) ^ ((fiEnable && (1532 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_3_io_in_control_0_shift_b <=( _mesh_1_3_io_out_control_0_shift) ^ ((fiEnable && (1533 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_3_io_in_control_0_dataflow_b <=( _mesh_1_3_io_out_control_0_dataflow) ^ ((fiEnable && (1534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_3_io_in_control_0_propagate_b <=( _mesh_1_3_io_out_control_0_propagate) ^ ((fiEnable && (1535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_3_io_out_valid_0) begin
			b_99_0 <=( _mesh_2_3_io_out_b_0) ^ ((fiEnable && (1536 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1123_0 <=( _mesh_2_3_io_out_c_0) ^ ((fiEnable && (1537 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_3_io_in_control_0_shift_b <=( _mesh_2_3_io_out_control_0_shift) ^ ((fiEnable && (1538 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_3_io_in_control_0_dataflow_b <=( _mesh_2_3_io_out_control_0_dataflow) ^ ((fiEnable && (1539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_3_io_in_control_0_propagate_b <=( _mesh_2_3_io_out_control_0_propagate) ^ ((fiEnable && (1540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_3_io_out_valid_0) begin
			b_100_0 <=( _mesh_3_3_io_out_b_0) ^ ((fiEnable && (1541 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1124_0 <=( _mesh_3_3_io_out_c_0) ^ ((fiEnable && (1542 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_3_io_in_control_0_shift_b <=( _mesh_3_3_io_out_control_0_shift) ^ ((fiEnable && (1543 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_3_io_in_control_0_dataflow_b <=( _mesh_3_3_io_out_control_0_dataflow) ^ ((fiEnable && (1544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_3_io_in_control_0_propagate_b <=( _mesh_3_3_io_out_control_0_propagate) ^ ((fiEnable && (1545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_3_io_out_valid_0) begin
			b_101_0 <=( _mesh_4_3_io_out_b_0) ^ ((fiEnable && (1546 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1125_0 <=( _mesh_4_3_io_out_c_0) ^ ((fiEnable && (1547 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_3_io_in_control_0_shift_b <=( _mesh_4_3_io_out_control_0_shift) ^ ((fiEnable && (1548 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_3_io_in_control_0_dataflow_b <=( _mesh_4_3_io_out_control_0_dataflow) ^ ((fiEnable && (1549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_3_io_in_control_0_propagate_b <=( _mesh_4_3_io_out_control_0_propagate) ^ ((fiEnable && (1550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_3_io_out_valid_0) begin
			b_102_0 <=( _mesh_5_3_io_out_b_0) ^ ((fiEnable && (1551 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1126_0 <=( _mesh_5_3_io_out_c_0) ^ ((fiEnable && (1552 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_3_io_in_control_0_shift_b <=( _mesh_5_3_io_out_control_0_shift) ^ ((fiEnable && (1553 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_3_io_in_control_0_dataflow_b <=( _mesh_5_3_io_out_control_0_dataflow) ^ ((fiEnable && (1554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_3_io_in_control_0_propagate_b <=( _mesh_5_3_io_out_control_0_propagate) ^ ((fiEnable && (1555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_3_io_out_valid_0) begin
			b_103_0 <=( _mesh_6_3_io_out_b_0) ^ ((fiEnable && (1556 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1127_0 <=( _mesh_6_3_io_out_c_0) ^ ((fiEnable && (1557 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_3_io_in_control_0_shift_b <=( _mesh_6_3_io_out_control_0_shift) ^ ((fiEnable && (1558 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_3_io_in_control_0_dataflow_b <=( _mesh_6_3_io_out_control_0_dataflow) ^ ((fiEnable && (1559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_3_io_in_control_0_propagate_b <=( _mesh_6_3_io_out_control_0_propagate) ^ ((fiEnable && (1560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_3_io_out_valid_0) begin
			b_104_0 <=( _mesh_7_3_io_out_b_0) ^ ((fiEnable && (1561 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1128_0 <=( _mesh_7_3_io_out_c_0) ^ ((fiEnable && (1562 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_3_io_in_control_0_shift_b <=( _mesh_7_3_io_out_control_0_shift) ^ ((fiEnable && (1563 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_3_io_in_control_0_dataflow_b <=( _mesh_7_3_io_out_control_0_dataflow) ^ ((fiEnable && (1564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_3_io_in_control_0_propagate_b <=( _mesh_7_3_io_out_control_0_propagate) ^ ((fiEnable && (1565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_3_io_out_valid_0) begin
			b_105_0 <=( _mesh_8_3_io_out_b_0) ^ ((fiEnable && (1566 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1129_0 <=( _mesh_8_3_io_out_c_0) ^ ((fiEnable && (1567 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_3_io_in_control_0_shift_b <=( _mesh_8_3_io_out_control_0_shift) ^ ((fiEnable && (1568 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_3_io_in_control_0_dataflow_b <=( _mesh_8_3_io_out_control_0_dataflow) ^ ((fiEnable && (1569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_3_io_in_control_0_propagate_b <=( _mesh_8_3_io_out_control_0_propagate) ^ ((fiEnable && (1570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_3_io_out_valid_0) begin
			b_106_0 <=( _mesh_9_3_io_out_b_0) ^ ((fiEnable && (1571 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1130_0 <=( _mesh_9_3_io_out_c_0) ^ ((fiEnable && (1572 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_3_io_in_control_0_shift_b <=( _mesh_9_3_io_out_control_0_shift) ^ ((fiEnable && (1573 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_3_io_in_control_0_dataflow_b <=( _mesh_9_3_io_out_control_0_dataflow) ^ ((fiEnable && (1574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_3_io_in_control_0_propagate_b <=( _mesh_9_3_io_out_control_0_propagate) ^ ((fiEnable && (1575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_3_io_out_valid_0) begin
			b_107_0 <=( _mesh_10_3_io_out_b_0) ^ ((fiEnable && (1576 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1131_0 <=( _mesh_10_3_io_out_c_0) ^ ((fiEnable && (1577 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_3_io_in_control_0_shift_b <=( _mesh_10_3_io_out_control_0_shift) ^ ((fiEnable && (1578 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_3_io_in_control_0_dataflow_b <=( _mesh_10_3_io_out_control_0_dataflow) ^ ((fiEnable && (1579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_3_io_in_control_0_propagate_b <=( _mesh_10_3_io_out_control_0_propagate) ^ ((fiEnable && (1580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_3_io_out_valid_0) begin
			b_108_0 <=( _mesh_11_3_io_out_b_0) ^ ((fiEnable && (1581 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1132_0 <=( _mesh_11_3_io_out_c_0) ^ ((fiEnable && (1582 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_3_io_in_control_0_shift_b <=( _mesh_11_3_io_out_control_0_shift) ^ ((fiEnable && (1583 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_3_io_in_control_0_dataflow_b <=( _mesh_11_3_io_out_control_0_dataflow) ^ ((fiEnable && (1584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_3_io_in_control_0_propagate_b <=( _mesh_11_3_io_out_control_0_propagate) ^ ((fiEnable && (1585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_3_io_out_valid_0) begin
			b_109_0 <=( _mesh_12_3_io_out_b_0) ^ ((fiEnable && (1586 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1133_0 <=( _mesh_12_3_io_out_c_0) ^ ((fiEnable && (1587 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_3_io_in_control_0_shift_b <=( _mesh_12_3_io_out_control_0_shift) ^ ((fiEnable && (1588 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_3_io_in_control_0_dataflow_b <=( _mesh_12_3_io_out_control_0_dataflow) ^ ((fiEnable && (1589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_3_io_in_control_0_propagate_b <=( _mesh_12_3_io_out_control_0_propagate) ^ ((fiEnable && (1590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_3_io_out_valid_0) begin
			b_110_0 <=( _mesh_13_3_io_out_b_0) ^ ((fiEnable && (1591 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1134_0 <=( _mesh_13_3_io_out_c_0) ^ ((fiEnable && (1592 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_3_io_in_control_0_shift_b <=( _mesh_13_3_io_out_control_0_shift) ^ ((fiEnable && (1593 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_3_io_in_control_0_dataflow_b <=( _mesh_13_3_io_out_control_0_dataflow) ^ ((fiEnable && (1594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_3_io_in_control_0_propagate_b <=( _mesh_13_3_io_out_control_0_propagate) ^ ((fiEnable && (1595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_3_io_out_valid_0) begin
			b_111_0 <=( _mesh_14_3_io_out_b_0) ^ ((fiEnable && (1596 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1135_0 <=( _mesh_14_3_io_out_c_0) ^ ((fiEnable && (1597 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_3_io_in_control_0_shift_b <=( _mesh_14_3_io_out_control_0_shift) ^ ((fiEnable && (1598 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_3_io_in_control_0_dataflow_b <=( _mesh_14_3_io_out_control_0_dataflow) ^ ((fiEnable && (1599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_3_io_in_control_0_propagate_b <=( _mesh_14_3_io_out_control_0_propagate) ^ ((fiEnable && (1600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_3_io_out_valid_0) begin
			b_112_0 <=( _mesh_15_3_io_out_b_0) ^ ((fiEnable && (1601 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1136_0 <=( _mesh_15_3_io_out_c_0) ^ ((fiEnable && (1602 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_3_io_in_control_0_shift_b <=( _mesh_15_3_io_out_control_0_shift) ^ ((fiEnable && (1603 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_3_io_in_control_0_dataflow_b <=( _mesh_15_3_io_out_control_0_dataflow) ^ ((fiEnable && (1604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_3_io_in_control_0_propagate_b <=( _mesh_15_3_io_out_control_0_propagate) ^ ((fiEnable && (1605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_3_io_out_valid_0) begin
			b_113_0 <=( _mesh_16_3_io_out_b_0) ^ ((fiEnable && (1606 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1137_0 <=( _mesh_16_3_io_out_c_0) ^ ((fiEnable && (1607 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_3_io_in_control_0_shift_b <=( _mesh_16_3_io_out_control_0_shift) ^ ((fiEnable && (1608 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_3_io_in_control_0_dataflow_b <=( _mesh_16_3_io_out_control_0_dataflow) ^ ((fiEnable && (1609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_3_io_in_control_0_propagate_b <=( _mesh_16_3_io_out_control_0_propagate) ^ ((fiEnable && (1610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_3_io_out_valid_0) begin
			b_114_0 <=( _mesh_17_3_io_out_b_0) ^ ((fiEnable && (1611 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1138_0 <=( _mesh_17_3_io_out_c_0) ^ ((fiEnable && (1612 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_3_io_in_control_0_shift_b <=( _mesh_17_3_io_out_control_0_shift) ^ ((fiEnable && (1613 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_3_io_in_control_0_dataflow_b <=( _mesh_17_3_io_out_control_0_dataflow) ^ ((fiEnable && (1614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_3_io_in_control_0_propagate_b <=( _mesh_17_3_io_out_control_0_propagate) ^ ((fiEnable && (1615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_3_io_out_valid_0) begin
			b_115_0 <=( _mesh_18_3_io_out_b_0) ^ ((fiEnable && (1616 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1139_0 <=( _mesh_18_3_io_out_c_0) ^ ((fiEnable && (1617 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_3_io_in_control_0_shift_b <=( _mesh_18_3_io_out_control_0_shift) ^ ((fiEnable && (1618 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_3_io_in_control_0_dataflow_b <=( _mesh_18_3_io_out_control_0_dataflow) ^ ((fiEnable && (1619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_3_io_in_control_0_propagate_b <=( _mesh_18_3_io_out_control_0_propagate) ^ ((fiEnable && (1620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_3_io_out_valid_0) begin
			b_116_0 <=( _mesh_19_3_io_out_b_0) ^ ((fiEnable && (1621 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1140_0 <=( _mesh_19_3_io_out_c_0) ^ ((fiEnable && (1622 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_3_io_in_control_0_shift_b <=( _mesh_19_3_io_out_control_0_shift) ^ ((fiEnable && (1623 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_3_io_in_control_0_dataflow_b <=( _mesh_19_3_io_out_control_0_dataflow) ^ ((fiEnable && (1624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_3_io_in_control_0_propagate_b <=( _mesh_19_3_io_out_control_0_propagate) ^ ((fiEnable && (1625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_3_io_out_valid_0) begin
			b_117_0 <=( _mesh_20_3_io_out_b_0) ^ ((fiEnable && (1626 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1141_0 <=( _mesh_20_3_io_out_c_0) ^ ((fiEnable && (1627 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_3_io_in_control_0_shift_b <=( _mesh_20_3_io_out_control_0_shift) ^ ((fiEnable && (1628 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_3_io_in_control_0_dataflow_b <=( _mesh_20_3_io_out_control_0_dataflow) ^ ((fiEnable && (1629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_3_io_in_control_0_propagate_b <=( _mesh_20_3_io_out_control_0_propagate) ^ ((fiEnable && (1630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_3_io_out_valid_0) begin
			b_118_0 <=( _mesh_21_3_io_out_b_0) ^ ((fiEnable && (1631 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1142_0 <=( _mesh_21_3_io_out_c_0) ^ ((fiEnable && (1632 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_3_io_in_control_0_shift_b <=( _mesh_21_3_io_out_control_0_shift) ^ ((fiEnable && (1633 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_3_io_in_control_0_dataflow_b <=( _mesh_21_3_io_out_control_0_dataflow) ^ ((fiEnable && (1634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_3_io_in_control_0_propagate_b <=( _mesh_21_3_io_out_control_0_propagate) ^ ((fiEnable && (1635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_3_io_out_valid_0) begin
			b_119_0 <=( _mesh_22_3_io_out_b_0) ^ ((fiEnable && (1636 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1143_0 <=( _mesh_22_3_io_out_c_0) ^ ((fiEnable && (1637 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_3_io_in_control_0_shift_b <=( _mesh_22_3_io_out_control_0_shift) ^ ((fiEnable && (1638 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_3_io_in_control_0_dataflow_b <=( _mesh_22_3_io_out_control_0_dataflow) ^ ((fiEnable && (1639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_3_io_in_control_0_propagate_b <=( _mesh_22_3_io_out_control_0_propagate) ^ ((fiEnable && (1640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_3_io_out_valid_0) begin
			b_120_0 <=( _mesh_23_3_io_out_b_0) ^ ((fiEnable && (1641 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1144_0 <=( _mesh_23_3_io_out_c_0) ^ ((fiEnable && (1642 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_3_io_in_control_0_shift_b <=( _mesh_23_3_io_out_control_0_shift) ^ ((fiEnable && (1643 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_3_io_in_control_0_dataflow_b <=( _mesh_23_3_io_out_control_0_dataflow) ^ ((fiEnable && (1644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_3_io_in_control_0_propagate_b <=( _mesh_23_3_io_out_control_0_propagate) ^ ((fiEnable && (1645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_3_io_out_valid_0) begin
			b_121_0 <=( _mesh_24_3_io_out_b_0) ^ ((fiEnable && (1646 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1145_0 <=( _mesh_24_3_io_out_c_0) ^ ((fiEnable && (1647 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_3_io_in_control_0_shift_b <=( _mesh_24_3_io_out_control_0_shift) ^ ((fiEnable && (1648 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_3_io_in_control_0_dataflow_b <=( _mesh_24_3_io_out_control_0_dataflow) ^ ((fiEnable && (1649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_3_io_in_control_0_propagate_b <=( _mesh_24_3_io_out_control_0_propagate) ^ ((fiEnable && (1650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_3_io_out_valid_0) begin
			b_122_0 <=( _mesh_25_3_io_out_b_0) ^ ((fiEnable && (1651 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1146_0 <=( _mesh_25_3_io_out_c_0) ^ ((fiEnable && (1652 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_3_io_in_control_0_shift_b <=( _mesh_25_3_io_out_control_0_shift) ^ ((fiEnable && (1653 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_3_io_in_control_0_dataflow_b <=( _mesh_25_3_io_out_control_0_dataflow) ^ ((fiEnable && (1654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_3_io_in_control_0_propagate_b <=( _mesh_25_3_io_out_control_0_propagate) ^ ((fiEnable && (1655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_3_io_out_valid_0) begin
			b_123_0 <=( _mesh_26_3_io_out_b_0) ^ ((fiEnable && (1656 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1147_0 <=( _mesh_26_3_io_out_c_0) ^ ((fiEnable && (1657 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_3_io_in_control_0_shift_b <=( _mesh_26_3_io_out_control_0_shift) ^ ((fiEnable && (1658 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_3_io_in_control_0_dataflow_b <=( _mesh_26_3_io_out_control_0_dataflow) ^ ((fiEnable && (1659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_3_io_in_control_0_propagate_b <=( _mesh_26_3_io_out_control_0_propagate) ^ ((fiEnable && (1660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_3_io_out_valid_0) begin
			b_124_0 <=( _mesh_27_3_io_out_b_0) ^ ((fiEnable && (1661 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1148_0 <=( _mesh_27_3_io_out_c_0) ^ ((fiEnable && (1662 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_3_io_in_control_0_shift_b <=( _mesh_27_3_io_out_control_0_shift) ^ ((fiEnable && (1663 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_3_io_in_control_0_dataflow_b <=( _mesh_27_3_io_out_control_0_dataflow) ^ ((fiEnable && (1664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_3_io_in_control_0_propagate_b <=( _mesh_27_3_io_out_control_0_propagate) ^ ((fiEnable && (1665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_3_io_out_valid_0) begin
			b_125_0 <=( _mesh_28_3_io_out_b_0) ^ ((fiEnable && (1666 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1149_0 <=( _mesh_28_3_io_out_c_0) ^ ((fiEnable && (1667 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_3_io_in_control_0_shift_b <=( _mesh_28_3_io_out_control_0_shift) ^ ((fiEnable && (1668 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_3_io_in_control_0_dataflow_b <=( _mesh_28_3_io_out_control_0_dataflow) ^ ((fiEnable && (1669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_3_io_in_control_0_propagate_b <=( _mesh_28_3_io_out_control_0_propagate) ^ ((fiEnable && (1670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_3_io_out_valid_0) begin
			b_126_0 <=( _mesh_29_3_io_out_b_0) ^ ((fiEnable && (1671 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1150_0 <=( _mesh_29_3_io_out_c_0) ^ ((fiEnable && (1672 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_3_io_in_control_0_shift_b <=( _mesh_29_3_io_out_control_0_shift) ^ ((fiEnable && (1673 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_3_io_in_control_0_dataflow_b <=( _mesh_29_3_io_out_control_0_dataflow) ^ ((fiEnable && (1674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_3_io_in_control_0_propagate_b <=( _mesh_29_3_io_out_control_0_propagate) ^ ((fiEnable && (1675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_3_io_out_valid_0) begin
			b_127_0 <=( _mesh_30_3_io_out_b_0) ^ ((fiEnable && (1676 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1151_0 <=( _mesh_30_3_io_out_c_0) ^ ((fiEnable && (1677 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_3_io_in_control_0_shift_b <=( _mesh_30_3_io_out_control_0_shift) ^ ((fiEnable && (1678 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_3_io_in_control_0_dataflow_b <=( _mesh_30_3_io_out_control_0_dataflow) ^ ((fiEnable && (1679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_3_io_in_control_0_propagate_b <=( _mesh_30_3_io_out_control_0_propagate) ^ ((fiEnable && (1680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_4_0) begin
			b_128_0 <=( io_in_b_4_0) ^ ((fiEnable && (1681 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1152_0 <=( io_in_d_4_0) ^ ((fiEnable && (1682 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_4_io_in_control_0_shift_b <=( io_in_control_4_0_shift) ^ ((fiEnable && (1683 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_4_io_in_control_0_dataflow_b <=( io_in_control_4_0_dataflow) ^ ((fiEnable && (1684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_4_io_in_control_0_propagate_b <=( io_in_control_4_0_propagate) ^ ((fiEnable && (1685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_4_io_out_valid_0) begin
			b_129_0 <=( _mesh_0_4_io_out_b_0) ^ ((fiEnable && (1686 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1153_0 <=( _mesh_0_4_io_out_c_0) ^ ((fiEnable && (1687 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_4_io_in_control_0_shift_b <=( _mesh_0_4_io_out_control_0_shift) ^ ((fiEnable && (1688 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_4_io_in_control_0_dataflow_b <=( _mesh_0_4_io_out_control_0_dataflow) ^ ((fiEnable && (1689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_4_io_in_control_0_propagate_b <=( _mesh_0_4_io_out_control_0_propagate) ^ ((fiEnable && (1690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_4_io_out_valid_0) begin
			b_130_0 <=( _mesh_1_4_io_out_b_0) ^ ((fiEnable && (1691 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1154_0 <=( _mesh_1_4_io_out_c_0) ^ ((fiEnable && (1692 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_4_io_in_control_0_shift_b <=( _mesh_1_4_io_out_control_0_shift) ^ ((fiEnable && (1693 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_4_io_in_control_0_dataflow_b <=( _mesh_1_4_io_out_control_0_dataflow) ^ ((fiEnable && (1694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_4_io_in_control_0_propagate_b <=( _mesh_1_4_io_out_control_0_propagate) ^ ((fiEnable && (1695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_4_io_out_valid_0) begin
			b_131_0 <=( _mesh_2_4_io_out_b_0) ^ ((fiEnable && (1696 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1155_0 <=( _mesh_2_4_io_out_c_0) ^ ((fiEnable && (1697 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_4_io_in_control_0_shift_b <=( _mesh_2_4_io_out_control_0_shift) ^ ((fiEnable && (1698 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_4_io_in_control_0_dataflow_b <=( _mesh_2_4_io_out_control_0_dataflow) ^ ((fiEnable && (1699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_4_io_in_control_0_propagate_b <=( _mesh_2_4_io_out_control_0_propagate) ^ ((fiEnable && (1700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_4_io_out_valid_0) begin
			b_132_0 <=( _mesh_3_4_io_out_b_0) ^ ((fiEnable && (1701 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1156_0 <=( _mesh_3_4_io_out_c_0) ^ ((fiEnable && (1702 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_4_io_in_control_0_shift_b <=( _mesh_3_4_io_out_control_0_shift) ^ ((fiEnable && (1703 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_4_io_in_control_0_dataflow_b <=( _mesh_3_4_io_out_control_0_dataflow) ^ ((fiEnable && (1704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_4_io_in_control_0_propagate_b <=( _mesh_3_4_io_out_control_0_propagate) ^ ((fiEnable && (1705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_4_io_out_valid_0) begin
			b_133_0 <=( _mesh_4_4_io_out_b_0) ^ ((fiEnable && (1706 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1157_0 <=( _mesh_4_4_io_out_c_0) ^ ((fiEnable && (1707 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_4_io_in_control_0_shift_b <=( _mesh_4_4_io_out_control_0_shift) ^ ((fiEnable && (1708 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_4_io_in_control_0_dataflow_b <=( _mesh_4_4_io_out_control_0_dataflow) ^ ((fiEnable && (1709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_4_io_in_control_0_propagate_b <=( _mesh_4_4_io_out_control_0_propagate) ^ ((fiEnable && (1710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_4_io_out_valid_0) begin
			b_134_0 <=( _mesh_5_4_io_out_b_0) ^ ((fiEnable && (1711 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1158_0 <=( _mesh_5_4_io_out_c_0) ^ ((fiEnable && (1712 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_4_io_in_control_0_shift_b <=( _mesh_5_4_io_out_control_0_shift) ^ ((fiEnable && (1713 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_4_io_in_control_0_dataflow_b <=( _mesh_5_4_io_out_control_0_dataflow) ^ ((fiEnable && (1714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_4_io_in_control_0_propagate_b <=( _mesh_5_4_io_out_control_0_propagate) ^ ((fiEnable && (1715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_4_io_out_valid_0) begin
			b_135_0 <=( _mesh_6_4_io_out_b_0) ^ ((fiEnable && (1716 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1159_0 <=( _mesh_6_4_io_out_c_0) ^ ((fiEnable && (1717 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_4_io_in_control_0_shift_b <=( _mesh_6_4_io_out_control_0_shift) ^ ((fiEnable && (1718 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_4_io_in_control_0_dataflow_b <=( _mesh_6_4_io_out_control_0_dataflow) ^ ((fiEnable && (1719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_4_io_in_control_0_propagate_b <=( _mesh_6_4_io_out_control_0_propagate) ^ ((fiEnable && (1720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_4_io_out_valid_0) begin
			b_136_0 <=( _mesh_7_4_io_out_b_0) ^ ((fiEnable && (1721 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1160_0 <=( _mesh_7_4_io_out_c_0) ^ ((fiEnable && (1722 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_4_io_in_control_0_shift_b <=( _mesh_7_4_io_out_control_0_shift) ^ ((fiEnable && (1723 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_4_io_in_control_0_dataflow_b <=( _mesh_7_4_io_out_control_0_dataflow) ^ ((fiEnable && (1724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_4_io_in_control_0_propagate_b <=( _mesh_7_4_io_out_control_0_propagate) ^ ((fiEnable && (1725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_4_io_out_valid_0) begin
			b_137_0 <=( _mesh_8_4_io_out_b_0) ^ ((fiEnable && (1726 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1161_0 <=( _mesh_8_4_io_out_c_0) ^ ((fiEnable && (1727 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_4_io_in_control_0_shift_b <=( _mesh_8_4_io_out_control_0_shift) ^ ((fiEnable && (1728 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_4_io_in_control_0_dataflow_b <=( _mesh_8_4_io_out_control_0_dataflow) ^ ((fiEnable && (1729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_4_io_in_control_0_propagate_b <=( _mesh_8_4_io_out_control_0_propagate) ^ ((fiEnable && (1730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_4_io_out_valid_0) begin
			b_138_0 <=( _mesh_9_4_io_out_b_0) ^ ((fiEnable && (1731 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1162_0 <=( _mesh_9_4_io_out_c_0) ^ ((fiEnable && (1732 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_4_io_in_control_0_shift_b <=( _mesh_9_4_io_out_control_0_shift) ^ ((fiEnable && (1733 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_4_io_in_control_0_dataflow_b <=( _mesh_9_4_io_out_control_0_dataflow) ^ ((fiEnable && (1734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_4_io_in_control_0_propagate_b <=( _mesh_9_4_io_out_control_0_propagate) ^ ((fiEnable && (1735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_4_io_out_valid_0) begin
			b_139_0 <=( _mesh_10_4_io_out_b_0) ^ ((fiEnable && (1736 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1163_0 <=( _mesh_10_4_io_out_c_0) ^ ((fiEnable && (1737 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_4_io_in_control_0_shift_b <=( _mesh_10_4_io_out_control_0_shift) ^ ((fiEnable && (1738 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_4_io_in_control_0_dataflow_b <=( _mesh_10_4_io_out_control_0_dataflow) ^ ((fiEnable && (1739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_4_io_in_control_0_propagate_b <=( _mesh_10_4_io_out_control_0_propagate) ^ ((fiEnable && (1740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_4_io_out_valid_0) begin
			b_140_0 <=( _mesh_11_4_io_out_b_0) ^ ((fiEnable && (1741 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1164_0 <=( _mesh_11_4_io_out_c_0) ^ ((fiEnable && (1742 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_4_io_in_control_0_shift_b <=( _mesh_11_4_io_out_control_0_shift) ^ ((fiEnable && (1743 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_4_io_in_control_0_dataflow_b <=( _mesh_11_4_io_out_control_0_dataflow) ^ ((fiEnable && (1744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_4_io_in_control_0_propagate_b <=( _mesh_11_4_io_out_control_0_propagate) ^ ((fiEnable && (1745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_4_io_out_valid_0) begin
			b_141_0 <=( _mesh_12_4_io_out_b_0) ^ ((fiEnable && (1746 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1165_0 <=( _mesh_12_4_io_out_c_0) ^ ((fiEnable && (1747 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_4_io_in_control_0_shift_b <=( _mesh_12_4_io_out_control_0_shift) ^ ((fiEnable && (1748 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_4_io_in_control_0_dataflow_b <=( _mesh_12_4_io_out_control_0_dataflow) ^ ((fiEnable && (1749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_4_io_in_control_0_propagate_b <=( _mesh_12_4_io_out_control_0_propagate) ^ ((fiEnable && (1750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_4_io_out_valid_0) begin
			b_142_0 <=( _mesh_13_4_io_out_b_0) ^ ((fiEnable && (1751 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1166_0 <=( _mesh_13_4_io_out_c_0) ^ ((fiEnable && (1752 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_4_io_in_control_0_shift_b <=( _mesh_13_4_io_out_control_0_shift) ^ ((fiEnable && (1753 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_4_io_in_control_0_dataflow_b <=( _mesh_13_4_io_out_control_0_dataflow) ^ ((fiEnable && (1754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_4_io_in_control_0_propagate_b <=( _mesh_13_4_io_out_control_0_propagate) ^ ((fiEnable && (1755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_4_io_out_valid_0) begin
			b_143_0 <=( _mesh_14_4_io_out_b_0) ^ ((fiEnable && (1756 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1167_0 <=( _mesh_14_4_io_out_c_0) ^ ((fiEnable && (1757 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_4_io_in_control_0_shift_b <=( _mesh_14_4_io_out_control_0_shift) ^ ((fiEnable && (1758 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_4_io_in_control_0_dataflow_b <=( _mesh_14_4_io_out_control_0_dataflow) ^ ((fiEnable && (1759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_4_io_in_control_0_propagate_b <=( _mesh_14_4_io_out_control_0_propagate) ^ ((fiEnable && (1760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_4_io_out_valid_0) begin
			b_144_0 <=( _mesh_15_4_io_out_b_0) ^ ((fiEnable && (1761 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1168_0 <=( _mesh_15_4_io_out_c_0) ^ ((fiEnable && (1762 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_4_io_in_control_0_shift_b <=( _mesh_15_4_io_out_control_0_shift) ^ ((fiEnable && (1763 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_4_io_in_control_0_dataflow_b <=( _mesh_15_4_io_out_control_0_dataflow) ^ ((fiEnable && (1764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_4_io_in_control_0_propagate_b <=( _mesh_15_4_io_out_control_0_propagate) ^ ((fiEnable && (1765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_4_io_out_valid_0) begin
			b_145_0 <=( _mesh_16_4_io_out_b_0) ^ ((fiEnable && (1766 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1169_0 <=( _mesh_16_4_io_out_c_0) ^ ((fiEnable && (1767 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_4_io_in_control_0_shift_b <=( _mesh_16_4_io_out_control_0_shift) ^ ((fiEnable && (1768 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_4_io_in_control_0_dataflow_b <=( _mesh_16_4_io_out_control_0_dataflow) ^ ((fiEnable && (1769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_4_io_in_control_0_propagate_b <=( _mesh_16_4_io_out_control_0_propagate) ^ ((fiEnable && (1770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_4_io_out_valid_0) begin
			b_146_0 <=( _mesh_17_4_io_out_b_0) ^ ((fiEnable && (1771 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1170_0 <=( _mesh_17_4_io_out_c_0) ^ ((fiEnable && (1772 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_4_io_in_control_0_shift_b <=( _mesh_17_4_io_out_control_0_shift) ^ ((fiEnable && (1773 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_4_io_in_control_0_dataflow_b <=( _mesh_17_4_io_out_control_0_dataflow) ^ ((fiEnable && (1774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_4_io_in_control_0_propagate_b <=( _mesh_17_4_io_out_control_0_propagate) ^ ((fiEnable && (1775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_4_io_out_valid_0) begin
			b_147_0 <=( _mesh_18_4_io_out_b_0) ^ ((fiEnable && (1776 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1171_0 <=( _mesh_18_4_io_out_c_0) ^ ((fiEnable && (1777 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_4_io_in_control_0_shift_b <=( _mesh_18_4_io_out_control_0_shift) ^ ((fiEnable && (1778 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_4_io_in_control_0_dataflow_b <=( _mesh_18_4_io_out_control_0_dataflow) ^ ((fiEnable && (1779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_4_io_in_control_0_propagate_b <=( _mesh_18_4_io_out_control_0_propagate) ^ ((fiEnable && (1780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_4_io_out_valid_0) begin
			b_148_0 <=( _mesh_19_4_io_out_b_0) ^ ((fiEnable && (1781 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1172_0 <=( _mesh_19_4_io_out_c_0) ^ ((fiEnable && (1782 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_4_io_in_control_0_shift_b <=( _mesh_19_4_io_out_control_0_shift) ^ ((fiEnable && (1783 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_4_io_in_control_0_dataflow_b <=( _mesh_19_4_io_out_control_0_dataflow) ^ ((fiEnable && (1784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_4_io_in_control_0_propagate_b <=( _mesh_19_4_io_out_control_0_propagate) ^ ((fiEnable && (1785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_4_io_out_valid_0) begin
			b_149_0 <=( _mesh_20_4_io_out_b_0) ^ ((fiEnable && (1786 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1173_0 <=( _mesh_20_4_io_out_c_0) ^ ((fiEnable && (1787 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_4_io_in_control_0_shift_b <=( _mesh_20_4_io_out_control_0_shift) ^ ((fiEnable && (1788 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_4_io_in_control_0_dataflow_b <=( _mesh_20_4_io_out_control_0_dataflow) ^ ((fiEnable && (1789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_4_io_in_control_0_propagate_b <=( _mesh_20_4_io_out_control_0_propagate) ^ ((fiEnable && (1790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_4_io_out_valid_0) begin
			b_150_0 <=( _mesh_21_4_io_out_b_0) ^ ((fiEnable && (1791 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1174_0 <=( _mesh_21_4_io_out_c_0) ^ ((fiEnable && (1792 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_4_io_in_control_0_shift_b <=( _mesh_21_4_io_out_control_0_shift) ^ ((fiEnable && (1793 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_4_io_in_control_0_dataflow_b <=( _mesh_21_4_io_out_control_0_dataflow) ^ ((fiEnable && (1794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_4_io_in_control_0_propagate_b <=( _mesh_21_4_io_out_control_0_propagate) ^ ((fiEnable && (1795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_4_io_out_valid_0) begin
			b_151_0 <=( _mesh_22_4_io_out_b_0) ^ ((fiEnable && (1796 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1175_0 <=( _mesh_22_4_io_out_c_0) ^ ((fiEnable && (1797 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_4_io_in_control_0_shift_b <=( _mesh_22_4_io_out_control_0_shift) ^ ((fiEnable && (1798 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_4_io_in_control_0_dataflow_b <=( _mesh_22_4_io_out_control_0_dataflow) ^ ((fiEnable && (1799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_4_io_in_control_0_propagate_b <=( _mesh_22_4_io_out_control_0_propagate) ^ ((fiEnable && (1800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_4_io_out_valid_0) begin
			b_152_0 <=( _mesh_23_4_io_out_b_0) ^ ((fiEnable && (1801 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1176_0 <=( _mesh_23_4_io_out_c_0) ^ ((fiEnable && (1802 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_4_io_in_control_0_shift_b <=( _mesh_23_4_io_out_control_0_shift) ^ ((fiEnable && (1803 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_4_io_in_control_0_dataflow_b <=( _mesh_23_4_io_out_control_0_dataflow) ^ ((fiEnable && (1804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_4_io_in_control_0_propagate_b <=( _mesh_23_4_io_out_control_0_propagate) ^ ((fiEnable && (1805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_4_io_out_valid_0) begin
			b_153_0 <=( _mesh_24_4_io_out_b_0) ^ ((fiEnable && (1806 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1177_0 <=( _mesh_24_4_io_out_c_0) ^ ((fiEnable && (1807 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_4_io_in_control_0_shift_b <=( _mesh_24_4_io_out_control_0_shift) ^ ((fiEnable && (1808 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_4_io_in_control_0_dataflow_b <=( _mesh_24_4_io_out_control_0_dataflow) ^ ((fiEnable && (1809 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_4_io_in_control_0_propagate_b <=( _mesh_24_4_io_out_control_0_propagate) ^ ((fiEnable && (1810 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_4_io_out_valid_0) begin
			b_154_0 <=( _mesh_25_4_io_out_b_0) ^ ((fiEnable && (1811 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1178_0 <=( _mesh_25_4_io_out_c_0) ^ ((fiEnable && (1812 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_4_io_in_control_0_shift_b <=( _mesh_25_4_io_out_control_0_shift) ^ ((fiEnable && (1813 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_4_io_in_control_0_dataflow_b <=( _mesh_25_4_io_out_control_0_dataflow) ^ ((fiEnable && (1814 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_4_io_in_control_0_propagate_b <=( _mesh_25_4_io_out_control_0_propagate) ^ ((fiEnable && (1815 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_4_io_out_valid_0) begin
			b_155_0 <=( _mesh_26_4_io_out_b_0) ^ ((fiEnable && (1816 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1179_0 <=( _mesh_26_4_io_out_c_0) ^ ((fiEnable && (1817 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_4_io_in_control_0_shift_b <=( _mesh_26_4_io_out_control_0_shift) ^ ((fiEnable && (1818 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_4_io_in_control_0_dataflow_b <=( _mesh_26_4_io_out_control_0_dataflow) ^ ((fiEnable && (1819 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_4_io_in_control_0_propagate_b <=( _mesh_26_4_io_out_control_0_propagate) ^ ((fiEnable && (1820 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_4_io_out_valid_0) begin
			b_156_0 <=( _mesh_27_4_io_out_b_0) ^ ((fiEnable && (1821 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1180_0 <=( _mesh_27_4_io_out_c_0) ^ ((fiEnable && (1822 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_4_io_in_control_0_shift_b <=( _mesh_27_4_io_out_control_0_shift) ^ ((fiEnable && (1823 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_4_io_in_control_0_dataflow_b <=( _mesh_27_4_io_out_control_0_dataflow) ^ ((fiEnable && (1824 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_4_io_in_control_0_propagate_b <=( _mesh_27_4_io_out_control_0_propagate) ^ ((fiEnable && (1825 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_4_io_out_valid_0) begin
			b_157_0 <=( _mesh_28_4_io_out_b_0) ^ ((fiEnable && (1826 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1181_0 <=( _mesh_28_4_io_out_c_0) ^ ((fiEnable && (1827 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_4_io_in_control_0_shift_b <=( _mesh_28_4_io_out_control_0_shift) ^ ((fiEnable && (1828 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_4_io_in_control_0_dataflow_b <=( _mesh_28_4_io_out_control_0_dataflow) ^ ((fiEnable && (1829 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_4_io_in_control_0_propagate_b <=( _mesh_28_4_io_out_control_0_propagate) ^ ((fiEnable && (1830 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_4_io_out_valid_0) begin
			b_158_0 <=( _mesh_29_4_io_out_b_0) ^ ((fiEnable && (1831 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1182_0 <=( _mesh_29_4_io_out_c_0) ^ ((fiEnable && (1832 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_4_io_in_control_0_shift_b <=( _mesh_29_4_io_out_control_0_shift) ^ ((fiEnable && (1833 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_4_io_in_control_0_dataflow_b <=( _mesh_29_4_io_out_control_0_dataflow) ^ ((fiEnable && (1834 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_4_io_in_control_0_propagate_b <=( _mesh_29_4_io_out_control_0_propagate) ^ ((fiEnable && (1835 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_4_io_out_valid_0) begin
			b_159_0 <=( _mesh_30_4_io_out_b_0) ^ ((fiEnable && (1836 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1183_0 <=( _mesh_30_4_io_out_c_0) ^ ((fiEnable && (1837 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_4_io_in_control_0_shift_b <=( _mesh_30_4_io_out_control_0_shift) ^ ((fiEnable && (1838 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_4_io_in_control_0_dataflow_b <=( _mesh_30_4_io_out_control_0_dataflow) ^ ((fiEnable && (1839 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_4_io_in_control_0_propagate_b <=( _mesh_30_4_io_out_control_0_propagate) ^ ((fiEnable && (1840 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_5_0) begin
			b_160_0 <=( io_in_b_5_0) ^ ((fiEnable && (1841 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1184_0 <=( io_in_d_5_0) ^ ((fiEnable && (1842 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_5_io_in_control_0_shift_b <=( io_in_control_5_0_shift) ^ ((fiEnable && (1843 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_5_io_in_control_0_dataflow_b <=( io_in_control_5_0_dataflow) ^ ((fiEnable && (1844 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_5_io_in_control_0_propagate_b <=( io_in_control_5_0_propagate) ^ ((fiEnable && (1845 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_5_io_out_valid_0) begin
			b_161_0 <=( _mesh_0_5_io_out_b_0) ^ ((fiEnable && (1846 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1185_0 <=( _mesh_0_5_io_out_c_0) ^ ((fiEnable && (1847 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_5_io_in_control_0_shift_b <=( _mesh_0_5_io_out_control_0_shift) ^ ((fiEnable && (1848 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_5_io_in_control_0_dataflow_b <=( _mesh_0_5_io_out_control_0_dataflow) ^ ((fiEnable && (1849 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_5_io_in_control_0_propagate_b <=( _mesh_0_5_io_out_control_0_propagate) ^ ((fiEnable && (1850 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_5_io_out_valid_0) begin
			b_162_0 <=( _mesh_1_5_io_out_b_0) ^ ((fiEnable && (1851 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1186_0 <=( _mesh_1_5_io_out_c_0) ^ ((fiEnable && (1852 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_5_io_in_control_0_shift_b <=( _mesh_1_5_io_out_control_0_shift) ^ ((fiEnable && (1853 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_5_io_in_control_0_dataflow_b <=( _mesh_1_5_io_out_control_0_dataflow) ^ ((fiEnable && (1854 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_5_io_in_control_0_propagate_b <=( _mesh_1_5_io_out_control_0_propagate) ^ ((fiEnable && (1855 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_5_io_out_valid_0) begin
			b_163_0 <=( _mesh_2_5_io_out_b_0) ^ ((fiEnable && (1856 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1187_0 <=( _mesh_2_5_io_out_c_0) ^ ((fiEnable && (1857 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_5_io_in_control_0_shift_b <=( _mesh_2_5_io_out_control_0_shift) ^ ((fiEnable && (1858 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_5_io_in_control_0_dataflow_b <=( _mesh_2_5_io_out_control_0_dataflow) ^ ((fiEnable && (1859 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_5_io_in_control_0_propagate_b <=( _mesh_2_5_io_out_control_0_propagate) ^ ((fiEnable && (1860 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_5_io_out_valid_0) begin
			b_164_0 <=( _mesh_3_5_io_out_b_0) ^ ((fiEnable && (1861 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1188_0 <=( _mesh_3_5_io_out_c_0) ^ ((fiEnable && (1862 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_5_io_in_control_0_shift_b <=( _mesh_3_5_io_out_control_0_shift) ^ ((fiEnable && (1863 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_5_io_in_control_0_dataflow_b <=( _mesh_3_5_io_out_control_0_dataflow) ^ ((fiEnable && (1864 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_5_io_in_control_0_propagate_b <=( _mesh_3_5_io_out_control_0_propagate) ^ ((fiEnable && (1865 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_5_io_out_valid_0) begin
			b_165_0 <=( _mesh_4_5_io_out_b_0) ^ ((fiEnable && (1866 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1189_0 <=( _mesh_4_5_io_out_c_0) ^ ((fiEnable && (1867 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_5_io_in_control_0_shift_b <=( _mesh_4_5_io_out_control_0_shift) ^ ((fiEnable && (1868 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_5_io_in_control_0_dataflow_b <=( _mesh_4_5_io_out_control_0_dataflow) ^ ((fiEnable && (1869 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_5_io_in_control_0_propagate_b <=( _mesh_4_5_io_out_control_0_propagate) ^ ((fiEnable && (1870 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_5_io_out_valid_0) begin
			b_166_0 <=( _mesh_5_5_io_out_b_0) ^ ((fiEnable && (1871 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1190_0 <=( _mesh_5_5_io_out_c_0) ^ ((fiEnable && (1872 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_5_io_in_control_0_shift_b <=( _mesh_5_5_io_out_control_0_shift) ^ ((fiEnable && (1873 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_5_io_in_control_0_dataflow_b <=( _mesh_5_5_io_out_control_0_dataflow) ^ ((fiEnable && (1874 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_5_io_in_control_0_propagate_b <=( _mesh_5_5_io_out_control_0_propagate) ^ ((fiEnable && (1875 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_5_io_out_valid_0) begin
			b_167_0 <=( _mesh_6_5_io_out_b_0) ^ ((fiEnable && (1876 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1191_0 <=( _mesh_6_5_io_out_c_0) ^ ((fiEnable && (1877 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_5_io_in_control_0_shift_b <=( _mesh_6_5_io_out_control_0_shift) ^ ((fiEnable && (1878 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_5_io_in_control_0_dataflow_b <=( _mesh_6_5_io_out_control_0_dataflow) ^ ((fiEnable && (1879 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_5_io_in_control_0_propagate_b <=( _mesh_6_5_io_out_control_0_propagate) ^ ((fiEnable && (1880 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_5_io_out_valid_0) begin
			b_168_0 <=( _mesh_7_5_io_out_b_0) ^ ((fiEnable && (1881 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1192_0 <=( _mesh_7_5_io_out_c_0) ^ ((fiEnable && (1882 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_5_io_in_control_0_shift_b <=( _mesh_7_5_io_out_control_0_shift) ^ ((fiEnable && (1883 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_5_io_in_control_0_dataflow_b <=( _mesh_7_5_io_out_control_0_dataflow) ^ ((fiEnable && (1884 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_5_io_in_control_0_propagate_b <=( _mesh_7_5_io_out_control_0_propagate) ^ ((fiEnable && (1885 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_5_io_out_valid_0) begin
			b_169_0 <=( _mesh_8_5_io_out_b_0) ^ ((fiEnable && (1886 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1193_0 <=( _mesh_8_5_io_out_c_0) ^ ((fiEnable && (1887 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_5_io_in_control_0_shift_b <=( _mesh_8_5_io_out_control_0_shift) ^ ((fiEnable && (1888 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_5_io_in_control_0_dataflow_b <=( _mesh_8_5_io_out_control_0_dataflow) ^ ((fiEnable && (1889 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_5_io_in_control_0_propagate_b <=( _mesh_8_5_io_out_control_0_propagate) ^ ((fiEnable && (1890 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_5_io_out_valid_0) begin
			b_170_0 <=( _mesh_9_5_io_out_b_0) ^ ((fiEnable && (1891 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1194_0 <=( _mesh_9_5_io_out_c_0) ^ ((fiEnable && (1892 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_5_io_in_control_0_shift_b <=( _mesh_9_5_io_out_control_0_shift) ^ ((fiEnable && (1893 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_5_io_in_control_0_dataflow_b <=( _mesh_9_5_io_out_control_0_dataflow) ^ ((fiEnable && (1894 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_5_io_in_control_0_propagate_b <=( _mesh_9_5_io_out_control_0_propagate) ^ ((fiEnable && (1895 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_5_io_out_valid_0) begin
			b_171_0 <=( _mesh_10_5_io_out_b_0) ^ ((fiEnable && (1896 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1195_0 <=( _mesh_10_5_io_out_c_0) ^ ((fiEnable && (1897 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_5_io_in_control_0_shift_b <=( _mesh_10_5_io_out_control_0_shift) ^ ((fiEnable && (1898 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_5_io_in_control_0_dataflow_b <=( _mesh_10_5_io_out_control_0_dataflow) ^ ((fiEnable && (1899 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_5_io_in_control_0_propagate_b <=( _mesh_10_5_io_out_control_0_propagate) ^ ((fiEnable && (1900 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_5_io_out_valid_0) begin
			b_172_0 <=( _mesh_11_5_io_out_b_0) ^ ((fiEnable && (1901 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1196_0 <=( _mesh_11_5_io_out_c_0) ^ ((fiEnable && (1902 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_5_io_in_control_0_shift_b <=( _mesh_11_5_io_out_control_0_shift) ^ ((fiEnable && (1903 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_5_io_in_control_0_dataflow_b <=( _mesh_11_5_io_out_control_0_dataflow) ^ ((fiEnable && (1904 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_5_io_in_control_0_propagate_b <=( _mesh_11_5_io_out_control_0_propagate) ^ ((fiEnable && (1905 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_5_io_out_valid_0) begin
			b_173_0 <=( _mesh_12_5_io_out_b_0) ^ ((fiEnable && (1906 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1197_0 <=( _mesh_12_5_io_out_c_0) ^ ((fiEnable && (1907 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_5_io_in_control_0_shift_b <=( _mesh_12_5_io_out_control_0_shift) ^ ((fiEnable && (1908 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_5_io_in_control_0_dataflow_b <=( _mesh_12_5_io_out_control_0_dataflow) ^ ((fiEnable && (1909 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_5_io_in_control_0_propagate_b <=( _mesh_12_5_io_out_control_0_propagate) ^ ((fiEnable && (1910 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_5_io_out_valid_0) begin
			b_174_0 <=( _mesh_13_5_io_out_b_0) ^ ((fiEnable && (1911 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1198_0 <=( _mesh_13_5_io_out_c_0) ^ ((fiEnable && (1912 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_5_io_in_control_0_shift_b <=( _mesh_13_5_io_out_control_0_shift) ^ ((fiEnable && (1913 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_5_io_in_control_0_dataflow_b <=( _mesh_13_5_io_out_control_0_dataflow) ^ ((fiEnable && (1914 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_5_io_in_control_0_propagate_b <=( _mesh_13_5_io_out_control_0_propagate) ^ ((fiEnable && (1915 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_5_io_out_valid_0) begin
			b_175_0 <=( _mesh_14_5_io_out_b_0) ^ ((fiEnable && (1916 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1199_0 <=( _mesh_14_5_io_out_c_0) ^ ((fiEnable && (1917 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_5_io_in_control_0_shift_b <=( _mesh_14_5_io_out_control_0_shift) ^ ((fiEnable && (1918 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_5_io_in_control_0_dataflow_b <=( _mesh_14_5_io_out_control_0_dataflow) ^ ((fiEnable && (1919 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_5_io_in_control_0_propagate_b <=( _mesh_14_5_io_out_control_0_propagate) ^ ((fiEnable && (1920 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_5_io_out_valid_0) begin
			b_176_0 <=( _mesh_15_5_io_out_b_0) ^ ((fiEnable && (1921 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1200_0 <=( _mesh_15_5_io_out_c_0) ^ ((fiEnable && (1922 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_5_io_in_control_0_shift_b <=( _mesh_15_5_io_out_control_0_shift) ^ ((fiEnable && (1923 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_5_io_in_control_0_dataflow_b <=( _mesh_15_5_io_out_control_0_dataflow) ^ ((fiEnable && (1924 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_5_io_in_control_0_propagate_b <=( _mesh_15_5_io_out_control_0_propagate) ^ ((fiEnable && (1925 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_5_io_out_valid_0) begin
			b_177_0 <=( _mesh_16_5_io_out_b_0) ^ ((fiEnable && (1926 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1201_0 <=( _mesh_16_5_io_out_c_0) ^ ((fiEnable && (1927 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_5_io_in_control_0_shift_b <=( _mesh_16_5_io_out_control_0_shift) ^ ((fiEnable && (1928 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_5_io_in_control_0_dataflow_b <=( _mesh_16_5_io_out_control_0_dataflow) ^ ((fiEnable && (1929 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_5_io_in_control_0_propagate_b <=( _mesh_16_5_io_out_control_0_propagate) ^ ((fiEnable && (1930 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_5_io_out_valid_0) begin
			b_178_0 <=( _mesh_17_5_io_out_b_0) ^ ((fiEnable && (1931 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1202_0 <=( _mesh_17_5_io_out_c_0) ^ ((fiEnable && (1932 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_5_io_in_control_0_shift_b <=( _mesh_17_5_io_out_control_0_shift) ^ ((fiEnable && (1933 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_5_io_in_control_0_dataflow_b <=( _mesh_17_5_io_out_control_0_dataflow) ^ ((fiEnable && (1934 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_5_io_in_control_0_propagate_b <=( _mesh_17_5_io_out_control_0_propagate) ^ ((fiEnable && (1935 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_5_io_out_valid_0) begin
			b_179_0 <=( _mesh_18_5_io_out_b_0) ^ ((fiEnable && (1936 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1203_0 <=( _mesh_18_5_io_out_c_0) ^ ((fiEnable && (1937 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_5_io_in_control_0_shift_b <=( _mesh_18_5_io_out_control_0_shift) ^ ((fiEnable && (1938 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_5_io_in_control_0_dataflow_b <=( _mesh_18_5_io_out_control_0_dataflow) ^ ((fiEnable && (1939 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_5_io_in_control_0_propagate_b <=( _mesh_18_5_io_out_control_0_propagate) ^ ((fiEnable && (1940 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_5_io_out_valid_0) begin
			b_180_0 <=( _mesh_19_5_io_out_b_0) ^ ((fiEnable && (1941 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1204_0 <=( _mesh_19_5_io_out_c_0) ^ ((fiEnable && (1942 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_5_io_in_control_0_shift_b <=( _mesh_19_5_io_out_control_0_shift) ^ ((fiEnable && (1943 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_5_io_in_control_0_dataflow_b <=( _mesh_19_5_io_out_control_0_dataflow) ^ ((fiEnable && (1944 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_5_io_in_control_0_propagate_b <=( _mesh_19_5_io_out_control_0_propagate) ^ ((fiEnable && (1945 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_5_io_out_valid_0) begin
			b_181_0 <=( _mesh_20_5_io_out_b_0) ^ ((fiEnable && (1946 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1205_0 <=( _mesh_20_5_io_out_c_0) ^ ((fiEnable && (1947 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_5_io_in_control_0_shift_b <=( _mesh_20_5_io_out_control_0_shift) ^ ((fiEnable && (1948 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_5_io_in_control_0_dataflow_b <=( _mesh_20_5_io_out_control_0_dataflow) ^ ((fiEnable && (1949 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_5_io_in_control_0_propagate_b <=( _mesh_20_5_io_out_control_0_propagate) ^ ((fiEnable && (1950 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_5_io_out_valid_0) begin
			b_182_0 <=( _mesh_21_5_io_out_b_0) ^ ((fiEnable && (1951 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1206_0 <=( _mesh_21_5_io_out_c_0) ^ ((fiEnable && (1952 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_5_io_in_control_0_shift_b <=( _mesh_21_5_io_out_control_0_shift) ^ ((fiEnable && (1953 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_5_io_in_control_0_dataflow_b <=( _mesh_21_5_io_out_control_0_dataflow) ^ ((fiEnable && (1954 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_5_io_in_control_0_propagate_b <=( _mesh_21_5_io_out_control_0_propagate) ^ ((fiEnable && (1955 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_5_io_out_valid_0) begin
			b_183_0 <=( _mesh_22_5_io_out_b_0) ^ ((fiEnable && (1956 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1207_0 <=( _mesh_22_5_io_out_c_0) ^ ((fiEnable && (1957 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_5_io_in_control_0_shift_b <=( _mesh_22_5_io_out_control_0_shift) ^ ((fiEnable && (1958 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_5_io_in_control_0_dataflow_b <=( _mesh_22_5_io_out_control_0_dataflow) ^ ((fiEnable && (1959 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_5_io_in_control_0_propagate_b <=( _mesh_22_5_io_out_control_0_propagate) ^ ((fiEnable && (1960 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_5_io_out_valid_0) begin
			b_184_0 <=( _mesh_23_5_io_out_b_0) ^ ((fiEnable && (1961 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1208_0 <=( _mesh_23_5_io_out_c_0) ^ ((fiEnable && (1962 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_5_io_in_control_0_shift_b <=( _mesh_23_5_io_out_control_0_shift) ^ ((fiEnable && (1963 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_5_io_in_control_0_dataflow_b <=( _mesh_23_5_io_out_control_0_dataflow) ^ ((fiEnable && (1964 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_5_io_in_control_0_propagate_b <=( _mesh_23_5_io_out_control_0_propagate) ^ ((fiEnable && (1965 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_5_io_out_valid_0) begin
			b_185_0 <=( _mesh_24_5_io_out_b_0) ^ ((fiEnable && (1966 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1209_0 <=( _mesh_24_5_io_out_c_0) ^ ((fiEnable && (1967 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_5_io_in_control_0_shift_b <=( _mesh_24_5_io_out_control_0_shift) ^ ((fiEnable && (1968 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_5_io_in_control_0_dataflow_b <=( _mesh_24_5_io_out_control_0_dataflow) ^ ((fiEnable && (1969 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_5_io_in_control_0_propagate_b <=( _mesh_24_5_io_out_control_0_propagate) ^ ((fiEnable && (1970 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_5_io_out_valid_0) begin
			b_186_0 <=( _mesh_25_5_io_out_b_0) ^ ((fiEnable && (1971 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1210_0 <=( _mesh_25_5_io_out_c_0) ^ ((fiEnable && (1972 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_5_io_in_control_0_shift_b <=( _mesh_25_5_io_out_control_0_shift) ^ ((fiEnable && (1973 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_5_io_in_control_0_dataflow_b <=( _mesh_25_5_io_out_control_0_dataflow) ^ ((fiEnable && (1974 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_5_io_in_control_0_propagate_b <=( _mesh_25_5_io_out_control_0_propagate) ^ ((fiEnable && (1975 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_5_io_out_valid_0) begin
			b_187_0 <=( _mesh_26_5_io_out_b_0) ^ ((fiEnable && (1976 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1211_0 <=( _mesh_26_5_io_out_c_0) ^ ((fiEnable && (1977 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_5_io_in_control_0_shift_b <=( _mesh_26_5_io_out_control_0_shift) ^ ((fiEnable && (1978 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_5_io_in_control_0_dataflow_b <=( _mesh_26_5_io_out_control_0_dataflow) ^ ((fiEnable && (1979 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_5_io_in_control_0_propagate_b <=( _mesh_26_5_io_out_control_0_propagate) ^ ((fiEnable && (1980 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_5_io_out_valid_0) begin
			b_188_0 <=( _mesh_27_5_io_out_b_0) ^ ((fiEnable && (1981 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1212_0 <=( _mesh_27_5_io_out_c_0) ^ ((fiEnable && (1982 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_5_io_in_control_0_shift_b <=( _mesh_27_5_io_out_control_0_shift) ^ ((fiEnable && (1983 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_5_io_in_control_0_dataflow_b <=( _mesh_27_5_io_out_control_0_dataflow) ^ ((fiEnable && (1984 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_5_io_in_control_0_propagate_b <=( _mesh_27_5_io_out_control_0_propagate) ^ ((fiEnable && (1985 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_5_io_out_valid_0) begin
			b_189_0 <=( _mesh_28_5_io_out_b_0) ^ ((fiEnable && (1986 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1213_0 <=( _mesh_28_5_io_out_c_0) ^ ((fiEnable && (1987 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_5_io_in_control_0_shift_b <=( _mesh_28_5_io_out_control_0_shift) ^ ((fiEnable && (1988 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_5_io_in_control_0_dataflow_b <=( _mesh_28_5_io_out_control_0_dataflow) ^ ((fiEnable && (1989 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_5_io_in_control_0_propagate_b <=( _mesh_28_5_io_out_control_0_propagate) ^ ((fiEnable && (1990 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_5_io_out_valid_0) begin
			b_190_0 <=( _mesh_29_5_io_out_b_0) ^ ((fiEnable && (1991 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1214_0 <=( _mesh_29_5_io_out_c_0) ^ ((fiEnable && (1992 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_5_io_in_control_0_shift_b <=( _mesh_29_5_io_out_control_0_shift) ^ ((fiEnable && (1993 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_5_io_in_control_0_dataflow_b <=( _mesh_29_5_io_out_control_0_dataflow) ^ ((fiEnable && (1994 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_5_io_in_control_0_propagate_b <=( _mesh_29_5_io_out_control_0_propagate) ^ ((fiEnable && (1995 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_5_io_out_valid_0) begin
			b_191_0 <=( _mesh_30_5_io_out_b_0) ^ ((fiEnable && (1996 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1215_0 <=( _mesh_30_5_io_out_c_0) ^ ((fiEnable && (1997 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_5_io_in_control_0_shift_b <=( _mesh_30_5_io_out_control_0_shift) ^ ((fiEnable && (1998 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_5_io_in_control_0_dataflow_b <=( _mesh_30_5_io_out_control_0_dataflow) ^ ((fiEnable && (1999 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_5_io_in_control_0_propagate_b <=( _mesh_30_5_io_out_control_0_propagate) ^ ((fiEnable && (2000 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_6_0) begin
			b_192_0 <=( io_in_b_6_0) ^ ((fiEnable && (2001 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1216_0 <=( io_in_d_6_0) ^ ((fiEnable && (2002 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_6_io_in_control_0_shift_b <=( io_in_control_6_0_shift) ^ ((fiEnable && (2003 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_6_io_in_control_0_dataflow_b <=( io_in_control_6_0_dataflow) ^ ((fiEnable && (2004 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_6_io_in_control_0_propagate_b <=( io_in_control_6_0_propagate) ^ ((fiEnable && (2005 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_6_io_out_valid_0) begin
			b_193_0 <=( _mesh_0_6_io_out_b_0) ^ ((fiEnable && (2006 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1217_0 <=( _mesh_0_6_io_out_c_0) ^ ((fiEnable && (2007 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_6_io_in_control_0_shift_b <=( _mesh_0_6_io_out_control_0_shift) ^ ((fiEnable && (2008 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_6_io_in_control_0_dataflow_b <=( _mesh_0_6_io_out_control_0_dataflow) ^ ((fiEnable && (2009 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_6_io_in_control_0_propagate_b <=( _mesh_0_6_io_out_control_0_propagate) ^ ((fiEnable && (2010 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_6_io_out_valid_0) begin
			b_194_0 <=( _mesh_1_6_io_out_b_0) ^ ((fiEnable && (2011 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1218_0 <=( _mesh_1_6_io_out_c_0) ^ ((fiEnable && (2012 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_6_io_in_control_0_shift_b <=( _mesh_1_6_io_out_control_0_shift) ^ ((fiEnable && (2013 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_6_io_in_control_0_dataflow_b <=( _mesh_1_6_io_out_control_0_dataflow) ^ ((fiEnable && (2014 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_6_io_in_control_0_propagate_b <=( _mesh_1_6_io_out_control_0_propagate) ^ ((fiEnable && (2015 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_6_io_out_valid_0) begin
			b_195_0 <=( _mesh_2_6_io_out_b_0) ^ ((fiEnable && (2016 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1219_0 <=( _mesh_2_6_io_out_c_0) ^ ((fiEnable && (2017 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_6_io_in_control_0_shift_b <=( _mesh_2_6_io_out_control_0_shift) ^ ((fiEnable && (2018 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_6_io_in_control_0_dataflow_b <=( _mesh_2_6_io_out_control_0_dataflow) ^ ((fiEnable && (2019 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_6_io_in_control_0_propagate_b <=( _mesh_2_6_io_out_control_0_propagate) ^ ((fiEnable && (2020 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_6_io_out_valid_0) begin
			b_196_0 <=( _mesh_3_6_io_out_b_0) ^ ((fiEnable && (2021 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1220_0 <=( _mesh_3_6_io_out_c_0) ^ ((fiEnable && (2022 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_6_io_in_control_0_shift_b <=( _mesh_3_6_io_out_control_0_shift) ^ ((fiEnable && (2023 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_6_io_in_control_0_dataflow_b <=( _mesh_3_6_io_out_control_0_dataflow) ^ ((fiEnable && (2024 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_6_io_in_control_0_propagate_b <=( _mesh_3_6_io_out_control_0_propagate) ^ ((fiEnable && (2025 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_6_io_out_valid_0) begin
			b_197_0 <=( _mesh_4_6_io_out_b_0) ^ ((fiEnable && (2026 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1221_0 <=( _mesh_4_6_io_out_c_0) ^ ((fiEnable && (2027 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_6_io_in_control_0_shift_b <=( _mesh_4_6_io_out_control_0_shift) ^ ((fiEnable && (2028 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_6_io_in_control_0_dataflow_b <=( _mesh_4_6_io_out_control_0_dataflow) ^ ((fiEnable && (2029 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_6_io_in_control_0_propagate_b <=( _mesh_4_6_io_out_control_0_propagate) ^ ((fiEnable && (2030 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_6_io_out_valid_0) begin
			b_198_0 <=( _mesh_5_6_io_out_b_0) ^ ((fiEnable && (2031 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1222_0 <=( _mesh_5_6_io_out_c_0) ^ ((fiEnable && (2032 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_6_io_in_control_0_shift_b <=( _mesh_5_6_io_out_control_0_shift) ^ ((fiEnable && (2033 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_6_io_in_control_0_dataflow_b <=( _mesh_5_6_io_out_control_0_dataflow) ^ ((fiEnable && (2034 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_6_io_in_control_0_propagate_b <=( _mesh_5_6_io_out_control_0_propagate) ^ ((fiEnable && (2035 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_6_io_out_valid_0) begin
			b_199_0 <=( _mesh_6_6_io_out_b_0) ^ ((fiEnable && (2036 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1223_0 <=( _mesh_6_6_io_out_c_0) ^ ((fiEnable && (2037 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_6_io_in_control_0_shift_b <=( _mesh_6_6_io_out_control_0_shift) ^ ((fiEnable && (2038 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_6_io_in_control_0_dataflow_b <=( _mesh_6_6_io_out_control_0_dataflow) ^ ((fiEnable && (2039 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_6_io_in_control_0_propagate_b <=( _mesh_6_6_io_out_control_0_propagate) ^ ((fiEnable && (2040 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_6_io_out_valid_0) begin
			b_200_0 <=( _mesh_7_6_io_out_b_0) ^ ((fiEnable && (2041 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1224_0 <=( _mesh_7_6_io_out_c_0) ^ ((fiEnable && (2042 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_6_io_in_control_0_shift_b <=( _mesh_7_6_io_out_control_0_shift) ^ ((fiEnable && (2043 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_6_io_in_control_0_dataflow_b <=( _mesh_7_6_io_out_control_0_dataflow) ^ ((fiEnable && (2044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_6_io_in_control_0_propagate_b <=( _mesh_7_6_io_out_control_0_propagate) ^ ((fiEnable && (2045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_6_io_out_valid_0) begin
			b_201_0 <=( _mesh_8_6_io_out_b_0) ^ ((fiEnable && (2046 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1225_0 <=( _mesh_8_6_io_out_c_0) ^ ((fiEnable && (2047 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_6_io_in_control_0_shift_b <=( _mesh_8_6_io_out_control_0_shift) ^ ((fiEnable && (2048 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_6_io_in_control_0_dataflow_b <=( _mesh_8_6_io_out_control_0_dataflow) ^ ((fiEnable && (2049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_6_io_in_control_0_propagate_b <=( _mesh_8_6_io_out_control_0_propagate) ^ ((fiEnable && (2050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_6_io_out_valid_0) begin
			b_202_0 <=( _mesh_9_6_io_out_b_0) ^ ((fiEnable && (2051 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1226_0 <=( _mesh_9_6_io_out_c_0) ^ ((fiEnable && (2052 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_6_io_in_control_0_shift_b <=( _mesh_9_6_io_out_control_0_shift) ^ ((fiEnable && (2053 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_6_io_in_control_0_dataflow_b <=( _mesh_9_6_io_out_control_0_dataflow) ^ ((fiEnable && (2054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_6_io_in_control_0_propagate_b <=( _mesh_9_6_io_out_control_0_propagate) ^ ((fiEnable && (2055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_6_io_out_valid_0) begin
			b_203_0 <=( _mesh_10_6_io_out_b_0) ^ ((fiEnable && (2056 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1227_0 <=( _mesh_10_6_io_out_c_0) ^ ((fiEnable && (2057 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_6_io_in_control_0_shift_b <=( _mesh_10_6_io_out_control_0_shift) ^ ((fiEnable && (2058 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_6_io_in_control_0_dataflow_b <=( _mesh_10_6_io_out_control_0_dataflow) ^ ((fiEnable && (2059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_6_io_in_control_0_propagate_b <=( _mesh_10_6_io_out_control_0_propagate) ^ ((fiEnable && (2060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_6_io_out_valid_0) begin
			b_204_0 <=( _mesh_11_6_io_out_b_0) ^ ((fiEnable && (2061 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1228_0 <=( _mesh_11_6_io_out_c_0) ^ ((fiEnable && (2062 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_6_io_in_control_0_shift_b <=( _mesh_11_6_io_out_control_0_shift) ^ ((fiEnable && (2063 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_6_io_in_control_0_dataflow_b <=( _mesh_11_6_io_out_control_0_dataflow) ^ ((fiEnable && (2064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_6_io_in_control_0_propagate_b <=( _mesh_11_6_io_out_control_0_propagate) ^ ((fiEnable && (2065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_6_io_out_valid_0) begin
			b_205_0 <=( _mesh_12_6_io_out_b_0) ^ ((fiEnable && (2066 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1229_0 <=( _mesh_12_6_io_out_c_0) ^ ((fiEnable && (2067 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_6_io_in_control_0_shift_b <=( _mesh_12_6_io_out_control_0_shift) ^ ((fiEnable && (2068 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_6_io_in_control_0_dataflow_b <=( _mesh_12_6_io_out_control_0_dataflow) ^ ((fiEnable && (2069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_6_io_in_control_0_propagate_b <=( _mesh_12_6_io_out_control_0_propagate) ^ ((fiEnable && (2070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_6_io_out_valid_0) begin
			b_206_0 <=( _mesh_13_6_io_out_b_0) ^ ((fiEnable && (2071 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1230_0 <=( _mesh_13_6_io_out_c_0) ^ ((fiEnable && (2072 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_6_io_in_control_0_shift_b <=( _mesh_13_6_io_out_control_0_shift) ^ ((fiEnable && (2073 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_6_io_in_control_0_dataflow_b <=( _mesh_13_6_io_out_control_0_dataflow) ^ ((fiEnable && (2074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_6_io_in_control_0_propagate_b <=( _mesh_13_6_io_out_control_0_propagate) ^ ((fiEnable && (2075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_6_io_out_valid_0) begin
			b_207_0 <=( _mesh_14_6_io_out_b_0) ^ ((fiEnable && (2076 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1231_0 <=( _mesh_14_6_io_out_c_0) ^ ((fiEnable && (2077 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_6_io_in_control_0_shift_b <=( _mesh_14_6_io_out_control_0_shift) ^ ((fiEnable && (2078 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_6_io_in_control_0_dataflow_b <=( _mesh_14_6_io_out_control_0_dataflow) ^ ((fiEnable && (2079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_6_io_in_control_0_propagate_b <=( _mesh_14_6_io_out_control_0_propagate) ^ ((fiEnable && (2080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_6_io_out_valid_0) begin
			b_208_0 <=( _mesh_15_6_io_out_b_0) ^ ((fiEnable && (2081 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1232_0 <=( _mesh_15_6_io_out_c_0) ^ ((fiEnable && (2082 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_6_io_in_control_0_shift_b <=( _mesh_15_6_io_out_control_0_shift) ^ ((fiEnable && (2083 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_6_io_in_control_0_dataflow_b <=( _mesh_15_6_io_out_control_0_dataflow) ^ ((fiEnable && (2084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_6_io_in_control_0_propagate_b <=( _mesh_15_6_io_out_control_0_propagate) ^ ((fiEnable && (2085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_6_io_out_valid_0) begin
			b_209_0 <=( _mesh_16_6_io_out_b_0) ^ ((fiEnable && (2086 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1233_0 <=( _mesh_16_6_io_out_c_0) ^ ((fiEnable && (2087 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_6_io_in_control_0_shift_b <=( _mesh_16_6_io_out_control_0_shift) ^ ((fiEnable && (2088 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_6_io_in_control_0_dataflow_b <=( _mesh_16_6_io_out_control_0_dataflow) ^ ((fiEnable && (2089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_6_io_in_control_0_propagate_b <=( _mesh_16_6_io_out_control_0_propagate) ^ ((fiEnable && (2090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_6_io_out_valid_0) begin
			b_210_0 <=( _mesh_17_6_io_out_b_0) ^ ((fiEnable && (2091 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1234_0 <=( _mesh_17_6_io_out_c_0) ^ ((fiEnable && (2092 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_6_io_in_control_0_shift_b <=( _mesh_17_6_io_out_control_0_shift) ^ ((fiEnable && (2093 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_6_io_in_control_0_dataflow_b <=( _mesh_17_6_io_out_control_0_dataflow) ^ ((fiEnable && (2094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_6_io_in_control_0_propagate_b <=( _mesh_17_6_io_out_control_0_propagate) ^ ((fiEnable && (2095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_6_io_out_valid_0) begin
			b_211_0 <=( _mesh_18_6_io_out_b_0) ^ ((fiEnable && (2096 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1235_0 <=( _mesh_18_6_io_out_c_0) ^ ((fiEnable && (2097 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_6_io_in_control_0_shift_b <=( _mesh_18_6_io_out_control_0_shift) ^ ((fiEnable && (2098 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_6_io_in_control_0_dataflow_b <=( _mesh_18_6_io_out_control_0_dataflow) ^ ((fiEnable && (2099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_6_io_in_control_0_propagate_b <=( _mesh_18_6_io_out_control_0_propagate) ^ ((fiEnable && (2100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_6_io_out_valid_0) begin
			b_212_0 <=( _mesh_19_6_io_out_b_0) ^ ((fiEnable && (2101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1236_0 <=( _mesh_19_6_io_out_c_0) ^ ((fiEnable && (2102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_6_io_in_control_0_shift_b <=( _mesh_19_6_io_out_control_0_shift) ^ ((fiEnable && (2103 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_6_io_in_control_0_dataflow_b <=( _mesh_19_6_io_out_control_0_dataflow) ^ ((fiEnable && (2104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_6_io_in_control_0_propagate_b <=( _mesh_19_6_io_out_control_0_propagate) ^ ((fiEnable && (2105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_6_io_out_valid_0) begin
			b_213_0 <=( _mesh_20_6_io_out_b_0) ^ ((fiEnable && (2106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1237_0 <=( _mesh_20_6_io_out_c_0) ^ ((fiEnable && (2107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_6_io_in_control_0_shift_b <=( _mesh_20_6_io_out_control_0_shift) ^ ((fiEnable && (2108 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_6_io_in_control_0_dataflow_b <=( _mesh_20_6_io_out_control_0_dataflow) ^ ((fiEnable && (2109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_6_io_in_control_0_propagate_b <=( _mesh_20_6_io_out_control_0_propagate) ^ ((fiEnable && (2110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_6_io_out_valid_0) begin
			b_214_0 <=( _mesh_21_6_io_out_b_0) ^ ((fiEnable && (2111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1238_0 <=( _mesh_21_6_io_out_c_0) ^ ((fiEnable && (2112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_6_io_in_control_0_shift_b <=( _mesh_21_6_io_out_control_0_shift) ^ ((fiEnable && (2113 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_6_io_in_control_0_dataflow_b <=( _mesh_21_6_io_out_control_0_dataflow) ^ ((fiEnable && (2114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_6_io_in_control_0_propagate_b <=( _mesh_21_6_io_out_control_0_propagate) ^ ((fiEnable && (2115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_6_io_out_valid_0) begin
			b_215_0 <=( _mesh_22_6_io_out_b_0) ^ ((fiEnable && (2116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1239_0 <=( _mesh_22_6_io_out_c_0) ^ ((fiEnable && (2117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_6_io_in_control_0_shift_b <=( _mesh_22_6_io_out_control_0_shift) ^ ((fiEnable && (2118 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_6_io_in_control_0_dataflow_b <=( _mesh_22_6_io_out_control_0_dataflow) ^ ((fiEnable && (2119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_6_io_in_control_0_propagate_b <=( _mesh_22_6_io_out_control_0_propagate) ^ ((fiEnable && (2120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_6_io_out_valid_0) begin
			b_216_0 <=( _mesh_23_6_io_out_b_0) ^ ((fiEnable && (2121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1240_0 <=( _mesh_23_6_io_out_c_0) ^ ((fiEnable && (2122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_6_io_in_control_0_shift_b <=( _mesh_23_6_io_out_control_0_shift) ^ ((fiEnable && (2123 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_6_io_in_control_0_dataflow_b <=( _mesh_23_6_io_out_control_0_dataflow) ^ ((fiEnable && (2124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_6_io_in_control_0_propagate_b <=( _mesh_23_6_io_out_control_0_propagate) ^ ((fiEnable && (2125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_6_io_out_valid_0) begin
			b_217_0 <=( _mesh_24_6_io_out_b_0) ^ ((fiEnable && (2126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1241_0 <=( _mesh_24_6_io_out_c_0) ^ ((fiEnable && (2127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_6_io_in_control_0_shift_b <=( _mesh_24_6_io_out_control_0_shift) ^ ((fiEnable && (2128 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_6_io_in_control_0_dataflow_b <=( _mesh_24_6_io_out_control_0_dataflow) ^ ((fiEnable && (2129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_6_io_in_control_0_propagate_b <=( _mesh_24_6_io_out_control_0_propagate) ^ ((fiEnable && (2130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_6_io_out_valid_0) begin
			b_218_0 <=( _mesh_25_6_io_out_b_0) ^ ((fiEnable && (2131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1242_0 <=( _mesh_25_6_io_out_c_0) ^ ((fiEnable && (2132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_6_io_in_control_0_shift_b <=( _mesh_25_6_io_out_control_0_shift) ^ ((fiEnable && (2133 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_6_io_in_control_0_dataflow_b <=( _mesh_25_6_io_out_control_0_dataflow) ^ ((fiEnable && (2134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_6_io_in_control_0_propagate_b <=( _mesh_25_6_io_out_control_0_propagate) ^ ((fiEnable && (2135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_6_io_out_valid_0) begin
			b_219_0 <=( _mesh_26_6_io_out_b_0) ^ ((fiEnable && (2136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1243_0 <=( _mesh_26_6_io_out_c_0) ^ ((fiEnable && (2137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_6_io_in_control_0_shift_b <=( _mesh_26_6_io_out_control_0_shift) ^ ((fiEnable && (2138 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_6_io_in_control_0_dataflow_b <=( _mesh_26_6_io_out_control_0_dataflow) ^ ((fiEnable && (2139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_6_io_in_control_0_propagate_b <=( _mesh_26_6_io_out_control_0_propagate) ^ ((fiEnable && (2140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_6_io_out_valid_0) begin
			b_220_0 <=( _mesh_27_6_io_out_b_0) ^ ((fiEnable && (2141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1244_0 <=( _mesh_27_6_io_out_c_0) ^ ((fiEnable && (2142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_6_io_in_control_0_shift_b <=( _mesh_27_6_io_out_control_0_shift) ^ ((fiEnable && (2143 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_6_io_in_control_0_dataflow_b <=( _mesh_27_6_io_out_control_0_dataflow) ^ ((fiEnable && (2144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_6_io_in_control_0_propagate_b <=( _mesh_27_6_io_out_control_0_propagate) ^ ((fiEnable && (2145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_6_io_out_valid_0) begin
			b_221_0 <=( _mesh_28_6_io_out_b_0) ^ ((fiEnable && (2146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1245_0 <=( _mesh_28_6_io_out_c_0) ^ ((fiEnable && (2147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_6_io_in_control_0_shift_b <=( _mesh_28_6_io_out_control_0_shift) ^ ((fiEnable && (2148 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_6_io_in_control_0_dataflow_b <=( _mesh_28_6_io_out_control_0_dataflow) ^ ((fiEnable && (2149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_6_io_in_control_0_propagate_b <=( _mesh_28_6_io_out_control_0_propagate) ^ ((fiEnable && (2150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_6_io_out_valid_0) begin
			b_222_0 <=( _mesh_29_6_io_out_b_0) ^ ((fiEnable && (2151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1246_0 <=( _mesh_29_6_io_out_c_0) ^ ((fiEnable && (2152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_6_io_in_control_0_shift_b <=( _mesh_29_6_io_out_control_0_shift) ^ ((fiEnable && (2153 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_6_io_in_control_0_dataflow_b <=( _mesh_29_6_io_out_control_0_dataflow) ^ ((fiEnable && (2154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_6_io_in_control_0_propagate_b <=( _mesh_29_6_io_out_control_0_propagate) ^ ((fiEnable && (2155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_6_io_out_valid_0) begin
			b_223_0 <=( _mesh_30_6_io_out_b_0) ^ ((fiEnable && (2156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1247_0 <=( _mesh_30_6_io_out_c_0) ^ ((fiEnable && (2157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_6_io_in_control_0_shift_b <=( _mesh_30_6_io_out_control_0_shift) ^ ((fiEnable && (2158 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_6_io_in_control_0_dataflow_b <=( _mesh_30_6_io_out_control_0_dataflow) ^ ((fiEnable && (2159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_6_io_in_control_0_propagate_b <=( _mesh_30_6_io_out_control_0_propagate) ^ ((fiEnable && (2160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_7_0) begin
			b_224_0 <=( io_in_b_7_0) ^ ((fiEnable && (2161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1248_0 <=( io_in_d_7_0) ^ ((fiEnable && (2162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_7_io_in_control_0_shift_b <=( io_in_control_7_0_shift) ^ ((fiEnable && (2163 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_7_io_in_control_0_dataflow_b <=( io_in_control_7_0_dataflow) ^ ((fiEnable && (2164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_7_io_in_control_0_propagate_b <=( io_in_control_7_0_propagate) ^ ((fiEnable && (2165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_7_io_out_valid_0) begin
			b_225_0 <=( _mesh_0_7_io_out_b_0) ^ ((fiEnable && (2166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1249_0 <=( _mesh_0_7_io_out_c_0) ^ ((fiEnable && (2167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_7_io_in_control_0_shift_b <=( _mesh_0_7_io_out_control_0_shift) ^ ((fiEnable && (2168 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_7_io_in_control_0_dataflow_b <=( _mesh_0_7_io_out_control_0_dataflow) ^ ((fiEnable && (2169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_7_io_in_control_0_propagate_b <=( _mesh_0_7_io_out_control_0_propagate) ^ ((fiEnable && (2170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_7_io_out_valid_0) begin
			b_226_0 <=( _mesh_1_7_io_out_b_0) ^ ((fiEnable && (2171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1250_0 <=( _mesh_1_7_io_out_c_0) ^ ((fiEnable && (2172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_7_io_in_control_0_shift_b <=( _mesh_1_7_io_out_control_0_shift) ^ ((fiEnable && (2173 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_7_io_in_control_0_dataflow_b <=( _mesh_1_7_io_out_control_0_dataflow) ^ ((fiEnable && (2174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_7_io_in_control_0_propagate_b <=( _mesh_1_7_io_out_control_0_propagate) ^ ((fiEnable && (2175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_7_io_out_valid_0) begin
			b_227_0 <=( _mesh_2_7_io_out_b_0) ^ ((fiEnable && (2176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1251_0 <=( _mesh_2_7_io_out_c_0) ^ ((fiEnable && (2177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_7_io_in_control_0_shift_b <=( _mesh_2_7_io_out_control_0_shift) ^ ((fiEnable && (2178 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_7_io_in_control_0_dataflow_b <=( _mesh_2_7_io_out_control_0_dataflow) ^ ((fiEnable && (2179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_7_io_in_control_0_propagate_b <=( _mesh_2_7_io_out_control_0_propagate) ^ ((fiEnable && (2180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_7_io_out_valid_0) begin
			b_228_0 <=( _mesh_3_7_io_out_b_0) ^ ((fiEnable && (2181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1252_0 <=( _mesh_3_7_io_out_c_0) ^ ((fiEnable && (2182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_7_io_in_control_0_shift_b <=( _mesh_3_7_io_out_control_0_shift) ^ ((fiEnable && (2183 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_7_io_in_control_0_dataflow_b <=( _mesh_3_7_io_out_control_0_dataflow) ^ ((fiEnable && (2184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_7_io_in_control_0_propagate_b <=( _mesh_3_7_io_out_control_0_propagate) ^ ((fiEnable && (2185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_7_io_out_valid_0) begin
			b_229_0 <=( _mesh_4_7_io_out_b_0) ^ ((fiEnable && (2186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1253_0 <=( _mesh_4_7_io_out_c_0) ^ ((fiEnable && (2187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_7_io_in_control_0_shift_b <=( _mesh_4_7_io_out_control_0_shift) ^ ((fiEnable && (2188 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_7_io_in_control_0_dataflow_b <=( _mesh_4_7_io_out_control_0_dataflow) ^ ((fiEnable && (2189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_7_io_in_control_0_propagate_b <=( _mesh_4_7_io_out_control_0_propagate) ^ ((fiEnable && (2190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_7_io_out_valid_0) begin
			b_230_0 <=( _mesh_5_7_io_out_b_0) ^ ((fiEnable && (2191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1254_0 <=( _mesh_5_7_io_out_c_0) ^ ((fiEnable && (2192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_7_io_in_control_0_shift_b <=( _mesh_5_7_io_out_control_0_shift) ^ ((fiEnable && (2193 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_7_io_in_control_0_dataflow_b <=( _mesh_5_7_io_out_control_0_dataflow) ^ ((fiEnable && (2194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_7_io_in_control_0_propagate_b <=( _mesh_5_7_io_out_control_0_propagate) ^ ((fiEnable && (2195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_7_io_out_valid_0) begin
			b_231_0 <=( _mesh_6_7_io_out_b_0) ^ ((fiEnable && (2196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1255_0 <=( _mesh_6_7_io_out_c_0) ^ ((fiEnable && (2197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_7_io_in_control_0_shift_b <=( _mesh_6_7_io_out_control_0_shift) ^ ((fiEnable && (2198 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_7_io_in_control_0_dataflow_b <=( _mesh_6_7_io_out_control_0_dataflow) ^ ((fiEnable && (2199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_7_io_in_control_0_propagate_b <=( _mesh_6_7_io_out_control_0_propagate) ^ ((fiEnable && (2200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_7_io_out_valid_0) begin
			b_232_0 <=( _mesh_7_7_io_out_b_0) ^ ((fiEnable && (2201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1256_0 <=( _mesh_7_7_io_out_c_0) ^ ((fiEnable && (2202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_7_io_in_control_0_shift_b <=( _mesh_7_7_io_out_control_0_shift) ^ ((fiEnable && (2203 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_7_io_in_control_0_dataflow_b <=( _mesh_7_7_io_out_control_0_dataflow) ^ ((fiEnable && (2204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_7_io_in_control_0_propagate_b <=( _mesh_7_7_io_out_control_0_propagate) ^ ((fiEnable && (2205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_7_io_out_valid_0) begin
			b_233_0 <=( _mesh_8_7_io_out_b_0) ^ ((fiEnable && (2206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1257_0 <=( _mesh_8_7_io_out_c_0) ^ ((fiEnable && (2207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_7_io_in_control_0_shift_b <=( _mesh_8_7_io_out_control_0_shift) ^ ((fiEnable && (2208 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_7_io_in_control_0_dataflow_b <=( _mesh_8_7_io_out_control_0_dataflow) ^ ((fiEnable && (2209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_7_io_in_control_0_propagate_b <=( _mesh_8_7_io_out_control_0_propagate) ^ ((fiEnable && (2210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_7_io_out_valid_0) begin
			b_234_0 <=( _mesh_9_7_io_out_b_0) ^ ((fiEnable && (2211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1258_0 <=( _mesh_9_7_io_out_c_0) ^ ((fiEnable && (2212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_7_io_in_control_0_shift_b <=( _mesh_9_7_io_out_control_0_shift) ^ ((fiEnable && (2213 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_7_io_in_control_0_dataflow_b <=( _mesh_9_7_io_out_control_0_dataflow) ^ ((fiEnable && (2214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_7_io_in_control_0_propagate_b <=( _mesh_9_7_io_out_control_0_propagate) ^ ((fiEnable && (2215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_7_io_out_valid_0) begin
			b_235_0 <=( _mesh_10_7_io_out_b_0) ^ ((fiEnable && (2216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1259_0 <=( _mesh_10_7_io_out_c_0) ^ ((fiEnable && (2217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_7_io_in_control_0_shift_b <=( _mesh_10_7_io_out_control_0_shift) ^ ((fiEnable && (2218 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_7_io_in_control_0_dataflow_b <=( _mesh_10_7_io_out_control_0_dataflow) ^ ((fiEnable && (2219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_7_io_in_control_0_propagate_b <=( _mesh_10_7_io_out_control_0_propagate) ^ ((fiEnable && (2220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_7_io_out_valid_0) begin
			b_236_0 <=( _mesh_11_7_io_out_b_0) ^ ((fiEnable && (2221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1260_0 <=( _mesh_11_7_io_out_c_0) ^ ((fiEnable && (2222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_7_io_in_control_0_shift_b <=( _mesh_11_7_io_out_control_0_shift) ^ ((fiEnable && (2223 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_7_io_in_control_0_dataflow_b <=( _mesh_11_7_io_out_control_0_dataflow) ^ ((fiEnable && (2224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_7_io_in_control_0_propagate_b <=( _mesh_11_7_io_out_control_0_propagate) ^ ((fiEnable && (2225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_7_io_out_valid_0) begin
			b_237_0 <=( _mesh_12_7_io_out_b_0) ^ ((fiEnable && (2226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1261_0 <=( _mesh_12_7_io_out_c_0) ^ ((fiEnable && (2227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_7_io_in_control_0_shift_b <=( _mesh_12_7_io_out_control_0_shift) ^ ((fiEnable && (2228 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_7_io_in_control_0_dataflow_b <=( _mesh_12_7_io_out_control_0_dataflow) ^ ((fiEnable && (2229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_7_io_in_control_0_propagate_b <=( _mesh_12_7_io_out_control_0_propagate) ^ ((fiEnable && (2230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_7_io_out_valid_0) begin
			b_238_0 <=( _mesh_13_7_io_out_b_0) ^ ((fiEnable && (2231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1262_0 <=( _mesh_13_7_io_out_c_0) ^ ((fiEnable && (2232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_7_io_in_control_0_shift_b <=( _mesh_13_7_io_out_control_0_shift) ^ ((fiEnable && (2233 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_7_io_in_control_0_dataflow_b <=( _mesh_13_7_io_out_control_0_dataflow) ^ ((fiEnable && (2234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_7_io_in_control_0_propagate_b <=( _mesh_13_7_io_out_control_0_propagate) ^ ((fiEnable && (2235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_7_io_out_valid_0) begin
			b_239_0 <=( _mesh_14_7_io_out_b_0) ^ ((fiEnable && (2236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1263_0 <=( _mesh_14_7_io_out_c_0) ^ ((fiEnable && (2237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_7_io_in_control_0_shift_b <=( _mesh_14_7_io_out_control_0_shift) ^ ((fiEnable && (2238 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_7_io_in_control_0_dataflow_b <=( _mesh_14_7_io_out_control_0_dataflow) ^ ((fiEnable && (2239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_7_io_in_control_0_propagate_b <=( _mesh_14_7_io_out_control_0_propagate) ^ ((fiEnable && (2240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_7_io_out_valid_0) begin
			b_240_0 <=( _mesh_15_7_io_out_b_0) ^ ((fiEnable && (2241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1264_0 <=( _mesh_15_7_io_out_c_0) ^ ((fiEnable && (2242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_7_io_in_control_0_shift_b <=( _mesh_15_7_io_out_control_0_shift) ^ ((fiEnable && (2243 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_7_io_in_control_0_dataflow_b <=( _mesh_15_7_io_out_control_0_dataflow) ^ ((fiEnable && (2244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_7_io_in_control_0_propagate_b <=( _mesh_15_7_io_out_control_0_propagate) ^ ((fiEnable && (2245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_7_io_out_valid_0) begin
			b_241_0 <=( _mesh_16_7_io_out_b_0) ^ ((fiEnable && (2246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1265_0 <=( _mesh_16_7_io_out_c_0) ^ ((fiEnable && (2247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_7_io_in_control_0_shift_b <=( _mesh_16_7_io_out_control_0_shift) ^ ((fiEnable && (2248 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_7_io_in_control_0_dataflow_b <=( _mesh_16_7_io_out_control_0_dataflow) ^ ((fiEnable && (2249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_7_io_in_control_0_propagate_b <=( _mesh_16_7_io_out_control_0_propagate) ^ ((fiEnable && (2250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_7_io_out_valid_0) begin
			b_242_0 <=( _mesh_17_7_io_out_b_0) ^ ((fiEnable && (2251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1266_0 <=( _mesh_17_7_io_out_c_0) ^ ((fiEnable && (2252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_7_io_in_control_0_shift_b <=( _mesh_17_7_io_out_control_0_shift) ^ ((fiEnable && (2253 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_7_io_in_control_0_dataflow_b <=( _mesh_17_7_io_out_control_0_dataflow) ^ ((fiEnable && (2254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_7_io_in_control_0_propagate_b <=( _mesh_17_7_io_out_control_0_propagate) ^ ((fiEnable && (2255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_7_io_out_valid_0) begin
			b_243_0 <=( _mesh_18_7_io_out_b_0) ^ ((fiEnable && (2256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1267_0 <=( _mesh_18_7_io_out_c_0) ^ ((fiEnable && (2257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_7_io_in_control_0_shift_b <=( _mesh_18_7_io_out_control_0_shift) ^ ((fiEnable && (2258 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_7_io_in_control_0_dataflow_b <=( _mesh_18_7_io_out_control_0_dataflow) ^ ((fiEnable && (2259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_7_io_in_control_0_propagate_b <=( _mesh_18_7_io_out_control_0_propagate) ^ ((fiEnable && (2260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_7_io_out_valid_0) begin
			b_244_0 <=( _mesh_19_7_io_out_b_0) ^ ((fiEnable && (2261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1268_0 <=( _mesh_19_7_io_out_c_0) ^ ((fiEnable && (2262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_7_io_in_control_0_shift_b <=( _mesh_19_7_io_out_control_0_shift) ^ ((fiEnable && (2263 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_7_io_in_control_0_dataflow_b <=( _mesh_19_7_io_out_control_0_dataflow) ^ ((fiEnable && (2264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_7_io_in_control_0_propagate_b <=( _mesh_19_7_io_out_control_0_propagate) ^ ((fiEnable && (2265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_7_io_out_valid_0) begin
			b_245_0 <=( _mesh_20_7_io_out_b_0) ^ ((fiEnable && (2266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1269_0 <=( _mesh_20_7_io_out_c_0) ^ ((fiEnable && (2267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_7_io_in_control_0_shift_b <=( _mesh_20_7_io_out_control_0_shift) ^ ((fiEnable && (2268 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_7_io_in_control_0_dataflow_b <=( _mesh_20_7_io_out_control_0_dataflow) ^ ((fiEnable && (2269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_7_io_in_control_0_propagate_b <=( _mesh_20_7_io_out_control_0_propagate) ^ ((fiEnable && (2270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_7_io_out_valid_0) begin
			b_246_0 <=( _mesh_21_7_io_out_b_0) ^ ((fiEnable && (2271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1270_0 <=( _mesh_21_7_io_out_c_0) ^ ((fiEnable && (2272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_7_io_in_control_0_shift_b <=( _mesh_21_7_io_out_control_0_shift) ^ ((fiEnable && (2273 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_7_io_in_control_0_dataflow_b <=( _mesh_21_7_io_out_control_0_dataflow) ^ ((fiEnable && (2274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_7_io_in_control_0_propagate_b <=( _mesh_21_7_io_out_control_0_propagate) ^ ((fiEnable && (2275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_7_io_out_valid_0) begin
			b_247_0 <=( _mesh_22_7_io_out_b_0) ^ ((fiEnable && (2276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1271_0 <=( _mesh_22_7_io_out_c_0) ^ ((fiEnable && (2277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_7_io_in_control_0_shift_b <=( _mesh_22_7_io_out_control_0_shift) ^ ((fiEnable && (2278 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_7_io_in_control_0_dataflow_b <=( _mesh_22_7_io_out_control_0_dataflow) ^ ((fiEnable && (2279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_7_io_in_control_0_propagate_b <=( _mesh_22_7_io_out_control_0_propagate) ^ ((fiEnable && (2280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_7_io_out_valid_0) begin
			b_248_0 <=( _mesh_23_7_io_out_b_0) ^ ((fiEnable && (2281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1272_0 <=( _mesh_23_7_io_out_c_0) ^ ((fiEnable && (2282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_7_io_in_control_0_shift_b <=( _mesh_23_7_io_out_control_0_shift) ^ ((fiEnable && (2283 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_7_io_in_control_0_dataflow_b <=( _mesh_23_7_io_out_control_0_dataflow) ^ ((fiEnable && (2284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_7_io_in_control_0_propagate_b <=( _mesh_23_7_io_out_control_0_propagate) ^ ((fiEnable && (2285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_7_io_out_valid_0) begin
			b_249_0 <=( _mesh_24_7_io_out_b_0) ^ ((fiEnable && (2286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1273_0 <=( _mesh_24_7_io_out_c_0) ^ ((fiEnable && (2287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_7_io_in_control_0_shift_b <=( _mesh_24_7_io_out_control_0_shift) ^ ((fiEnable && (2288 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_7_io_in_control_0_dataflow_b <=( _mesh_24_7_io_out_control_0_dataflow) ^ ((fiEnable && (2289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_7_io_in_control_0_propagate_b <=( _mesh_24_7_io_out_control_0_propagate) ^ ((fiEnable && (2290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_7_io_out_valid_0) begin
			b_250_0 <=( _mesh_25_7_io_out_b_0) ^ ((fiEnable && (2291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1274_0 <=( _mesh_25_7_io_out_c_0) ^ ((fiEnable && (2292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_7_io_in_control_0_shift_b <=( _mesh_25_7_io_out_control_0_shift) ^ ((fiEnable && (2293 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_7_io_in_control_0_dataflow_b <=( _mesh_25_7_io_out_control_0_dataflow) ^ ((fiEnable && (2294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_7_io_in_control_0_propagate_b <=( _mesh_25_7_io_out_control_0_propagate) ^ ((fiEnable && (2295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_7_io_out_valid_0) begin
			b_251_0 <=( _mesh_26_7_io_out_b_0) ^ ((fiEnable && (2296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1275_0 <=( _mesh_26_7_io_out_c_0) ^ ((fiEnable && (2297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_7_io_in_control_0_shift_b <=( _mesh_26_7_io_out_control_0_shift) ^ ((fiEnable && (2298 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_7_io_in_control_0_dataflow_b <=( _mesh_26_7_io_out_control_0_dataflow) ^ ((fiEnable && (2299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_7_io_in_control_0_propagate_b <=( _mesh_26_7_io_out_control_0_propagate) ^ ((fiEnable && (2300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_7_io_out_valid_0) begin
			b_252_0 <=( _mesh_27_7_io_out_b_0) ^ ((fiEnable && (2301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1276_0 <=( _mesh_27_7_io_out_c_0) ^ ((fiEnable && (2302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_7_io_in_control_0_shift_b <=( _mesh_27_7_io_out_control_0_shift) ^ ((fiEnable && (2303 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_7_io_in_control_0_dataflow_b <=( _mesh_27_7_io_out_control_0_dataflow) ^ ((fiEnable && (2304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_7_io_in_control_0_propagate_b <=( _mesh_27_7_io_out_control_0_propagate) ^ ((fiEnable && (2305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_7_io_out_valid_0) begin
			b_253_0 <=( _mesh_28_7_io_out_b_0) ^ ((fiEnable && (2306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1277_0 <=( _mesh_28_7_io_out_c_0) ^ ((fiEnable && (2307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_7_io_in_control_0_shift_b <=( _mesh_28_7_io_out_control_0_shift) ^ ((fiEnable && (2308 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_7_io_in_control_0_dataflow_b <=( _mesh_28_7_io_out_control_0_dataflow) ^ ((fiEnable && (2309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_7_io_in_control_0_propagate_b <=( _mesh_28_7_io_out_control_0_propagate) ^ ((fiEnable && (2310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_7_io_out_valid_0) begin
			b_254_0 <=( _mesh_29_7_io_out_b_0) ^ ((fiEnable && (2311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1278_0 <=( _mesh_29_7_io_out_c_0) ^ ((fiEnable && (2312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_7_io_in_control_0_shift_b <=( _mesh_29_7_io_out_control_0_shift) ^ ((fiEnable && (2313 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_7_io_in_control_0_dataflow_b <=( _mesh_29_7_io_out_control_0_dataflow) ^ ((fiEnable && (2314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_7_io_in_control_0_propagate_b <=( _mesh_29_7_io_out_control_0_propagate) ^ ((fiEnable && (2315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_7_io_out_valid_0) begin
			b_255_0 <=( _mesh_30_7_io_out_b_0) ^ ((fiEnable && (2316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1279_0 <=( _mesh_30_7_io_out_c_0) ^ ((fiEnable && (2317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_7_io_in_control_0_shift_b <=( _mesh_30_7_io_out_control_0_shift) ^ ((fiEnable && (2318 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_7_io_in_control_0_dataflow_b <=( _mesh_30_7_io_out_control_0_dataflow) ^ ((fiEnable && (2319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_7_io_in_control_0_propagate_b <=( _mesh_30_7_io_out_control_0_propagate) ^ ((fiEnable && (2320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_8_0) begin
			b_256_0 <=( io_in_b_8_0) ^ ((fiEnable && (2321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1280_0 <=( io_in_d_8_0) ^ ((fiEnable && (2322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_8_io_in_control_0_shift_b <=( io_in_control_8_0_shift) ^ ((fiEnable && (2323 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_8_io_in_control_0_dataflow_b <=( io_in_control_8_0_dataflow) ^ ((fiEnable && (2324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_8_io_in_control_0_propagate_b <=( io_in_control_8_0_propagate) ^ ((fiEnable && (2325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_8_io_out_valid_0) begin
			b_257_0 <=( _mesh_0_8_io_out_b_0) ^ ((fiEnable && (2326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1281_0 <=( _mesh_0_8_io_out_c_0) ^ ((fiEnable && (2327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_8_io_in_control_0_shift_b <=( _mesh_0_8_io_out_control_0_shift) ^ ((fiEnable && (2328 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_8_io_in_control_0_dataflow_b <=( _mesh_0_8_io_out_control_0_dataflow) ^ ((fiEnable && (2329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_8_io_in_control_0_propagate_b <=( _mesh_0_8_io_out_control_0_propagate) ^ ((fiEnable && (2330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_8_io_out_valid_0) begin
			b_258_0 <=( _mesh_1_8_io_out_b_0) ^ ((fiEnable && (2331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1282_0 <=( _mesh_1_8_io_out_c_0) ^ ((fiEnable && (2332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_8_io_in_control_0_shift_b <=( _mesh_1_8_io_out_control_0_shift) ^ ((fiEnable && (2333 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_8_io_in_control_0_dataflow_b <=( _mesh_1_8_io_out_control_0_dataflow) ^ ((fiEnable && (2334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_8_io_in_control_0_propagate_b <=( _mesh_1_8_io_out_control_0_propagate) ^ ((fiEnable && (2335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_8_io_out_valid_0) begin
			b_259_0 <=( _mesh_2_8_io_out_b_0) ^ ((fiEnable && (2336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1283_0 <=( _mesh_2_8_io_out_c_0) ^ ((fiEnable && (2337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_8_io_in_control_0_shift_b <=( _mesh_2_8_io_out_control_0_shift) ^ ((fiEnable && (2338 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_8_io_in_control_0_dataflow_b <=( _mesh_2_8_io_out_control_0_dataflow) ^ ((fiEnable && (2339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_8_io_in_control_0_propagate_b <=( _mesh_2_8_io_out_control_0_propagate) ^ ((fiEnable && (2340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_8_io_out_valid_0) begin
			b_260_0 <=( _mesh_3_8_io_out_b_0) ^ ((fiEnable && (2341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1284_0 <=( _mesh_3_8_io_out_c_0) ^ ((fiEnable && (2342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_8_io_in_control_0_shift_b <=( _mesh_3_8_io_out_control_0_shift) ^ ((fiEnable && (2343 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_8_io_in_control_0_dataflow_b <=( _mesh_3_8_io_out_control_0_dataflow) ^ ((fiEnable && (2344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_8_io_in_control_0_propagate_b <=( _mesh_3_8_io_out_control_0_propagate) ^ ((fiEnable && (2345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_8_io_out_valid_0) begin
			b_261_0 <=( _mesh_4_8_io_out_b_0) ^ ((fiEnable && (2346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1285_0 <=( _mesh_4_8_io_out_c_0) ^ ((fiEnable && (2347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_8_io_in_control_0_shift_b <=( _mesh_4_8_io_out_control_0_shift) ^ ((fiEnable && (2348 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_8_io_in_control_0_dataflow_b <=( _mesh_4_8_io_out_control_0_dataflow) ^ ((fiEnable && (2349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_8_io_in_control_0_propagate_b <=( _mesh_4_8_io_out_control_0_propagate) ^ ((fiEnable && (2350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_8_io_out_valid_0) begin
			b_262_0 <=( _mesh_5_8_io_out_b_0) ^ ((fiEnable && (2351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1286_0 <=( _mesh_5_8_io_out_c_0) ^ ((fiEnable && (2352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_8_io_in_control_0_shift_b <=( _mesh_5_8_io_out_control_0_shift) ^ ((fiEnable && (2353 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_8_io_in_control_0_dataflow_b <=( _mesh_5_8_io_out_control_0_dataflow) ^ ((fiEnable && (2354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_8_io_in_control_0_propagate_b <=( _mesh_5_8_io_out_control_0_propagate) ^ ((fiEnable && (2355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_8_io_out_valid_0) begin
			b_263_0 <=( _mesh_6_8_io_out_b_0) ^ ((fiEnable && (2356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1287_0 <=( _mesh_6_8_io_out_c_0) ^ ((fiEnable && (2357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_8_io_in_control_0_shift_b <=( _mesh_6_8_io_out_control_0_shift) ^ ((fiEnable && (2358 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_8_io_in_control_0_dataflow_b <=( _mesh_6_8_io_out_control_0_dataflow) ^ ((fiEnable && (2359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_8_io_in_control_0_propagate_b <=( _mesh_6_8_io_out_control_0_propagate) ^ ((fiEnable && (2360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_8_io_out_valid_0) begin
			b_264_0 <=( _mesh_7_8_io_out_b_0) ^ ((fiEnable && (2361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1288_0 <=( _mesh_7_8_io_out_c_0) ^ ((fiEnable && (2362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_8_io_in_control_0_shift_b <=( _mesh_7_8_io_out_control_0_shift) ^ ((fiEnable && (2363 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_8_io_in_control_0_dataflow_b <=( _mesh_7_8_io_out_control_0_dataflow) ^ ((fiEnable && (2364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_8_io_in_control_0_propagate_b <=( _mesh_7_8_io_out_control_0_propagate) ^ ((fiEnable && (2365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_8_io_out_valid_0) begin
			b_265_0 <=( _mesh_8_8_io_out_b_0) ^ ((fiEnable && (2366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1289_0 <=( _mesh_8_8_io_out_c_0) ^ ((fiEnable && (2367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_8_io_in_control_0_shift_b <=( _mesh_8_8_io_out_control_0_shift) ^ ((fiEnable && (2368 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_8_io_in_control_0_dataflow_b <=( _mesh_8_8_io_out_control_0_dataflow) ^ ((fiEnable && (2369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_8_io_in_control_0_propagate_b <=( _mesh_8_8_io_out_control_0_propagate) ^ ((fiEnable && (2370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_8_io_out_valid_0) begin
			b_266_0 <=( _mesh_9_8_io_out_b_0) ^ ((fiEnable && (2371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1290_0 <=( _mesh_9_8_io_out_c_0) ^ ((fiEnable && (2372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_8_io_in_control_0_shift_b <=( _mesh_9_8_io_out_control_0_shift) ^ ((fiEnable && (2373 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_8_io_in_control_0_dataflow_b <=( _mesh_9_8_io_out_control_0_dataflow) ^ ((fiEnable && (2374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_8_io_in_control_0_propagate_b <=( _mesh_9_8_io_out_control_0_propagate) ^ ((fiEnable && (2375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_8_io_out_valid_0) begin
			b_267_0 <=( _mesh_10_8_io_out_b_0) ^ ((fiEnable && (2376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1291_0 <=( _mesh_10_8_io_out_c_0) ^ ((fiEnable && (2377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_8_io_in_control_0_shift_b <=( _mesh_10_8_io_out_control_0_shift) ^ ((fiEnable && (2378 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_8_io_in_control_0_dataflow_b <=( _mesh_10_8_io_out_control_0_dataflow) ^ ((fiEnable && (2379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_8_io_in_control_0_propagate_b <=( _mesh_10_8_io_out_control_0_propagate) ^ ((fiEnable && (2380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_8_io_out_valid_0) begin
			b_268_0 <=( _mesh_11_8_io_out_b_0) ^ ((fiEnable && (2381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1292_0 <=( _mesh_11_8_io_out_c_0) ^ ((fiEnable && (2382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_8_io_in_control_0_shift_b <=( _mesh_11_8_io_out_control_0_shift) ^ ((fiEnable && (2383 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_8_io_in_control_0_dataflow_b <=( _mesh_11_8_io_out_control_0_dataflow) ^ ((fiEnable && (2384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_8_io_in_control_0_propagate_b <=( _mesh_11_8_io_out_control_0_propagate) ^ ((fiEnable && (2385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_8_io_out_valid_0) begin
			b_269_0 <=( _mesh_12_8_io_out_b_0) ^ ((fiEnable && (2386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1293_0 <=( _mesh_12_8_io_out_c_0) ^ ((fiEnable && (2387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_8_io_in_control_0_shift_b <=( _mesh_12_8_io_out_control_0_shift) ^ ((fiEnable && (2388 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_8_io_in_control_0_dataflow_b <=( _mesh_12_8_io_out_control_0_dataflow) ^ ((fiEnable && (2389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_8_io_in_control_0_propagate_b <=( _mesh_12_8_io_out_control_0_propagate) ^ ((fiEnable && (2390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_8_io_out_valid_0) begin
			b_270_0 <=( _mesh_13_8_io_out_b_0) ^ ((fiEnable && (2391 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1294_0 <=( _mesh_13_8_io_out_c_0) ^ ((fiEnable && (2392 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_8_io_in_control_0_shift_b <=( _mesh_13_8_io_out_control_0_shift) ^ ((fiEnable && (2393 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_8_io_in_control_0_dataflow_b <=( _mesh_13_8_io_out_control_0_dataflow) ^ ((fiEnable && (2394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_8_io_in_control_0_propagate_b <=( _mesh_13_8_io_out_control_0_propagate) ^ ((fiEnable && (2395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_8_io_out_valid_0) begin
			b_271_0 <=( _mesh_14_8_io_out_b_0) ^ ((fiEnable && (2396 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1295_0 <=( _mesh_14_8_io_out_c_0) ^ ((fiEnable && (2397 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_8_io_in_control_0_shift_b <=( _mesh_14_8_io_out_control_0_shift) ^ ((fiEnable && (2398 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_8_io_in_control_0_dataflow_b <=( _mesh_14_8_io_out_control_0_dataflow) ^ ((fiEnable && (2399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_8_io_in_control_0_propagate_b <=( _mesh_14_8_io_out_control_0_propagate) ^ ((fiEnable && (2400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_8_io_out_valid_0) begin
			b_272_0 <=( _mesh_15_8_io_out_b_0) ^ ((fiEnable && (2401 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1296_0 <=( _mesh_15_8_io_out_c_0) ^ ((fiEnable && (2402 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_8_io_in_control_0_shift_b <=( _mesh_15_8_io_out_control_0_shift) ^ ((fiEnable && (2403 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_8_io_in_control_0_dataflow_b <=( _mesh_15_8_io_out_control_0_dataflow) ^ ((fiEnable && (2404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_8_io_in_control_0_propagate_b <=( _mesh_15_8_io_out_control_0_propagate) ^ ((fiEnable && (2405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_8_io_out_valid_0) begin
			b_273_0 <=( _mesh_16_8_io_out_b_0) ^ ((fiEnable && (2406 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1297_0 <=( _mesh_16_8_io_out_c_0) ^ ((fiEnable && (2407 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_8_io_in_control_0_shift_b <=( _mesh_16_8_io_out_control_0_shift) ^ ((fiEnable && (2408 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_8_io_in_control_0_dataflow_b <=( _mesh_16_8_io_out_control_0_dataflow) ^ ((fiEnable && (2409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_8_io_in_control_0_propagate_b <=( _mesh_16_8_io_out_control_0_propagate) ^ ((fiEnable && (2410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_8_io_out_valid_0) begin
			b_274_0 <=( _mesh_17_8_io_out_b_0) ^ ((fiEnable && (2411 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1298_0 <=( _mesh_17_8_io_out_c_0) ^ ((fiEnable && (2412 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_8_io_in_control_0_shift_b <=( _mesh_17_8_io_out_control_0_shift) ^ ((fiEnable && (2413 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_8_io_in_control_0_dataflow_b <=( _mesh_17_8_io_out_control_0_dataflow) ^ ((fiEnable && (2414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_8_io_in_control_0_propagate_b <=( _mesh_17_8_io_out_control_0_propagate) ^ ((fiEnable && (2415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_8_io_out_valid_0) begin
			b_275_0 <=( _mesh_18_8_io_out_b_0) ^ ((fiEnable && (2416 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1299_0 <=( _mesh_18_8_io_out_c_0) ^ ((fiEnable && (2417 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_8_io_in_control_0_shift_b <=( _mesh_18_8_io_out_control_0_shift) ^ ((fiEnable && (2418 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_8_io_in_control_0_dataflow_b <=( _mesh_18_8_io_out_control_0_dataflow) ^ ((fiEnable && (2419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_8_io_in_control_0_propagate_b <=( _mesh_18_8_io_out_control_0_propagate) ^ ((fiEnable && (2420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_8_io_out_valid_0) begin
			b_276_0 <=( _mesh_19_8_io_out_b_0) ^ ((fiEnable && (2421 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1300_0 <=( _mesh_19_8_io_out_c_0) ^ ((fiEnable && (2422 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_8_io_in_control_0_shift_b <=( _mesh_19_8_io_out_control_0_shift) ^ ((fiEnable && (2423 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_8_io_in_control_0_dataflow_b <=( _mesh_19_8_io_out_control_0_dataflow) ^ ((fiEnable && (2424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_8_io_in_control_0_propagate_b <=( _mesh_19_8_io_out_control_0_propagate) ^ ((fiEnable && (2425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_8_io_out_valid_0) begin
			b_277_0 <=( _mesh_20_8_io_out_b_0) ^ ((fiEnable && (2426 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1301_0 <=( _mesh_20_8_io_out_c_0) ^ ((fiEnable && (2427 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_8_io_in_control_0_shift_b <=( _mesh_20_8_io_out_control_0_shift) ^ ((fiEnable && (2428 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_8_io_in_control_0_dataflow_b <=( _mesh_20_8_io_out_control_0_dataflow) ^ ((fiEnable && (2429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_8_io_in_control_0_propagate_b <=( _mesh_20_8_io_out_control_0_propagate) ^ ((fiEnable && (2430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_8_io_out_valid_0) begin
			b_278_0 <=( _mesh_21_8_io_out_b_0) ^ ((fiEnable && (2431 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1302_0 <=( _mesh_21_8_io_out_c_0) ^ ((fiEnable && (2432 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_8_io_in_control_0_shift_b <=( _mesh_21_8_io_out_control_0_shift) ^ ((fiEnable && (2433 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_8_io_in_control_0_dataflow_b <=( _mesh_21_8_io_out_control_0_dataflow) ^ ((fiEnable && (2434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_8_io_in_control_0_propagate_b <=( _mesh_21_8_io_out_control_0_propagate) ^ ((fiEnable && (2435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_8_io_out_valid_0) begin
			b_279_0 <=( _mesh_22_8_io_out_b_0) ^ ((fiEnable && (2436 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1303_0 <=( _mesh_22_8_io_out_c_0) ^ ((fiEnable && (2437 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_8_io_in_control_0_shift_b <=( _mesh_22_8_io_out_control_0_shift) ^ ((fiEnable && (2438 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_8_io_in_control_0_dataflow_b <=( _mesh_22_8_io_out_control_0_dataflow) ^ ((fiEnable && (2439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_8_io_in_control_0_propagate_b <=( _mesh_22_8_io_out_control_0_propagate) ^ ((fiEnable && (2440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_8_io_out_valid_0) begin
			b_280_0 <=( _mesh_23_8_io_out_b_0) ^ ((fiEnable && (2441 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1304_0 <=( _mesh_23_8_io_out_c_0) ^ ((fiEnable && (2442 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_8_io_in_control_0_shift_b <=( _mesh_23_8_io_out_control_0_shift) ^ ((fiEnable && (2443 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_8_io_in_control_0_dataflow_b <=( _mesh_23_8_io_out_control_0_dataflow) ^ ((fiEnable && (2444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_8_io_in_control_0_propagate_b <=( _mesh_23_8_io_out_control_0_propagate) ^ ((fiEnable && (2445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_8_io_out_valid_0) begin
			b_281_0 <=( _mesh_24_8_io_out_b_0) ^ ((fiEnable && (2446 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1305_0 <=( _mesh_24_8_io_out_c_0) ^ ((fiEnable && (2447 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_8_io_in_control_0_shift_b <=( _mesh_24_8_io_out_control_0_shift) ^ ((fiEnable && (2448 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_8_io_in_control_0_dataflow_b <=( _mesh_24_8_io_out_control_0_dataflow) ^ ((fiEnable && (2449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_8_io_in_control_0_propagate_b <=( _mesh_24_8_io_out_control_0_propagate) ^ ((fiEnable && (2450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_8_io_out_valid_0) begin
			b_282_0 <=( _mesh_25_8_io_out_b_0) ^ ((fiEnable && (2451 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1306_0 <=( _mesh_25_8_io_out_c_0) ^ ((fiEnable && (2452 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_8_io_in_control_0_shift_b <=( _mesh_25_8_io_out_control_0_shift) ^ ((fiEnable && (2453 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_8_io_in_control_0_dataflow_b <=( _mesh_25_8_io_out_control_0_dataflow) ^ ((fiEnable && (2454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_8_io_in_control_0_propagate_b <=( _mesh_25_8_io_out_control_0_propagate) ^ ((fiEnable && (2455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_8_io_out_valid_0) begin
			b_283_0 <=( _mesh_26_8_io_out_b_0) ^ ((fiEnable && (2456 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1307_0 <=( _mesh_26_8_io_out_c_0) ^ ((fiEnable && (2457 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_8_io_in_control_0_shift_b <=( _mesh_26_8_io_out_control_0_shift) ^ ((fiEnable && (2458 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_8_io_in_control_0_dataflow_b <=( _mesh_26_8_io_out_control_0_dataflow) ^ ((fiEnable && (2459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_8_io_in_control_0_propagate_b <=( _mesh_26_8_io_out_control_0_propagate) ^ ((fiEnable && (2460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_8_io_out_valid_0) begin
			b_284_0 <=( _mesh_27_8_io_out_b_0) ^ ((fiEnable && (2461 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1308_0 <=( _mesh_27_8_io_out_c_0) ^ ((fiEnable && (2462 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_8_io_in_control_0_shift_b <=( _mesh_27_8_io_out_control_0_shift) ^ ((fiEnable && (2463 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_8_io_in_control_0_dataflow_b <=( _mesh_27_8_io_out_control_0_dataflow) ^ ((fiEnable && (2464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_8_io_in_control_0_propagate_b <=( _mesh_27_8_io_out_control_0_propagate) ^ ((fiEnable && (2465 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_8_io_out_valid_0) begin
			b_285_0 <=( _mesh_28_8_io_out_b_0) ^ ((fiEnable && (2466 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1309_0 <=( _mesh_28_8_io_out_c_0) ^ ((fiEnable && (2467 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_8_io_in_control_0_shift_b <=( _mesh_28_8_io_out_control_0_shift) ^ ((fiEnable && (2468 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_8_io_in_control_0_dataflow_b <=( _mesh_28_8_io_out_control_0_dataflow) ^ ((fiEnable && (2469 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_8_io_in_control_0_propagate_b <=( _mesh_28_8_io_out_control_0_propagate) ^ ((fiEnable && (2470 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_8_io_out_valid_0) begin
			b_286_0 <=( _mesh_29_8_io_out_b_0) ^ ((fiEnable && (2471 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1310_0 <=( _mesh_29_8_io_out_c_0) ^ ((fiEnable && (2472 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_8_io_in_control_0_shift_b <=( _mesh_29_8_io_out_control_0_shift) ^ ((fiEnable && (2473 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_8_io_in_control_0_dataflow_b <=( _mesh_29_8_io_out_control_0_dataflow) ^ ((fiEnable && (2474 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_8_io_in_control_0_propagate_b <=( _mesh_29_8_io_out_control_0_propagate) ^ ((fiEnable && (2475 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_8_io_out_valid_0) begin
			b_287_0 <=( _mesh_30_8_io_out_b_0) ^ ((fiEnable && (2476 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1311_0 <=( _mesh_30_8_io_out_c_0) ^ ((fiEnable && (2477 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_8_io_in_control_0_shift_b <=( _mesh_30_8_io_out_control_0_shift) ^ ((fiEnable && (2478 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_8_io_in_control_0_dataflow_b <=( _mesh_30_8_io_out_control_0_dataflow) ^ ((fiEnable && (2479 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_8_io_in_control_0_propagate_b <=( _mesh_30_8_io_out_control_0_propagate) ^ ((fiEnable && (2480 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_9_0) begin
			b_288_0 <=( io_in_b_9_0) ^ ((fiEnable && (2481 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1312_0 <=( io_in_d_9_0) ^ ((fiEnable && (2482 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_9_io_in_control_0_shift_b <=( io_in_control_9_0_shift) ^ ((fiEnable && (2483 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_9_io_in_control_0_dataflow_b <=( io_in_control_9_0_dataflow) ^ ((fiEnable && (2484 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_9_io_in_control_0_propagate_b <=( io_in_control_9_0_propagate) ^ ((fiEnable && (2485 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_9_io_out_valid_0) begin
			b_289_0 <=( _mesh_0_9_io_out_b_0) ^ ((fiEnable && (2486 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1313_0 <=( _mesh_0_9_io_out_c_0) ^ ((fiEnable && (2487 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_9_io_in_control_0_shift_b <=( _mesh_0_9_io_out_control_0_shift) ^ ((fiEnable && (2488 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_9_io_in_control_0_dataflow_b <=( _mesh_0_9_io_out_control_0_dataflow) ^ ((fiEnable && (2489 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_9_io_in_control_0_propagate_b <=( _mesh_0_9_io_out_control_0_propagate) ^ ((fiEnable && (2490 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_9_io_out_valid_0) begin
			b_290_0 <=( _mesh_1_9_io_out_b_0) ^ ((fiEnable && (2491 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1314_0 <=( _mesh_1_9_io_out_c_0) ^ ((fiEnable && (2492 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_9_io_in_control_0_shift_b <=( _mesh_1_9_io_out_control_0_shift) ^ ((fiEnable && (2493 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_9_io_in_control_0_dataflow_b <=( _mesh_1_9_io_out_control_0_dataflow) ^ ((fiEnable && (2494 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_9_io_in_control_0_propagate_b <=( _mesh_1_9_io_out_control_0_propagate) ^ ((fiEnable && (2495 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_9_io_out_valid_0) begin
			b_291_0 <=( _mesh_2_9_io_out_b_0) ^ ((fiEnable && (2496 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1315_0 <=( _mesh_2_9_io_out_c_0) ^ ((fiEnable && (2497 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_9_io_in_control_0_shift_b <=( _mesh_2_9_io_out_control_0_shift) ^ ((fiEnable && (2498 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_9_io_in_control_0_dataflow_b <=( _mesh_2_9_io_out_control_0_dataflow) ^ ((fiEnable && (2499 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_9_io_in_control_0_propagate_b <=( _mesh_2_9_io_out_control_0_propagate) ^ ((fiEnable && (2500 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_9_io_out_valid_0) begin
			b_292_0 <=( _mesh_3_9_io_out_b_0) ^ ((fiEnable && (2501 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1316_0 <=( _mesh_3_9_io_out_c_0) ^ ((fiEnable && (2502 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_9_io_in_control_0_shift_b <=( _mesh_3_9_io_out_control_0_shift) ^ ((fiEnable && (2503 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_9_io_in_control_0_dataflow_b <=( _mesh_3_9_io_out_control_0_dataflow) ^ ((fiEnable && (2504 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_9_io_in_control_0_propagate_b <=( _mesh_3_9_io_out_control_0_propagate) ^ ((fiEnable && (2505 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_9_io_out_valid_0) begin
			b_293_0 <=( _mesh_4_9_io_out_b_0) ^ ((fiEnable && (2506 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1317_0 <=( _mesh_4_9_io_out_c_0) ^ ((fiEnable && (2507 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_9_io_in_control_0_shift_b <=( _mesh_4_9_io_out_control_0_shift) ^ ((fiEnable && (2508 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_9_io_in_control_0_dataflow_b <=( _mesh_4_9_io_out_control_0_dataflow) ^ ((fiEnable && (2509 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_9_io_in_control_0_propagate_b <=( _mesh_4_9_io_out_control_0_propagate) ^ ((fiEnable && (2510 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_9_io_out_valid_0) begin
			b_294_0 <=( _mesh_5_9_io_out_b_0) ^ ((fiEnable && (2511 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1318_0 <=( _mesh_5_9_io_out_c_0) ^ ((fiEnable && (2512 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_9_io_in_control_0_shift_b <=( _mesh_5_9_io_out_control_0_shift) ^ ((fiEnable && (2513 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_9_io_in_control_0_dataflow_b <=( _mesh_5_9_io_out_control_0_dataflow) ^ ((fiEnable && (2514 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_9_io_in_control_0_propagate_b <=( _mesh_5_9_io_out_control_0_propagate) ^ ((fiEnable && (2515 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_9_io_out_valid_0) begin
			b_295_0 <=( _mesh_6_9_io_out_b_0) ^ ((fiEnable && (2516 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1319_0 <=( _mesh_6_9_io_out_c_0) ^ ((fiEnable && (2517 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_9_io_in_control_0_shift_b <=( _mesh_6_9_io_out_control_0_shift) ^ ((fiEnable && (2518 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_9_io_in_control_0_dataflow_b <=( _mesh_6_9_io_out_control_0_dataflow) ^ ((fiEnable && (2519 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_9_io_in_control_0_propagate_b <=( _mesh_6_9_io_out_control_0_propagate) ^ ((fiEnable && (2520 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_9_io_out_valid_0) begin
			b_296_0 <=( _mesh_7_9_io_out_b_0) ^ ((fiEnable && (2521 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1320_0 <=( _mesh_7_9_io_out_c_0) ^ ((fiEnable && (2522 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_9_io_in_control_0_shift_b <=( _mesh_7_9_io_out_control_0_shift) ^ ((fiEnable && (2523 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_9_io_in_control_0_dataflow_b <=( _mesh_7_9_io_out_control_0_dataflow) ^ ((fiEnable && (2524 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_9_io_in_control_0_propagate_b <=( _mesh_7_9_io_out_control_0_propagate) ^ ((fiEnable && (2525 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_9_io_out_valid_0) begin
			b_297_0 <=( _mesh_8_9_io_out_b_0) ^ ((fiEnable && (2526 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1321_0 <=( _mesh_8_9_io_out_c_0) ^ ((fiEnable && (2527 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_9_io_in_control_0_shift_b <=( _mesh_8_9_io_out_control_0_shift) ^ ((fiEnable && (2528 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_9_io_in_control_0_dataflow_b <=( _mesh_8_9_io_out_control_0_dataflow) ^ ((fiEnable && (2529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_9_io_in_control_0_propagate_b <=( _mesh_8_9_io_out_control_0_propagate) ^ ((fiEnable && (2530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_9_io_out_valid_0) begin
			b_298_0 <=( _mesh_9_9_io_out_b_0) ^ ((fiEnable && (2531 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1322_0 <=( _mesh_9_9_io_out_c_0) ^ ((fiEnable && (2532 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_9_io_in_control_0_shift_b <=( _mesh_9_9_io_out_control_0_shift) ^ ((fiEnable && (2533 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_9_io_in_control_0_dataflow_b <=( _mesh_9_9_io_out_control_0_dataflow) ^ ((fiEnable && (2534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_9_io_in_control_0_propagate_b <=( _mesh_9_9_io_out_control_0_propagate) ^ ((fiEnable && (2535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_9_io_out_valid_0) begin
			b_299_0 <=( _mesh_10_9_io_out_b_0) ^ ((fiEnable && (2536 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1323_0 <=( _mesh_10_9_io_out_c_0) ^ ((fiEnable && (2537 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_9_io_in_control_0_shift_b <=( _mesh_10_9_io_out_control_0_shift) ^ ((fiEnable && (2538 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_9_io_in_control_0_dataflow_b <=( _mesh_10_9_io_out_control_0_dataflow) ^ ((fiEnable && (2539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_9_io_in_control_0_propagate_b <=( _mesh_10_9_io_out_control_0_propagate) ^ ((fiEnable && (2540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_9_io_out_valid_0) begin
			b_300_0 <=( _mesh_11_9_io_out_b_0) ^ ((fiEnable && (2541 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1324_0 <=( _mesh_11_9_io_out_c_0) ^ ((fiEnable && (2542 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_9_io_in_control_0_shift_b <=( _mesh_11_9_io_out_control_0_shift) ^ ((fiEnable && (2543 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_9_io_in_control_0_dataflow_b <=( _mesh_11_9_io_out_control_0_dataflow) ^ ((fiEnable && (2544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_9_io_in_control_0_propagate_b <=( _mesh_11_9_io_out_control_0_propagate) ^ ((fiEnable && (2545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_9_io_out_valid_0) begin
			b_301_0 <=( _mesh_12_9_io_out_b_0) ^ ((fiEnable && (2546 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1325_0 <=( _mesh_12_9_io_out_c_0) ^ ((fiEnable && (2547 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_9_io_in_control_0_shift_b <=( _mesh_12_9_io_out_control_0_shift) ^ ((fiEnable && (2548 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_9_io_in_control_0_dataflow_b <=( _mesh_12_9_io_out_control_0_dataflow) ^ ((fiEnable && (2549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_9_io_in_control_0_propagate_b <=( _mesh_12_9_io_out_control_0_propagate) ^ ((fiEnable && (2550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_9_io_out_valid_0) begin
			b_302_0 <=( _mesh_13_9_io_out_b_0) ^ ((fiEnable && (2551 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1326_0 <=( _mesh_13_9_io_out_c_0) ^ ((fiEnable && (2552 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_9_io_in_control_0_shift_b <=( _mesh_13_9_io_out_control_0_shift) ^ ((fiEnable && (2553 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_9_io_in_control_0_dataflow_b <=( _mesh_13_9_io_out_control_0_dataflow) ^ ((fiEnable && (2554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_9_io_in_control_0_propagate_b <=( _mesh_13_9_io_out_control_0_propagate) ^ ((fiEnable && (2555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_9_io_out_valid_0) begin
			b_303_0 <=( _mesh_14_9_io_out_b_0) ^ ((fiEnable && (2556 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1327_0 <=( _mesh_14_9_io_out_c_0) ^ ((fiEnable && (2557 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_9_io_in_control_0_shift_b <=( _mesh_14_9_io_out_control_0_shift) ^ ((fiEnable && (2558 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_9_io_in_control_0_dataflow_b <=( _mesh_14_9_io_out_control_0_dataflow) ^ ((fiEnable && (2559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_9_io_in_control_0_propagate_b <=( _mesh_14_9_io_out_control_0_propagate) ^ ((fiEnable && (2560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_9_io_out_valid_0) begin
			b_304_0 <=( _mesh_15_9_io_out_b_0) ^ ((fiEnable && (2561 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1328_0 <=( _mesh_15_9_io_out_c_0) ^ ((fiEnable && (2562 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_9_io_in_control_0_shift_b <=( _mesh_15_9_io_out_control_0_shift) ^ ((fiEnable && (2563 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_9_io_in_control_0_dataflow_b <=( _mesh_15_9_io_out_control_0_dataflow) ^ ((fiEnable && (2564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_9_io_in_control_0_propagate_b <=( _mesh_15_9_io_out_control_0_propagate) ^ ((fiEnable && (2565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_9_io_out_valid_0) begin
			b_305_0 <=( _mesh_16_9_io_out_b_0) ^ ((fiEnable && (2566 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1329_0 <=( _mesh_16_9_io_out_c_0) ^ ((fiEnable && (2567 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_9_io_in_control_0_shift_b <=( _mesh_16_9_io_out_control_0_shift) ^ ((fiEnable && (2568 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_9_io_in_control_0_dataflow_b <=( _mesh_16_9_io_out_control_0_dataflow) ^ ((fiEnable && (2569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_9_io_in_control_0_propagate_b <=( _mesh_16_9_io_out_control_0_propagate) ^ ((fiEnable && (2570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_9_io_out_valid_0) begin
			b_306_0 <=( _mesh_17_9_io_out_b_0) ^ ((fiEnable && (2571 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1330_0 <=( _mesh_17_9_io_out_c_0) ^ ((fiEnable && (2572 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_9_io_in_control_0_shift_b <=( _mesh_17_9_io_out_control_0_shift) ^ ((fiEnable && (2573 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_9_io_in_control_0_dataflow_b <=( _mesh_17_9_io_out_control_0_dataflow) ^ ((fiEnable && (2574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_9_io_in_control_0_propagate_b <=( _mesh_17_9_io_out_control_0_propagate) ^ ((fiEnable && (2575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_9_io_out_valid_0) begin
			b_307_0 <=( _mesh_18_9_io_out_b_0) ^ ((fiEnable && (2576 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1331_0 <=( _mesh_18_9_io_out_c_0) ^ ((fiEnable && (2577 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_9_io_in_control_0_shift_b <=( _mesh_18_9_io_out_control_0_shift) ^ ((fiEnable && (2578 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_9_io_in_control_0_dataflow_b <=( _mesh_18_9_io_out_control_0_dataflow) ^ ((fiEnable && (2579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_9_io_in_control_0_propagate_b <=( _mesh_18_9_io_out_control_0_propagate) ^ ((fiEnable && (2580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_9_io_out_valid_0) begin
			b_308_0 <=( _mesh_19_9_io_out_b_0) ^ ((fiEnable && (2581 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1332_0 <=( _mesh_19_9_io_out_c_0) ^ ((fiEnable && (2582 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_9_io_in_control_0_shift_b <=( _mesh_19_9_io_out_control_0_shift) ^ ((fiEnable && (2583 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_9_io_in_control_0_dataflow_b <=( _mesh_19_9_io_out_control_0_dataflow) ^ ((fiEnable && (2584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_9_io_in_control_0_propagate_b <=( _mesh_19_9_io_out_control_0_propagate) ^ ((fiEnable && (2585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_9_io_out_valid_0) begin
			b_309_0 <=( _mesh_20_9_io_out_b_0) ^ ((fiEnable && (2586 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1333_0 <=( _mesh_20_9_io_out_c_0) ^ ((fiEnable && (2587 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_9_io_in_control_0_shift_b <=( _mesh_20_9_io_out_control_0_shift) ^ ((fiEnable && (2588 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_9_io_in_control_0_dataflow_b <=( _mesh_20_9_io_out_control_0_dataflow) ^ ((fiEnable && (2589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_9_io_in_control_0_propagate_b <=( _mesh_20_9_io_out_control_0_propagate) ^ ((fiEnable && (2590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_9_io_out_valid_0) begin
			b_310_0 <=( _mesh_21_9_io_out_b_0) ^ ((fiEnable && (2591 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1334_0 <=( _mesh_21_9_io_out_c_0) ^ ((fiEnable && (2592 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_9_io_in_control_0_shift_b <=( _mesh_21_9_io_out_control_0_shift) ^ ((fiEnable && (2593 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_9_io_in_control_0_dataflow_b <=( _mesh_21_9_io_out_control_0_dataflow) ^ ((fiEnable && (2594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_9_io_in_control_0_propagate_b <=( _mesh_21_9_io_out_control_0_propagate) ^ ((fiEnable && (2595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_9_io_out_valid_0) begin
			b_311_0 <=( _mesh_22_9_io_out_b_0) ^ ((fiEnable && (2596 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1335_0 <=( _mesh_22_9_io_out_c_0) ^ ((fiEnable && (2597 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_9_io_in_control_0_shift_b <=( _mesh_22_9_io_out_control_0_shift) ^ ((fiEnable && (2598 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_9_io_in_control_0_dataflow_b <=( _mesh_22_9_io_out_control_0_dataflow) ^ ((fiEnable && (2599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_9_io_in_control_0_propagate_b <=( _mesh_22_9_io_out_control_0_propagate) ^ ((fiEnable && (2600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_9_io_out_valid_0) begin
			b_312_0 <=( _mesh_23_9_io_out_b_0) ^ ((fiEnable && (2601 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1336_0 <=( _mesh_23_9_io_out_c_0) ^ ((fiEnable && (2602 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_9_io_in_control_0_shift_b <=( _mesh_23_9_io_out_control_0_shift) ^ ((fiEnable && (2603 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_9_io_in_control_0_dataflow_b <=( _mesh_23_9_io_out_control_0_dataflow) ^ ((fiEnable && (2604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_9_io_in_control_0_propagate_b <=( _mesh_23_9_io_out_control_0_propagate) ^ ((fiEnable && (2605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_9_io_out_valid_0) begin
			b_313_0 <=( _mesh_24_9_io_out_b_0) ^ ((fiEnable && (2606 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1337_0 <=( _mesh_24_9_io_out_c_0) ^ ((fiEnable && (2607 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_9_io_in_control_0_shift_b <=( _mesh_24_9_io_out_control_0_shift) ^ ((fiEnable && (2608 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_9_io_in_control_0_dataflow_b <=( _mesh_24_9_io_out_control_0_dataflow) ^ ((fiEnable && (2609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_9_io_in_control_0_propagate_b <=( _mesh_24_9_io_out_control_0_propagate) ^ ((fiEnable && (2610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_9_io_out_valid_0) begin
			b_314_0 <=( _mesh_25_9_io_out_b_0) ^ ((fiEnable && (2611 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1338_0 <=( _mesh_25_9_io_out_c_0) ^ ((fiEnable && (2612 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_9_io_in_control_0_shift_b <=( _mesh_25_9_io_out_control_0_shift) ^ ((fiEnable && (2613 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_9_io_in_control_0_dataflow_b <=( _mesh_25_9_io_out_control_0_dataflow) ^ ((fiEnable && (2614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_9_io_in_control_0_propagate_b <=( _mesh_25_9_io_out_control_0_propagate) ^ ((fiEnable && (2615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_9_io_out_valid_0) begin
			b_315_0 <=( _mesh_26_9_io_out_b_0) ^ ((fiEnable && (2616 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1339_0 <=( _mesh_26_9_io_out_c_0) ^ ((fiEnable && (2617 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_9_io_in_control_0_shift_b <=( _mesh_26_9_io_out_control_0_shift) ^ ((fiEnable && (2618 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_9_io_in_control_0_dataflow_b <=( _mesh_26_9_io_out_control_0_dataflow) ^ ((fiEnable && (2619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_9_io_in_control_0_propagate_b <=( _mesh_26_9_io_out_control_0_propagate) ^ ((fiEnable && (2620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_9_io_out_valid_0) begin
			b_316_0 <=( _mesh_27_9_io_out_b_0) ^ ((fiEnable && (2621 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1340_0 <=( _mesh_27_9_io_out_c_0) ^ ((fiEnable && (2622 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_9_io_in_control_0_shift_b <=( _mesh_27_9_io_out_control_0_shift) ^ ((fiEnable && (2623 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_9_io_in_control_0_dataflow_b <=( _mesh_27_9_io_out_control_0_dataflow) ^ ((fiEnable && (2624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_9_io_in_control_0_propagate_b <=( _mesh_27_9_io_out_control_0_propagate) ^ ((fiEnable && (2625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_9_io_out_valid_0) begin
			b_317_0 <=( _mesh_28_9_io_out_b_0) ^ ((fiEnable && (2626 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1341_0 <=( _mesh_28_9_io_out_c_0) ^ ((fiEnable && (2627 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_9_io_in_control_0_shift_b <=( _mesh_28_9_io_out_control_0_shift) ^ ((fiEnable && (2628 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_9_io_in_control_0_dataflow_b <=( _mesh_28_9_io_out_control_0_dataflow) ^ ((fiEnable && (2629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_9_io_in_control_0_propagate_b <=( _mesh_28_9_io_out_control_0_propagate) ^ ((fiEnable && (2630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_9_io_out_valid_0) begin
			b_318_0 <=( _mesh_29_9_io_out_b_0) ^ ((fiEnable && (2631 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1342_0 <=( _mesh_29_9_io_out_c_0) ^ ((fiEnable && (2632 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_9_io_in_control_0_shift_b <=( _mesh_29_9_io_out_control_0_shift) ^ ((fiEnable && (2633 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_9_io_in_control_0_dataflow_b <=( _mesh_29_9_io_out_control_0_dataflow) ^ ((fiEnable && (2634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_9_io_in_control_0_propagate_b <=( _mesh_29_9_io_out_control_0_propagate) ^ ((fiEnable && (2635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_9_io_out_valid_0) begin
			b_319_0 <=( _mesh_30_9_io_out_b_0) ^ ((fiEnable && (2636 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1343_0 <=( _mesh_30_9_io_out_c_0) ^ ((fiEnable && (2637 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_9_io_in_control_0_shift_b <=( _mesh_30_9_io_out_control_0_shift) ^ ((fiEnable && (2638 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_9_io_in_control_0_dataflow_b <=( _mesh_30_9_io_out_control_0_dataflow) ^ ((fiEnable && (2639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_9_io_in_control_0_propagate_b <=( _mesh_30_9_io_out_control_0_propagate) ^ ((fiEnable && (2640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_10_0) begin
			b_320_0 <=( io_in_b_10_0) ^ ((fiEnable && (2641 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1344_0 <=( io_in_d_10_0) ^ ((fiEnable && (2642 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_10_io_in_control_0_shift_b <=( io_in_control_10_0_shift) ^ ((fiEnable && (2643 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_10_io_in_control_0_dataflow_b <=( io_in_control_10_0_dataflow) ^ ((fiEnable && (2644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_10_io_in_control_0_propagate_b <=( io_in_control_10_0_propagate) ^ ((fiEnable && (2645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_10_io_out_valid_0) begin
			b_321_0 <=( _mesh_0_10_io_out_b_0) ^ ((fiEnable && (2646 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1345_0 <=( _mesh_0_10_io_out_c_0) ^ ((fiEnable && (2647 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_10_io_in_control_0_shift_b <=( _mesh_0_10_io_out_control_0_shift) ^ ((fiEnable && (2648 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_10_io_in_control_0_dataflow_b <=( _mesh_0_10_io_out_control_0_dataflow) ^ ((fiEnable && (2649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_10_io_in_control_0_propagate_b <=( _mesh_0_10_io_out_control_0_propagate) ^ ((fiEnable && (2650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_10_io_out_valid_0) begin
			b_322_0 <=( _mesh_1_10_io_out_b_0) ^ ((fiEnable && (2651 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1346_0 <=( _mesh_1_10_io_out_c_0) ^ ((fiEnable && (2652 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_10_io_in_control_0_shift_b <=( _mesh_1_10_io_out_control_0_shift) ^ ((fiEnable && (2653 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_10_io_in_control_0_dataflow_b <=( _mesh_1_10_io_out_control_0_dataflow) ^ ((fiEnable && (2654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_10_io_in_control_0_propagate_b <=( _mesh_1_10_io_out_control_0_propagate) ^ ((fiEnable && (2655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_10_io_out_valid_0) begin
			b_323_0 <=( _mesh_2_10_io_out_b_0) ^ ((fiEnable && (2656 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1347_0 <=( _mesh_2_10_io_out_c_0) ^ ((fiEnable && (2657 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_10_io_in_control_0_shift_b <=( _mesh_2_10_io_out_control_0_shift) ^ ((fiEnable && (2658 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_10_io_in_control_0_dataflow_b <=( _mesh_2_10_io_out_control_0_dataflow) ^ ((fiEnable && (2659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_10_io_in_control_0_propagate_b <=( _mesh_2_10_io_out_control_0_propagate) ^ ((fiEnable && (2660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_10_io_out_valid_0) begin
			b_324_0 <=( _mesh_3_10_io_out_b_0) ^ ((fiEnable && (2661 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1348_0 <=( _mesh_3_10_io_out_c_0) ^ ((fiEnable && (2662 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_10_io_in_control_0_shift_b <=( _mesh_3_10_io_out_control_0_shift) ^ ((fiEnable && (2663 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_10_io_in_control_0_dataflow_b <=( _mesh_3_10_io_out_control_0_dataflow) ^ ((fiEnable && (2664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_10_io_in_control_0_propagate_b <=( _mesh_3_10_io_out_control_0_propagate) ^ ((fiEnable && (2665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_10_io_out_valid_0) begin
			b_325_0 <=( _mesh_4_10_io_out_b_0) ^ ((fiEnable && (2666 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1349_0 <=( _mesh_4_10_io_out_c_0) ^ ((fiEnable && (2667 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_10_io_in_control_0_shift_b <=( _mesh_4_10_io_out_control_0_shift) ^ ((fiEnable && (2668 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_10_io_in_control_0_dataflow_b <=( _mesh_4_10_io_out_control_0_dataflow) ^ ((fiEnable && (2669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_10_io_in_control_0_propagate_b <=( _mesh_4_10_io_out_control_0_propagate) ^ ((fiEnable && (2670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_10_io_out_valid_0) begin
			b_326_0 <=( _mesh_5_10_io_out_b_0) ^ ((fiEnable && (2671 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1350_0 <=( _mesh_5_10_io_out_c_0) ^ ((fiEnable && (2672 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_10_io_in_control_0_shift_b <=( _mesh_5_10_io_out_control_0_shift) ^ ((fiEnable && (2673 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_10_io_in_control_0_dataflow_b <=( _mesh_5_10_io_out_control_0_dataflow) ^ ((fiEnable && (2674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_10_io_in_control_0_propagate_b <=( _mesh_5_10_io_out_control_0_propagate) ^ ((fiEnable && (2675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_10_io_out_valid_0) begin
			b_327_0 <=( _mesh_6_10_io_out_b_0) ^ ((fiEnable && (2676 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1351_0 <=( _mesh_6_10_io_out_c_0) ^ ((fiEnable && (2677 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_10_io_in_control_0_shift_b <=( _mesh_6_10_io_out_control_0_shift) ^ ((fiEnable && (2678 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_10_io_in_control_0_dataflow_b <=( _mesh_6_10_io_out_control_0_dataflow) ^ ((fiEnable && (2679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_10_io_in_control_0_propagate_b <=( _mesh_6_10_io_out_control_0_propagate) ^ ((fiEnable && (2680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_10_io_out_valid_0) begin
			b_328_0 <=( _mesh_7_10_io_out_b_0) ^ ((fiEnable && (2681 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1352_0 <=( _mesh_7_10_io_out_c_0) ^ ((fiEnable && (2682 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_10_io_in_control_0_shift_b <=( _mesh_7_10_io_out_control_0_shift) ^ ((fiEnable && (2683 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_10_io_in_control_0_dataflow_b <=( _mesh_7_10_io_out_control_0_dataflow) ^ ((fiEnable && (2684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_10_io_in_control_0_propagate_b <=( _mesh_7_10_io_out_control_0_propagate) ^ ((fiEnable && (2685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_10_io_out_valid_0) begin
			b_329_0 <=( _mesh_8_10_io_out_b_0) ^ ((fiEnable && (2686 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1353_0 <=( _mesh_8_10_io_out_c_0) ^ ((fiEnable && (2687 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_10_io_in_control_0_shift_b <=( _mesh_8_10_io_out_control_0_shift) ^ ((fiEnable && (2688 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_10_io_in_control_0_dataflow_b <=( _mesh_8_10_io_out_control_0_dataflow) ^ ((fiEnable && (2689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_10_io_in_control_0_propagate_b <=( _mesh_8_10_io_out_control_0_propagate) ^ ((fiEnable && (2690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_10_io_out_valid_0) begin
			b_330_0 <=( _mesh_9_10_io_out_b_0) ^ ((fiEnable && (2691 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1354_0 <=( _mesh_9_10_io_out_c_0) ^ ((fiEnable && (2692 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_10_io_in_control_0_shift_b <=( _mesh_9_10_io_out_control_0_shift) ^ ((fiEnable && (2693 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_10_io_in_control_0_dataflow_b <=( _mesh_9_10_io_out_control_0_dataflow) ^ ((fiEnable && (2694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_10_io_in_control_0_propagate_b <=( _mesh_9_10_io_out_control_0_propagate) ^ ((fiEnable && (2695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_10_io_out_valid_0) begin
			b_331_0 <=( _mesh_10_10_io_out_b_0) ^ ((fiEnable && (2696 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1355_0 <=( _mesh_10_10_io_out_c_0) ^ ((fiEnable && (2697 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_10_io_in_control_0_shift_b <=( _mesh_10_10_io_out_control_0_shift) ^ ((fiEnable && (2698 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_10_io_in_control_0_dataflow_b <=( _mesh_10_10_io_out_control_0_dataflow) ^ ((fiEnable && (2699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_10_io_in_control_0_propagate_b <=( _mesh_10_10_io_out_control_0_propagate) ^ ((fiEnable && (2700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_10_io_out_valid_0) begin
			b_332_0 <=( _mesh_11_10_io_out_b_0) ^ ((fiEnable && (2701 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1356_0 <=( _mesh_11_10_io_out_c_0) ^ ((fiEnable && (2702 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_10_io_in_control_0_shift_b <=( _mesh_11_10_io_out_control_0_shift) ^ ((fiEnable && (2703 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_10_io_in_control_0_dataflow_b <=( _mesh_11_10_io_out_control_0_dataflow) ^ ((fiEnable && (2704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_10_io_in_control_0_propagate_b <=( _mesh_11_10_io_out_control_0_propagate) ^ ((fiEnable && (2705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_10_io_out_valid_0) begin
			b_333_0 <=( _mesh_12_10_io_out_b_0) ^ ((fiEnable && (2706 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1357_0 <=( _mesh_12_10_io_out_c_0) ^ ((fiEnable && (2707 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_10_io_in_control_0_shift_b <=( _mesh_12_10_io_out_control_0_shift) ^ ((fiEnable && (2708 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_10_io_in_control_0_dataflow_b <=( _mesh_12_10_io_out_control_0_dataflow) ^ ((fiEnable && (2709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_10_io_in_control_0_propagate_b <=( _mesh_12_10_io_out_control_0_propagate) ^ ((fiEnable && (2710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_10_io_out_valid_0) begin
			b_334_0 <=( _mesh_13_10_io_out_b_0) ^ ((fiEnable && (2711 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1358_0 <=( _mesh_13_10_io_out_c_0) ^ ((fiEnable && (2712 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_10_io_in_control_0_shift_b <=( _mesh_13_10_io_out_control_0_shift) ^ ((fiEnable && (2713 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_10_io_in_control_0_dataflow_b <=( _mesh_13_10_io_out_control_0_dataflow) ^ ((fiEnable && (2714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_10_io_in_control_0_propagate_b <=( _mesh_13_10_io_out_control_0_propagate) ^ ((fiEnable && (2715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_10_io_out_valid_0) begin
			b_335_0 <=( _mesh_14_10_io_out_b_0) ^ ((fiEnable && (2716 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1359_0 <=( _mesh_14_10_io_out_c_0) ^ ((fiEnable && (2717 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_10_io_in_control_0_shift_b <=( _mesh_14_10_io_out_control_0_shift) ^ ((fiEnable && (2718 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_10_io_in_control_0_dataflow_b <=( _mesh_14_10_io_out_control_0_dataflow) ^ ((fiEnable && (2719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_10_io_in_control_0_propagate_b <=( _mesh_14_10_io_out_control_0_propagate) ^ ((fiEnable && (2720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_10_io_out_valid_0) begin
			b_336_0 <=( _mesh_15_10_io_out_b_0) ^ ((fiEnable && (2721 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1360_0 <=( _mesh_15_10_io_out_c_0) ^ ((fiEnable && (2722 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_10_io_in_control_0_shift_b <=( _mesh_15_10_io_out_control_0_shift) ^ ((fiEnable && (2723 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_10_io_in_control_0_dataflow_b <=( _mesh_15_10_io_out_control_0_dataflow) ^ ((fiEnable && (2724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_10_io_in_control_0_propagate_b <=( _mesh_15_10_io_out_control_0_propagate) ^ ((fiEnable && (2725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_10_io_out_valid_0) begin
			b_337_0 <=( _mesh_16_10_io_out_b_0) ^ ((fiEnable && (2726 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1361_0 <=( _mesh_16_10_io_out_c_0) ^ ((fiEnable && (2727 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_10_io_in_control_0_shift_b <=( _mesh_16_10_io_out_control_0_shift) ^ ((fiEnable && (2728 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_10_io_in_control_0_dataflow_b <=( _mesh_16_10_io_out_control_0_dataflow) ^ ((fiEnable && (2729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_10_io_in_control_0_propagate_b <=( _mesh_16_10_io_out_control_0_propagate) ^ ((fiEnable && (2730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_10_io_out_valid_0) begin
			b_338_0 <=( _mesh_17_10_io_out_b_0) ^ ((fiEnable && (2731 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1362_0 <=( _mesh_17_10_io_out_c_0) ^ ((fiEnable && (2732 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_10_io_in_control_0_shift_b <=( _mesh_17_10_io_out_control_0_shift) ^ ((fiEnable && (2733 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_10_io_in_control_0_dataflow_b <=( _mesh_17_10_io_out_control_0_dataflow) ^ ((fiEnable && (2734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_10_io_in_control_0_propagate_b <=( _mesh_17_10_io_out_control_0_propagate) ^ ((fiEnable && (2735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_10_io_out_valid_0) begin
			b_339_0 <=( _mesh_18_10_io_out_b_0) ^ ((fiEnable && (2736 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1363_0 <=( _mesh_18_10_io_out_c_0) ^ ((fiEnable && (2737 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_10_io_in_control_0_shift_b <=( _mesh_18_10_io_out_control_0_shift) ^ ((fiEnable && (2738 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_10_io_in_control_0_dataflow_b <=( _mesh_18_10_io_out_control_0_dataflow) ^ ((fiEnable && (2739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_10_io_in_control_0_propagate_b <=( _mesh_18_10_io_out_control_0_propagate) ^ ((fiEnable && (2740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_10_io_out_valid_0) begin
			b_340_0 <=( _mesh_19_10_io_out_b_0) ^ ((fiEnable && (2741 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1364_0 <=( _mesh_19_10_io_out_c_0) ^ ((fiEnable && (2742 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_10_io_in_control_0_shift_b <=( _mesh_19_10_io_out_control_0_shift) ^ ((fiEnable && (2743 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_10_io_in_control_0_dataflow_b <=( _mesh_19_10_io_out_control_0_dataflow) ^ ((fiEnable && (2744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_10_io_in_control_0_propagate_b <=( _mesh_19_10_io_out_control_0_propagate) ^ ((fiEnable && (2745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_10_io_out_valid_0) begin
			b_341_0 <=( _mesh_20_10_io_out_b_0) ^ ((fiEnable && (2746 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1365_0 <=( _mesh_20_10_io_out_c_0) ^ ((fiEnable && (2747 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_10_io_in_control_0_shift_b <=( _mesh_20_10_io_out_control_0_shift) ^ ((fiEnable && (2748 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_10_io_in_control_0_dataflow_b <=( _mesh_20_10_io_out_control_0_dataflow) ^ ((fiEnable && (2749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_10_io_in_control_0_propagate_b <=( _mesh_20_10_io_out_control_0_propagate) ^ ((fiEnable && (2750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_10_io_out_valid_0) begin
			b_342_0 <=( _mesh_21_10_io_out_b_0) ^ ((fiEnable && (2751 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1366_0 <=( _mesh_21_10_io_out_c_0) ^ ((fiEnable && (2752 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_10_io_in_control_0_shift_b <=( _mesh_21_10_io_out_control_0_shift) ^ ((fiEnable && (2753 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_10_io_in_control_0_dataflow_b <=( _mesh_21_10_io_out_control_0_dataflow) ^ ((fiEnable && (2754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_10_io_in_control_0_propagate_b <=( _mesh_21_10_io_out_control_0_propagate) ^ ((fiEnable && (2755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_10_io_out_valid_0) begin
			b_343_0 <=( _mesh_22_10_io_out_b_0) ^ ((fiEnable && (2756 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1367_0 <=( _mesh_22_10_io_out_c_0) ^ ((fiEnable && (2757 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_10_io_in_control_0_shift_b <=( _mesh_22_10_io_out_control_0_shift) ^ ((fiEnable && (2758 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_10_io_in_control_0_dataflow_b <=( _mesh_22_10_io_out_control_0_dataflow) ^ ((fiEnable && (2759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_10_io_in_control_0_propagate_b <=( _mesh_22_10_io_out_control_0_propagate) ^ ((fiEnable && (2760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_10_io_out_valid_0) begin
			b_344_0 <=( _mesh_23_10_io_out_b_0) ^ ((fiEnable && (2761 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1368_0 <=( _mesh_23_10_io_out_c_0) ^ ((fiEnable && (2762 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_10_io_in_control_0_shift_b <=( _mesh_23_10_io_out_control_0_shift) ^ ((fiEnable && (2763 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_10_io_in_control_0_dataflow_b <=( _mesh_23_10_io_out_control_0_dataflow) ^ ((fiEnable && (2764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_10_io_in_control_0_propagate_b <=( _mesh_23_10_io_out_control_0_propagate) ^ ((fiEnable && (2765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_10_io_out_valid_0) begin
			b_345_0 <=( _mesh_24_10_io_out_b_0) ^ ((fiEnable && (2766 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1369_0 <=( _mesh_24_10_io_out_c_0) ^ ((fiEnable && (2767 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_10_io_in_control_0_shift_b <=( _mesh_24_10_io_out_control_0_shift) ^ ((fiEnable && (2768 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_10_io_in_control_0_dataflow_b <=( _mesh_24_10_io_out_control_0_dataflow) ^ ((fiEnable && (2769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_10_io_in_control_0_propagate_b <=( _mesh_24_10_io_out_control_0_propagate) ^ ((fiEnable && (2770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_10_io_out_valid_0) begin
			b_346_0 <=( _mesh_25_10_io_out_b_0) ^ ((fiEnable && (2771 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1370_0 <=( _mesh_25_10_io_out_c_0) ^ ((fiEnable && (2772 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_10_io_in_control_0_shift_b <=( _mesh_25_10_io_out_control_0_shift) ^ ((fiEnable && (2773 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_10_io_in_control_0_dataflow_b <=( _mesh_25_10_io_out_control_0_dataflow) ^ ((fiEnable && (2774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_10_io_in_control_0_propagate_b <=( _mesh_25_10_io_out_control_0_propagate) ^ ((fiEnable && (2775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_10_io_out_valid_0) begin
			b_347_0 <=( _mesh_26_10_io_out_b_0) ^ ((fiEnable && (2776 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1371_0 <=( _mesh_26_10_io_out_c_0) ^ ((fiEnable && (2777 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_10_io_in_control_0_shift_b <=( _mesh_26_10_io_out_control_0_shift) ^ ((fiEnable && (2778 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_10_io_in_control_0_dataflow_b <=( _mesh_26_10_io_out_control_0_dataflow) ^ ((fiEnable && (2779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_10_io_in_control_0_propagate_b <=( _mesh_26_10_io_out_control_0_propagate) ^ ((fiEnable && (2780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_10_io_out_valid_0) begin
			b_348_0 <=( _mesh_27_10_io_out_b_0) ^ ((fiEnable && (2781 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1372_0 <=( _mesh_27_10_io_out_c_0) ^ ((fiEnable && (2782 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_10_io_in_control_0_shift_b <=( _mesh_27_10_io_out_control_0_shift) ^ ((fiEnable && (2783 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_10_io_in_control_0_dataflow_b <=( _mesh_27_10_io_out_control_0_dataflow) ^ ((fiEnable && (2784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_10_io_in_control_0_propagate_b <=( _mesh_27_10_io_out_control_0_propagate) ^ ((fiEnable && (2785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_10_io_out_valid_0) begin
			b_349_0 <=( _mesh_28_10_io_out_b_0) ^ ((fiEnable && (2786 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1373_0 <=( _mesh_28_10_io_out_c_0) ^ ((fiEnable && (2787 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_10_io_in_control_0_shift_b <=( _mesh_28_10_io_out_control_0_shift) ^ ((fiEnable && (2788 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_10_io_in_control_0_dataflow_b <=( _mesh_28_10_io_out_control_0_dataflow) ^ ((fiEnable && (2789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_10_io_in_control_0_propagate_b <=( _mesh_28_10_io_out_control_0_propagate) ^ ((fiEnable && (2790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_10_io_out_valid_0) begin
			b_350_0 <=( _mesh_29_10_io_out_b_0) ^ ((fiEnable && (2791 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1374_0 <=( _mesh_29_10_io_out_c_0) ^ ((fiEnable && (2792 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_10_io_in_control_0_shift_b <=( _mesh_29_10_io_out_control_0_shift) ^ ((fiEnable && (2793 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_10_io_in_control_0_dataflow_b <=( _mesh_29_10_io_out_control_0_dataflow) ^ ((fiEnable && (2794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_10_io_in_control_0_propagate_b <=( _mesh_29_10_io_out_control_0_propagate) ^ ((fiEnable && (2795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_10_io_out_valid_0) begin
			b_351_0 <=( _mesh_30_10_io_out_b_0) ^ ((fiEnable && (2796 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1375_0 <=( _mesh_30_10_io_out_c_0) ^ ((fiEnable && (2797 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_10_io_in_control_0_shift_b <=( _mesh_30_10_io_out_control_0_shift) ^ ((fiEnable && (2798 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_10_io_in_control_0_dataflow_b <=( _mesh_30_10_io_out_control_0_dataflow) ^ ((fiEnable && (2799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_10_io_in_control_0_propagate_b <=( _mesh_30_10_io_out_control_0_propagate) ^ ((fiEnable && (2800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_11_0) begin
			b_352_0 <=( io_in_b_11_0) ^ ((fiEnable && (2801 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1376_0 <=( io_in_d_11_0) ^ ((fiEnable && (2802 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_11_io_in_control_0_shift_b <=( io_in_control_11_0_shift) ^ ((fiEnable && (2803 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_11_io_in_control_0_dataflow_b <=( io_in_control_11_0_dataflow) ^ ((fiEnable && (2804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_11_io_in_control_0_propagate_b <=( io_in_control_11_0_propagate) ^ ((fiEnable && (2805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_11_io_out_valid_0) begin
			b_353_0 <=( _mesh_0_11_io_out_b_0) ^ ((fiEnable && (2806 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1377_0 <=( _mesh_0_11_io_out_c_0) ^ ((fiEnable && (2807 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_11_io_in_control_0_shift_b <=( _mesh_0_11_io_out_control_0_shift) ^ ((fiEnable && (2808 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_11_io_in_control_0_dataflow_b <=( _mesh_0_11_io_out_control_0_dataflow) ^ ((fiEnable && (2809 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_11_io_in_control_0_propagate_b <=( _mesh_0_11_io_out_control_0_propagate) ^ ((fiEnable && (2810 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_11_io_out_valid_0) begin
			b_354_0 <=( _mesh_1_11_io_out_b_0) ^ ((fiEnable && (2811 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1378_0 <=( _mesh_1_11_io_out_c_0) ^ ((fiEnable && (2812 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_11_io_in_control_0_shift_b <=( _mesh_1_11_io_out_control_0_shift) ^ ((fiEnable && (2813 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_11_io_in_control_0_dataflow_b <=( _mesh_1_11_io_out_control_0_dataflow) ^ ((fiEnable && (2814 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_11_io_in_control_0_propagate_b <=( _mesh_1_11_io_out_control_0_propagate) ^ ((fiEnable && (2815 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_11_io_out_valid_0) begin
			b_355_0 <=( _mesh_2_11_io_out_b_0) ^ ((fiEnable && (2816 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1379_0 <=( _mesh_2_11_io_out_c_0) ^ ((fiEnable && (2817 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_11_io_in_control_0_shift_b <=( _mesh_2_11_io_out_control_0_shift) ^ ((fiEnable && (2818 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_11_io_in_control_0_dataflow_b <=( _mesh_2_11_io_out_control_0_dataflow) ^ ((fiEnable && (2819 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_11_io_in_control_0_propagate_b <=( _mesh_2_11_io_out_control_0_propagate) ^ ((fiEnable && (2820 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_11_io_out_valid_0) begin
			b_356_0 <=( _mesh_3_11_io_out_b_0) ^ ((fiEnable && (2821 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1380_0 <=( _mesh_3_11_io_out_c_0) ^ ((fiEnable && (2822 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_11_io_in_control_0_shift_b <=( _mesh_3_11_io_out_control_0_shift) ^ ((fiEnable && (2823 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_11_io_in_control_0_dataflow_b <=( _mesh_3_11_io_out_control_0_dataflow) ^ ((fiEnable && (2824 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_11_io_in_control_0_propagate_b <=( _mesh_3_11_io_out_control_0_propagate) ^ ((fiEnable && (2825 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_11_io_out_valid_0) begin
			b_357_0 <=( _mesh_4_11_io_out_b_0) ^ ((fiEnable && (2826 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1381_0 <=( _mesh_4_11_io_out_c_0) ^ ((fiEnable && (2827 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_11_io_in_control_0_shift_b <=( _mesh_4_11_io_out_control_0_shift) ^ ((fiEnable && (2828 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_11_io_in_control_0_dataflow_b <=( _mesh_4_11_io_out_control_0_dataflow) ^ ((fiEnable && (2829 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_11_io_in_control_0_propagate_b <=( _mesh_4_11_io_out_control_0_propagate) ^ ((fiEnable && (2830 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_11_io_out_valid_0) begin
			b_358_0 <=( _mesh_5_11_io_out_b_0) ^ ((fiEnable && (2831 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1382_0 <=( _mesh_5_11_io_out_c_0) ^ ((fiEnable && (2832 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_11_io_in_control_0_shift_b <=( _mesh_5_11_io_out_control_0_shift) ^ ((fiEnable && (2833 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_11_io_in_control_0_dataflow_b <=( _mesh_5_11_io_out_control_0_dataflow) ^ ((fiEnable && (2834 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_11_io_in_control_0_propagate_b <=( _mesh_5_11_io_out_control_0_propagate) ^ ((fiEnable && (2835 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_11_io_out_valid_0) begin
			b_359_0 <=( _mesh_6_11_io_out_b_0) ^ ((fiEnable && (2836 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1383_0 <=( _mesh_6_11_io_out_c_0) ^ ((fiEnable && (2837 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_11_io_in_control_0_shift_b <=( _mesh_6_11_io_out_control_0_shift) ^ ((fiEnable && (2838 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_11_io_in_control_0_dataflow_b <=( _mesh_6_11_io_out_control_0_dataflow) ^ ((fiEnable && (2839 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_11_io_in_control_0_propagate_b <=( _mesh_6_11_io_out_control_0_propagate) ^ ((fiEnable && (2840 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_11_io_out_valid_0) begin
			b_360_0 <=( _mesh_7_11_io_out_b_0) ^ ((fiEnable && (2841 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1384_0 <=( _mesh_7_11_io_out_c_0) ^ ((fiEnable && (2842 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_11_io_in_control_0_shift_b <=( _mesh_7_11_io_out_control_0_shift) ^ ((fiEnable && (2843 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_11_io_in_control_0_dataflow_b <=( _mesh_7_11_io_out_control_0_dataflow) ^ ((fiEnable && (2844 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_11_io_in_control_0_propagate_b <=( _mesh_7_11_io_out_control_0_propagate) ^ ((fiEnable && (2845 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_11_io_out_valid_0) begin
			b_361_0 <=( _mesh_8_11_io_out_b_0) ^ ((fiEnable && (2846 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1385_0 <=( _mesh_8_11_io_out_c_0) ^ ((fiEnable && (2847 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_11_io_in_control_0_shift_b <=( _mesh_8_11_io_out_control_0_shift) ^ ((fiEnable && (2848 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_11_io_in_control_0_dataflow_b <=( _mesh_8_11_io_out_control_0_dataflow) ^ ((fiEnable && (2849 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_11_io_in_control_0_propagate_b <=( _mesh_8_11_io_out_control_0_propagate) ^ ((fiEnable && (2850 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_11_io_out_valid_0) begin
			b_362_0 <=( _mesh_9_11_io_out_b_0) ^ ((fiEnable && (2851 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1386_0 <=( _mesh_9_11_io_out_c_0) ^ ((fiEnable && (2852 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_11_io_in_control_0_shift_b <=( _mesh_9_11_io_out_control_0_shift) ^ ((fiEnable && (2853 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_11_io_in_control_0_dataflow_b <=( _mesh_9_11_io_out_control_0_dataflow) ^ ((fiEnable && (2854 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_11_io_in_control_0_propagate_b <=( _mesh_9_11_io_out_control_0_propagate) ^ ((fiEnable && (2855 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_11_io_out_valid_0) begin
			b_363_0 <=( _mesh_10_11_io_out_b_0) ^ ((fiEnable && (2856 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1387_0 <=( _mesh_10_11_io_out_c_0) ^ ((fiEnable && (2857 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_11_io_in_control_0_shift_b <=( _mesh_10_11_io_out_control_0_shift) ^ ((fiEnable && (2858 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_11_io_in_control_0_dataflow_b <=( _mesh_10_11_io_out_control_0_dataflow) ^ ((fiEnable && (2859 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_11_io_in_control_0_propagate_b <=( _mesh_10_11_io_out_control_0_propagate) ^ ((fiEnable && (2860 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_11_io_out_valid_0) begin
			b_364_0 <=( _mesh_11_11_io_out_b_0) ^ ((fiEnable && (2861 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1388_0 <=( _mesh_11_11_io_out_c_0) ^ ((fiEnable && (2862 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_11_io_in_control_0_shift_b <=( _mesh_11_11_io_out_control_0_shift) ^ ((fiEnable && (2863 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_11_io_in_control_0_dataflow_b <=( _mesh_11_11_io_out_control_0_dataflow) ^ ((fiEnable && (2864 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_11_io_in_control_0_propagate_b <=( _mesh_11_11_io_out_control_0_propagate) ^ ((fiEnable && (2865 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_11_io_out_valid_0) begin
			b_365_0 <=( _mesh_12_11_io_out_b_0) ^ ((fiEnable && (2866 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1389_0 <=( _mesh_12_11_io_out_c_0) ^ ((fiEnable && (2867 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_11_io_in_control_0_shift_b <=( _mesh_12_11_io_out_control_0_shift) ^ ((fiEnable && (2868 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_11_io_in_control_0_dataflow_b <=( _mesh_12_11_io_out_control_0_dataflow) ^ ((fiEnable && (2869 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_11_io_in_control_0_propagate_b <=( _mesh_12_11_io_out_control_0_propagate) ^ ((fiEnable && (2870 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_11_io_out_valid_0) begin
			b_366_0 <=( _mesh_13_11_io_out_b_0) ^ ((fiEnable && (2871 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1390_0 <=( _mesh_13_11_io_out_c_0) ^ ((fiEnable && (2872 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_11_io_in_control_0_shift_b <=( _mesh_13_11_io_out_control_0_shift) ^ ((fiEnable && (2873 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_11_io_in_control_0_dataflow_b <=( _mesh_13_11_io_out_control_0_dataflow) ^ ((fiEnable && (2874 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_11_io_in_control_0_propagate_b <=( _mesh_13_11_io_out_control_0_propagate) ^ ((fiEnable && (2875 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_11_io_out_valid_0) begin
			b_367_0 <=( _mesh_14_11_io_out_b_0) ^ ((fiEnable && (2876 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1391_0 <=( _mesh_14_11_io_out_c_0) ^ ((fiEnable && (2877 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_11_io_in_control_0_shift_b <=( _mesh_14_11_io_out_control_0_shift) ^ ((fiEnable && (2878 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_11_io_in_control_0_dataflow_b <=( _mesh_14_11_io_out_control_0_dataflow) ^ ((fiEnable && (2879 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_11_io_in_control_0_propagate_b <=( _mesh_14_11_io_out_control_0_propagate) ^ ((fiEnable && (2880 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_11_io_out_valid_0) begin
			b_368_0 <=( _mesh_15_11_io_out_b_0) ^ ((fiEnable && (2881 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1392_0 <=( _mesh_15_11_io_out_c_0) ^ ((fiEnable && (2882 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_11_io_in_control_0_shift_b <=( _mesh_15_11_io_out_control_0_shift) ^ ((fiEnable && (2883 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_11_io_in_control_0_dataflow_b <=( _mesh_15_11_io_out_control_0_dataflow) ^ ((fiEnable && (2884 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_11_io_in_control_0_propagate_b <=( _mesh_15_11_io_out_control_0_propagate) ^ ((fiEnable && (2885 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_11_io_out_valid_0) begin
			b_369_0 <=( _mesh_16_11_io_out_b_0) ^ ((fiEnable && (2886 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1393_0 <=( _mesh_16_11_io_out_c_0) ^ ((fiEnable && (2887 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_11_io_in_control_0_shift_b <=( _mesh_16_11_io_out_control_0_shift) ^ ((fiEnable && (2888 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_11_io_in_control_0_dataflow_b <=( _mesh_16_11_io_out_control_0_dataflow) ^ ((fiEnable && (2889 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_11_io_in_control_0_propagate_b <=( _mesh_16_11_io_out_control_0_propagate) ^ ((fiEnable && (2890 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_11_io_out_valid_0) begin
			b_370_0 <=( _mesh_17_11_io_out_b_0) ^ ((fiEnable && (2891 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1394_0 <=( _mesh_17_11_io_out_c_0) ^ ((fiEnable && (2892 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_11_io_in_control_0_shift_b <=( _mesh_17_11_io_out_control_0_shift) ^ ((fiEnable && (2893 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_11_io_in_control_0_dataflow_b <=( _mesh_17_11_io_out_control_0_dataflow) ^ ((fiEnable && (2894 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_11_io_in_control_0_propagate_b <=( _mesh_17_11_io_out_control_0_propagate) ^ ((fiEnable && (2895 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_11_io_out_valid_0) begin
			b_371_0 <=( _mesh_18_11_io_out_b_0) ^ ((fiEnable && (2896 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1395_0 <=( _mesh_18_11_io_out_c_0) ^ ((fiEnable && (2897 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_11_io_in_control_0_shift_b <=( _mesh_18_11_io_out_control_0_shift) ^ ((fiEnable && (2898 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_11_io_in_control_0_dataflow_b <=( _mesh_18_11_io_out_control_0_dataflow) ^ ((fiEnable && (2899 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_11_io_in_control_0_propagate_b <=( _mesh_18_11_io_out_control_0_propagate) ^ ((fiEnable && (2900 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_11_io_out_valid_0) begin
			b_372_0 <=( _mesh_19_11_io_out_b_0) ^ ((fiEnable && (2901 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1396_0 <=( _mesh_19_11_io_out_c_0) ^ ((fiEnable && (2902 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_11_io_in_control_0_shift_b <=( _mesh_19_11_io_out_control_0_shift) ^ ((fiEnable && (2903 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_11_io_in_control_0_dataflow_b <=( _mesh_19_11_io_out_control_0_dataflow) ^ ((fiEnable && (2904 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_11_io_in_control_0_propagate_b <=( _mesh_19_11_io_out_control_0_propagate) ^ ((fiEnable && (2905 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_11_io_out_valid_0) begin
			b_373_0 <=( _mesh_20_11_io_out_b_0) ^ ((fiEnable && (2906 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1397_0 <=( _mesh_20_11_io_out_c_0) ^ ((fiEnable && (2907 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_11_io_in_control_0_shift_b <=( _mesh_20_11_io_out_control_0_shift) ^ ((fiEnable && (2908 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_11_io_in_control_0_dataflow_b <=( _mesh_20_11_io_out_control_0_dataflow) ^ ((fiEnable && (2909 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_11_io_in_control_0_propagate_b <=( _mesh_20_11_io_out_control_0_propagate) ^ ((fiEnable && (2910 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_11_io_out_valid_0) begin
			b_374_0 <=( _mesh_21_11_io_out_b_0) ^ ((fiEnable && (2911 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1398_0 <=( _mesh_21_11_io_out_c_0) ^ ((fiEnable && (2912 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_11_io_in_control_0_shift_b <=( _mesh_21_11_io_out_control_0_shift) ^ ((fiEnable && (2913 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_11_io_in_control_0_dataflow_b <=( _mesh_21_11_io_out_control_0_dataflow) ^ ((fiEnable && (2914 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_11_io_in_control_0_propagate_b <=( _mesh_21_11_io_out_control_0_propagate) ^ ((fiEnable && (2915 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_11_io_out_valid_0) begin
			b_375_0 <=( _mesh_22_11_io_out_b_0) ^ ((fiEnable && (2916 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1399_0 <=( _mesh_22_11_io_out_c_0) ^ ((fiEnable && (2917 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_11_io_in_control_0_shift_b <=( _mesh_22_11_io_out_control_0_shift) ^ ((fiEnable && (2918 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_11_io_in_control_0_dataflow_b <=( _mesh_22_11_io_out_control_0_dataflow) ^ ((fiEnable && (2919 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_11_io_in_control_0_propagate_b <=( _mesh_22_11_io_out_control_0_propagate) ^ ((fiEnable && (2920 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_11_io_out_valid_0) begin
			b_376_0 <=( _mesh_23_11_io_out_b_0) ^ ((fiEnable && (2921 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1400_0 <=( _mesh_23_11_io_out_c_0) ^ ((fiEnable && (2922 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_11_io_in_control_0_shift_b <=( _mesh_23_11_io_out_control_0_shift) ^ ((fiEnable && (2923 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_11_io_in_control_0_dataflow_b <=( _mesh_23_11_io_out_control_0_dataflow) ^ ((fiEnable && (2924 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_11_io_in_control_0_propagate_b <=( _mesh_23_11_io_out_control_0_propagate) ^ ((fiEnable && (2925 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_11_io_out_valid_0) begin
			b_377_0 <=( _mesh_24_11_io_out_b_0) ^ ((fiEnable && (2926 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1401_0 <=( _mesh_24_11_io_out_c_0) ^ ((fiEnable && (2927 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_11_io_in_control_0_shift_b <=( _mesh_24_11_io_out_control_0_shift) ^ ((fiEnable && (2928 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_11_io_in_control_0_dataflow_b <=( _mesh_24_11_io_out_control_0_dataflow) ^ ((fiEnable && (2929 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_11_io_in_control_0_propagate_b <=( _mesh_24_11_io_out_control_0_propagate) ^ ((fiEnable && (2930 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_11_io_out_valid_0) begin
			b_378_0 <=( _mesh_25_11_io_out_b_0) ^ ((fiEnable && (2931 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1402_0 <=( _mesh_25_11_io_out_c_0) ^ ((fiEnable && (2932 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_11_io_in_control_0_shift_b <=( _mesh_25_11_io_out_control_0_shift) ^ ((fiEnable && (2933 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_11_io_in_control_0_dataflow_b <=( _mesh_25_11_io_out_control_0_dataflow) ^ ((fiEnable && (2934 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_11_io_in_control_0_propagate_b <=( _mesh_25_11_io_out_control_0_propagate) ^ ((fiEnable && (2935 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_11_io_out_valid_0) begin
			b_379_0 <=( _mesh_26_11_io_out_b_0) ^ ((fiEnable && (2936 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1403_0 <=( _mesh_26_11_io_out_c_0) ^ ((fiEnable && (2937 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_11_io_in_control_0_shift_b <=( _mesh_26_11_io_out_control_0_shift) ^ ((fiEnable && (2938 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_11_io_in_control_0_dataflow_b <=( _mesh_26_11_io_out_control_0_dataflow) ^ ((fiEnable && (2939 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_11_io_in_control_0_propagate_b <=( _mesh_26_11_io_out_control_0_propagate) ^ ((fiEnable && (2940 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_11_io_out_valid_0) begin
			b_380_0 <=( _mesh_27_11_io_out_b_0) ^ ((fiEnable && (2941 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1404_0 <=( _mesh_27_11_io_out_c_0) ^ ((fiEnable && (2942 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_11_io_in_control_0_shift_b <=( _mesh_27_11_io_out_control_0_shift) ^ ((fiEnable && (2943 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_11_io_in_control_0_dataflow_b <=( _mesh_27_11_io_out_control_0_dataflow) ^ ((fiEnable && (2944 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_11_io_in_control_0_propagate_b <=( _mesh_27_11_io_out_control_0_propagate) ^ ((fiEnable && (2945 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_11_io_out_valid_0) begin
			b_381_0 <=( _mesh_28_11_io_out_b_0) ^ ((fiEnable && (2946 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1405_0 <=( _mesh_28_11_io_out_c_0) ^ ((fiEnable && (2947 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_11_io_in_control_0_shift_b <=( _mesh_28_11_io_out_control_0_shift) ^ ((fiEnable && (2948 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_11_io_in_control_0_dataflow_b <=( _mesh_28_11_io_out_control_0_dataflow) ^ ((fiEnable && (2949 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_11_io_in_control_0_propagate_b <=( _mesh_28_11_io_out_control_0_propagate) ^ ((fiEnable && (2950 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_11_io_out_valid_0) begin
			b_382_0 <=( _mesh_29_11_io_out_b_0) ^ ((fiEnable && (2951 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1406_0 <=( _mesh_29_11_io_out_c_0) ^ ((fiEnable && (2952 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_11_io_in_control_0_shift_b <=( _mesh_29_11_io_out_control_0_shift) ^ ((fiEnable && (2953 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_11_io_in_control_0_dataflow_b <=( _mesh_29_11_io_out_control_0_dataflow) ^ ((fiEnable && (2954 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_11_io_in_control_0_propagate_b <=( _mesh_29_11_io_out_control_0_propagate) ^ ((fiEnable && (2955 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_11_io_out_valid_0) begin
			b_383_0 <=( _mesh_30_11_io_out_b_0) ^ ((fiEnable && (2956 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1407_0 <=( _mesh_30_11_io_out_c_0) ^ ((fiEnable && (2957 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_11_io_in_control_0_shift_b <=( _mesh_30_11_io_out_control_0_shift) ^ ((fiEnable && (2958 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_11_io_in_control_0_dataflow_b <=( _mesh_30_11_io_out_control_0_dataflow) ^ ((fiEnable && (2959 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_11_io_in_control_0_propagate_b <=( _mesh_30_11_io_out_control_0_propagate) ^ ((fiEnable && (2960 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_12_0) begin
			b_384_0 <=( io_in_b_12_0) ^ ((fiEnable && (2961 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1408_0 <=( io_in_d_12_0) ^ ((fiEnable && (2962 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_12_io_in_control_0_shift_b <=( io_in_control_12_0_shift) ^ ((fiEnable && (2963 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_12_io_in_control_0_dataflow_b <=( io_in_control_12_0_dataflow) ^ ((fiEnable && (2964 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_12_io_in_control_0_propagate_b <=( io_in_control_12_0_propagate) ^ ((fiEnable && (2965 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_12_io_out_valid_0) begin
			b_385_0 <=( _mesh_0_12_io_out_b_0) ^ ((fiEnable && (2966 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1409_0 <=( _mesh_0_12_io_out_c_0) ^ ((fiEnable && (2967 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_12_io_in_control_0_shift_b <=( _mesh_0_12_io_out_control_0_shift) ^ ((fiEnable && (2968 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_12_io_in_control_0_dataflow_b <=( _mesh_0_12_io_out_control_0_dataflow) ^ ((fiEnable && (2969 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_12_io_in_control_0_propagate_b <=( _mesh_0_12_io_out_control_0_propagate) ^ ((fiEnable && (2970 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_12_io_out_valid_0) begin
			b_386_0 <=( _mesh_1_12_io_out_b_0) ^ ((fiEnable && (2971 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1410_0 <=( _mesh_1_12_io_out_c_0) ^ ((fiEnable && (2972 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_12_io_in_control_0_shift_b <=( _mesh_1_12_io_out_control_0_shift) ^ ((fiEnable && (2973 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_12_io_in_control_0_dataflow_b <=( _mesh_1_12_io_out_control_0_dataflow) ^ ((fiEnable && (2974 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_12_io_in_control_0_propagate_b <=( _mesh_1_12_io_out_control_0_propagate) ^ ((fiEnable && (2975 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_12_io_out_valid_0) begin
			b_387_0 <=( _mesh_2_12_io_out_b_0) ^ ((fiEnable && (2976 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1411_0 <=( _mesh_2_12_io_out_c_0) ^ ((fiEnable && (2977 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_12_io_in_control_0_shift_b <=( _mesh_2_12_io_out_control_0_shift) ^ ((fiEnable && (2978 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_12_io_in_control_0_dataflow_b <=( _mesh_2_12_io_out_control_0_dataflow) ^ ((fiEnable && (2979 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_12_io_in_control_0_propagate_b <=( _mesh_2_12_io_out_control_0_propagate) ^ ((fiEnable && (2980 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_12_io_out_valid_0) begin
			b_388_0 <=( _mesh_3_12_io_out_b_0) ^ ((fiEnable && (2981 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1412_0 <=( _mesh_3_12_io_out_c_0) ^ ((fiEnable && (2982 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_12_io_in_control_0_shift_b <=( _mesh_3_12_io_out_control_0_shift) ^ ((fiEnable && (2983 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_12_io_in_control_0_dataflow_b <=( _mesh_3_12_io_out_control_0_dataflow) ^ ((fiEnable && (2984 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_12_io_in_control_0_propagate_b <=( _mesh_3_12_io_out_control_0_propagate) ^ ((fiEnable && (2985 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_12_io_out_valid_0) begin
			b_389_0 <=( _mesh_4_12_io_out_b_0) ^ ((fiEnable && (2986 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1413_0 <=( _mesh_4_12_io_out_c_0) ^ ((fiEnable && (2987 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_12_io_in_control_0_shift_b <=( _mesh_4_12_io_out_control_0_shift) ^ ((fiEnable && (2988 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_12_io_in_control_0_dataflow_b <=( _mesh_4_12_io_out_control_0_dataflow) ^ ((fiEnable && (2989 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_12_io_in_control_0_propagate_b <=( _mesh_4_12_io_out_control_0_propagate) ^ ((fiEnable && (2990 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_12_io_out_valid_0) begin
			b_390_0 <=( _mesh_5_12_io_out_b_0) ^ ((fiEnable && (2991 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1414_0 <=( _mesh_5_12_io_out_c_0) ^ ((fiEnable && (2992 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_12_io_in_control_0_shift_b <=( _mesh_5_12_io_out_control_0_shift) ^ ((fiEnable && (2993 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_12_io_in_control_0_dataflow_b <=( _mesh_5_12_io_out_control_0_dataflow) ^ ((fiEnable && (2994 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_12_io_in_control_0_propagate_b <=( _mesh_5_12_io_out_control_0_propagate) ^ ((fiEnable && (2995 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_12_io_out_valid_0) begin
			b_391_0 <=( _mesh_6_12_io_out_b_0) ^ ((fiEnable && (2996 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1415_0 <=( _mesh_6_12_io_out_c_0) ^ ((fiEnable && (2997 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_12_io_in_control_0_shift_b <=( _mesh_6_12_io_out_control_0_shift) ^ ((fiEnable && (2998 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_12_io_in_control_0_dataflow_b <=( _mesh_6_12_io_out_control_0_dataflow) ^ ((fiEnable && (2999 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_12_io_in_control_0_propagate_b <=( _mesh_6_12_io_out_control_0_propagate) ^ ((fiEnable && (3000 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_12_io_out_valid_0) begin
			b_392_0 <=( _mesh_7_12_io_out_b_0) ^ ((fiEnable && (3001 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1416_0 <=( _mesh_7_12_io_out_c_0) ^ ((fiEnable && (3002 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_12_io_in_control_0_shift_b <=( _mesh_7_12_io_out_control_0_shift) ^ ((fiEnable && (3003 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_12_io_in_control_0_dataflow_b <=( _mesh_7_12_io_out_control_0_dataflow) ^ ((fiEnable && (3004 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_12_io_in_control_0_propagate_b <=( _mesh_7_12_io_out_control_0_propagate) ^ ((fiEnable && (3005 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_12_io_out_valid_0) begin
			b_393_0 <=( _mesh_8_12_io_out_b_0) ^ ((fiEnable && (3006 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1417_0 <=( _mesh_8_12_io_out_c_0) ^ ((fiEnable && (3007 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_12_io_in_control_0_shift_b <=( _mesh_8_12_io_out_control_0_shift) ^ ((fiEnable && (3008 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_12_io_in_control_0_dataflow_b <=( _mesh_8_12_io_out_control_0_dataflow) ^ ((fiEnable && (3009 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_12_io_in_control_0_propagate_b <=( _mesh_8_12_io_out_control_0_propagate) ^ ((fiEnable && (3010 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_12_io_out_valid_0) begin
			b_394_0 <=( _mesh_9_12_io_out_b_0) ^ ((fiEnable && (3011 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1418_0 <=( _mesh_9_12_io_out_c_0) ^ ((fiEnable && (3012 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_12_io_in_control_0_shift_b <=( _mesh_9_12_io_out_control_0_shift) ^ ((fiEnable && (3013 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_12_io_in_control_0_dataflow_b <=( _mesh_9_12_io_out_control_0_dataflow) ^ ((fiEnable && (3014 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_12_io_in_control_0_propagate_b <=( _mesh_9_12_io_out_control_0_propagate) ^ ((fiEnable && (3015 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_12_io_out_valid_0) begin
			b_395_0 <=( _mesh_10_12_io_out_b_0) ^ ((fiEnable && (3016 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1419_0 <=( _mesh_10_12_io_out_c_0) ^ ((fiEnable && (3017 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_12_io_in_control_0_shift_b <=( _mesh_10_12_io_out_control_0_shift) ^ ((fiEnable && (3018 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_12_io_in_control_0_dataflow_b <=( _mesh_10_12_io_out_control_0_dataflow) ^ ((fiEnable && (3019 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_12_io_in_control_0_propagate_b <=( _mesh_10_12_io_out_control_0_propagate) ^ ((fiEnable && (3020 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_12_io_out_valid_0) begin
			b_396_0 <=( _mesh_11_12_io_out_b_0) ^ ((fiEnable && (3021 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1420_0 <=( _mesh_11_12_io_out_c_0) ^ ((fiEnable && (3022 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_12_io_in_control_0_shift_b <=( _mesh_11_12_io_out_control_0_shift) ^ ((fiEnable && (3023 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_12_io_in_control_0_dataflow_b <=( _mesh_11_12_io_out_control_0_dataflow) ^ ((fiEnable && (3024 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_12_io_in_control_0_propagate_b <=( _mesh_11_12_io_out_control_0_propagate) ^ ((fiEnable && (3025 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_12_io_out_valid_0) begin
			b_397_0 <=( _mesh_12_12_io_out_b_0) ^ ((fiEnable && (3026 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1421_0 <=( _mesh_12_12_io_out_c_0) ^ ((fiEnable && (3027 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_12_io_in_control_0_shift_b <=( _mesh_12_12_io_out_control_0_shift) ^ ((fiEnable && (3028 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_12_io_in_control_0_dataflow_b <=( _mesh_12_12_io_out_control_0_dataflow) ^ ((fiEnable && (3029 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_12_io_in_control_0_propagate_b <=( _mesh_12_12_io_out_control_0_propagate) ^ ((fiEnable && (3030 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_12_io_out_valid_0) begin
			b_398_0 <=( _mesh_13_12_io_out_b_0) ^ ((fiEnable && (3031 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1422_0 <=( _mesh_13_12_io_out_c_0) ^ ((fiEnable && (3032 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_12_io_in_control_0_shift_b <=( _mesh_13_12_io_out_control_0_shift) ^ ((fiEnable && (3033 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_12_io_in_control_0_dataflow_b <=( _mesh_13_12_io_out_control_0_dataflow) ^ ((fiEnable && (3034 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_12_io_in_control_0_propagate_b <=( _mesh_13_12_io_out_control_0_propagate) ^ ((fiEnable && (3035 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_12_io_out_valid_0) begin
			b_399_0 <=( _mesh_14_12_io_out_b_0) ^ ((fiEnable && (3036 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1423_0 <=( _mesh_14_12_io_out_c_0) ^ ((fiEnable && (3037 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_12_io_in_control_0_shift_b <=( _mesh_14_12_io_out_control_0_shift) ^ ((fiEnable && (3038 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_12_io_in_control_0_dataflow_b <=( _mesh_14_12_io_out_control_0_dataflow) ^ ((fiEnable && (3039 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_12_io_in_control_0_propagate_b <=( _mesh_14_12_io_out_control_0_propagate) ^ ((fiEnable && (3040 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_12_io_out_valid_0) begin
			b_400_0 <=( _mesh_15_12_io_out_b_0) ^ ((fiEnable && (3041 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1424_0 <=( _mesh_15_12_io_out_c_0) ^ ((fiEnable && (3042 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_12_io_in_control_0_shift_b <=( _mesh_15_12_io_out_control_0_shift) ^ ((fiEnable && (3043 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_12_io_in_control_0_dataflow_b <=( _mesh_15_12_io_out_control_0_dataflow) ^ ((fiEnable && (3044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_12_io_in_control_0_propagate_b <=( _mesh_15_12_io_out_control_0_propagate) ^ ((fiEnable && (3045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_12_io_out_valid_0) begin
			b_401_0 <=( _mesh_16_12_io_out_b_0) ^ ((fiEnable && (3046 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1425_0 <=( _mesh_16_12_io_out_c_0) ^ ((fiEnable && (3047 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_12_io_in_control_0_shift_b <=( _mesh_16_12_io_out_control_0_shift) ^ ((fiEnable && (3048 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_12_io_in_control_0_dataflow_b <=( _mesh_16_12_io_out_control_0_dataflow) ^ ((fiEnable && (3049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_12_io_in_control_0_propagate_b <=( _mesh_16_12_io_out_control_0_propagate) ^ ((fiEnable && (3050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_12_io_out_valid_0) begin
			b_402_0 <=( _mesh_17_12_io_out_b_0) ^ ((fiEnable && (3051 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1426_0 <=( _mesh_17_12_io_out_c_0) ^ ((fiEnable && (3052 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_12_io_in_control_0_shift_b <=( _mesh_17_12_io_out_control_0_shift) ^ ((fiEnable && (3053 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_12_io_in_control_0_dataflow_b <=( _mesh_17_12_io_out_control_0_dataflow) ^ ((fiEnable && (3054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_12_io_in_control_0_propagate_b <=( _mesh_17_12_io_out_control_0_propagate) ^ ((fiEnable && (3055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_12_io_out_valid_0) begin
			b_403_0 <=( _mesh_18_12_io_out_b_0) ^ ((fiEnable && (3056 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1427_0 <=( _mesh_18_12_io_out_c_0) ^ ((fiEnable && (3057 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_12_io_in_control_0_shift_b <=( _mesh_18_12_io_out_control_0_shift) ^ ((fiEnable && (3058 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_12_io_in_control_0_dataflow_b <=( _mesh_18_12_io_out_control_0_dataflow) ^ ((fiEnable && (3059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_12_io_in_control_0_propagate_b <=( _mesh_18_12_io_out_control_0_propagate) ^ ((fiEnable && (3060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_12_io_out_valid_0) begin
			b_404_0 <=( _mesh_19_12_io_out_b_0) ^ ((fiEnable && (3061 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1428_0 <=( _mesh_19_12_io_out_c_0) ^ ((fiEnable && (3062 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_12_io_in_control_0_shift_b <=( _mesh_19_12_io_out_control_0_shift) ^ ((fiEnable && (3063 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_12_io_in_control_0_dataflow_b <=( _mesh_19_12_io_out_control_0_dataflow) ^ ((fiEnable && (3064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_12_io_in_control_0_propagate_b <=( _mesh_19_12_io_out_control_0_propagate) ^ ((fiEnable && (3065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_12_io_out_valid_0) begin
			b_405_0 <=( _mesh_20_12_io_out_b_0) ^ ((fiEnable && (3066 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1429_0 <=( _mesh_20_12_io_out_c_0) ^ ((fiEnable && (3067 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_12_io_in_control_0_shift_b <=( _mesh_20_12_io_out_control_0_shift) ^ ((fiEnable && (3068 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_12_io_in_control_0_dataflow_b <=( _mesh_20_12_io_out_control_0_dataflow) ^ ((fiEnable && (3069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_12_io_in_control_0_propagate_b <=( _mesh_20_12_io_out_control_0_propagate) ^ ((fiEnable && (3070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_12_io_out_valid_0) begin
			b_406_0 <=( _mesh_21_12_io_out_b_0) ^ ((fiEnable && (3071 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1430_0 <=( _mesh_21_12_io_out_c_0) ^ ((fiEnable && (3072 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_12_io_in_control_0_shift_b <=( _mesh_21_12_io_out_control_0_shift) ^ ((fiEnable && (3073 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_12_io_in_control_0_dataflow_b <=( _mesh_21_12_io_out_control_0_dataflow) ^ ((fiEnable && (3074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_12_io_in_control_0_propagate_b <=( _mesh_21_12_io_out_control_0_propagate) ^ ((fiEnable && (3075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_12_io_out_valid_0) begin
			b_407_0 <=( _mesh_22_12_io_out_b_0) ^ ((fiEnable && (3076 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1431_0 <=( _mesh_22_12_io_out_c_0) ^ ((fiEnable && (3077 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_12_io_in_control_0_shift_b <=( _mesh_22_12_io_out_control_0_shift) ^ ((fiEnable && (3078 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_12_io_in_control_0_dataflow_b <=( _mesh_22_12_io_out_control_0_dataflow) ^ ((fiEnable && (3079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_12_io_in_control_0_propagate_b <=( _mesh_22_12_io_out_control_0_propagate) ^ ((fiEnable && (3080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_12_io_out_valid_0) begin
			b_408_0 <=( _mesh_23_12_io_out_b_0) ^ ((fiEnable && (3081 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1432_0 <=( _mesh_23_12_io_out_c_0) ^ ((fiEnable && (3082 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_12_io_in_control_0_shift_b <=( _mesh_23_12_io_out_control_0_shift) ^ ((fiEnable && (3083 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_12_io_in_control_0_dataflow_b <=( _mesh_23_12_io_out_control_0_dataflow) ^ ((fiEnable && (3084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_12_io_in_control_0_propagate_b <=( _mesh_23_12_io_out_control_0_propagate) ^ ((fiEnable && (3085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_12_io_out_valid_0) begin
			b_409_0 <=( _mesh_24_12_io_out_b_0) ^ ((fiEnable && (3086 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1433_0 <=( _mesh_24_12_io_out_c_0) ^ ((fiEnable && (3087 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_12_io_in_control_0_shift_b <=( _mesh_24_12_io_out_control_0_shift) ^ ((fiEnable && (3088 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_12_io_in_control_0_dataflow_b <=( _mesh_24_12_io_out_control_0_dataflow) ^ ((fiEnable && (3089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_12_io_in_control_0_propagate_b <=( _mesh_24_12_io_out_control_0_propagate) ^ ((fiEnable && (3090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_12_io_out_valid_0) begin
			b_410_0 <=( _mesh_25_12_io_out_b_0) ^ ((fiEnable && (3091 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1434_0 <=( _mesh_25_12_io_out_c_0) ^ ((fiEnable && (3092 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_12_io_in_control_0_shift_b <=( _mesh_25_12_io_out_control_0_shift) ^ ((fiEnable && (3093 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_12_io_in_control_0_dataflow_b <=( _mesh_25_12_io_out_control_0_dataflow) ^ ((fiEnable && (3094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_12_io_in_control_0_propagate_b <=( _mesh_25_12_io_out_control_0_propagate) ^ ((fiEnable && (3095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_12_io_out_valid_0) begin
			b_411_0 <=( _mesh_26_12_io_out_b_0) ^ ((fiEnable && (3096 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1435_0 <=( _mesh_26_12_io_out_c_0) ^ ((fiEnable && (3097 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_12_io_in_control_0_shift_b <=( _mesh_26_12_io_out_control_0_shift) ^ ((fiEnable && (3098 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_12_io_in_control_0_dataflow_b <=( _mesh_26_12_io_out_control_0_dataflow) ^ ((fiEnable && (3099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_12_io_in_control_0_propagate_b <=( _mesh_26_12_io_out_control_0_propagate) ^ ((fiEnable && (3100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_12_io_out_valid_0) begin
			b_412_0 <=( _mesh_27_12_io_out_b_0) ^ ((fiEnable && (3101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1436_0 <=( _mesh_27_12_io_out_c_0) ^ ((fiEnable && (3102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_12_io_in_control_0_shift_b <=( _mesh_27_12_io_out_control_0_shift) ^ ((fiEnable && (3103 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_12_io_in_control_0_dataflow_b <=( _mesh_27_12_io_out_control_0_dataflow) ^ ((fiEnable && (3104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_12_io_in_control_0_propagate_b <=( _mesh_27_12_io_out_control_0_propagate) ^ ((fiEnable && (3105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_12_io_out_valid_0) begin
			b_413_0 <=( _mesh_28_12_io_out_b_0) ^ ((fiEnable && (3106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1437_0 <=( _mesh_28_12_io_out_c_0) ^ ((fiEnable && (3107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_12_io_in_control_0_shift_b <=( _mesh_28_12_io_out_control_0_shift) ^ ((fiEnable && (3108 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_12_io_in_control_0_dataflow_b <=( _mesh_28_12_io_out_control_0_dataflow) ^ ((fiEnable && (3109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_12_io_in_control_0_propagate_b <=( _mesh_28_12_io_out_control_0_propagate) ^ ((fiEnable && (3110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_12_io_out_valid_0) begin
			b_414_0 <=( _mesh_29_12_io_out_b_0) ^ ((fiEnable && (3111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1438_0 <=( _mesh_29_12_io_out_c_0) ^ ((fiEnable && (3112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_12_io_in_control_0_shift_b <=( _mesh_29_12_io_out_control_0_shift) ^ ((fiEnable && (3113 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_12_io_in_control_0_dataflow_b <=( _mesh_29_12_io_out_control_0_dataflow) ^ ((fiEnable && (3114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_12_io_in_control_0_propagate_b <=( _mesh_29_12_io_out_control_0_propagate) ^ ((fiEnable && (3115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_12_io_out_valid_0) begin
			b_415_0 <=( _mesh_30_12_io_out_b_0) ^ ((fiEnable && (3116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1439_0 <=( _mesh_30_12_io_out_c_0) ^ ((fiEnable && (3117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_12_io_in_control_0_shift_b <=( _mesh_30_12_io_out_control_0_shift) ^ ((fiEnable && (3118 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_12_io_in_control_0_dataflow_b <=( _mesh_30_12_io_out_control_0_dataflow) ^ ((fiEnable && (3119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_12_io_in_control_0_propagate_b <=( _mesh_30_12_io_out_control_0_propagate) ^ ((fiEnable && (3120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_13_0) begin
			b_416_0 <=( io_in_b_13_0) ^ ((fiEnable && (3121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1440_0 <=( io_in_d_13_0) ^ ((fiEnable && (3122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_13_io_in_control_0_shift_b <=( io_in_control_13_0_shift) ^ ((fiEnable && (3123 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_13_io_in_control_0_dataflow_b <=( io_in_control_13_0_dataflow) ^ ((fiEnable && (3124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_13_io_in_control_0_propagate_b <=( io_in_control_13_0_propagate) ^ ((fiEnable && (3125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_13_io_out_valid_0) begin
			b_417_0 <=( _mesh_0_13_io_out_b_0) ^ ((fiEnable && (3126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1441_0 <=( _mesh_0_13_io_out_c_0) ^ ((fiEnable && (3127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_13_io_in_control_0_shift_b <=( _mesh_0_13_io_out_control_0_shift) ^ ((fiEnable && (3128 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_13_io_in_control_0_dataflow_b <=( _mesh_0_13_io_out_control_0_dataflow) ^ ((fiEnable && (3129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_13_io_in_control_0_propagate_b <=( _mesh_0_13_io_out_control_0_propagate) ^ ((fiEnable && (3130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_13_io_out_valid_0) begin
			b_418_0 <=( _mesh_1_13_io_out_b_0) ^ ((fiEnable && (3131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1442_0 <=( _mesh_1_13_io_out_c_0) ^ ((fiEnable && (3132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_13_io_in_control_0_shift_b <=( _mesh_1_13_io_out_control_0_shift) ^ ((fiEnable && (3133 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_13_io_in_control_0_dataflow_b <=( _mesh_1_13_io_out_control_0_dataflow) ^ ((fiEnable && (3134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_13_io_in_control_0_propagate_b <=( _mesh_1_13_io_out_control_0_propagate) ^ ((fiEnable && (3135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_13_io_out_valid_0) begin
			b_419_0 <=( _mesh_2_13_io_out_b_0) ^ ((fiEnable && (3136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1443_0 <=( _mesh_2_13_io_out_c_0) ^ ((fiEnable && (3137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_13_io_in_control_0_shift_b <=( _mesh_2_13_io_out_control_0_shift) ^ ((fiEnable && (3138 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_13_io_in_control_0_dataflow_b <=( _mesh_2_13_io_out_control_0_dataflow) ^ ((fiEnable && (3139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_13_io_in_control_0_propagate_b <=( _mesh_2_13_io_out_control_0_propagate) ^ ((fiEnable && (3140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_13_io_out_valid_0) begin
			b_420_0 <=( _mesh_3_13_io_out_b_0) ^ ((fiEnable && (3141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1444_0 <=( _mesh_3_13_io_out_c_0) ^ ((fiEnable && (3142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_13_io_in_control_0_shift_b <=( _mesh_3_13_io_out_control_0_shift) ^ ((fiEnable && (3143 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_13_io_in_control_0_dataflow_b <=( _mesh_3_13_io_out_control_0_dataflow) ^ ((fiEnable && (3144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_13_io_in_control_0_propagate_b <=( _mesh_3_13_io_out_control_0_propagate) ^ ((fiEnable && (3145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_13_io_out_valid_0) begin
			b_421_0 <=( _mesh_4_13_io_out_b_0) ^ ((fiEnable && (3146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1445_0 <=( _mesh_4_13_io_out_c_0) ^ ((fiEnable && (3147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_13_io_in_control_0_shift_b <=( _mesh_4_13_io_out_control_0_shift) ^ ((fiEnable && (3148 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_13_io_in_control_0_dataflow_b <=( _mesh_4_13_io_out_control_0_dataflow) ^ ((fiEnable && (3149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_13_io_in_control_0_propagate_b <=( _mesh_4_13_io_out_control_0_propagate) ^ ((fiEnable && (3150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_13_io_out_valid_0) begin
			b_422_0 <=( _mesh_5_13_io_out_b_0) ^ ((fiEnable && (3151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1446_0 <=( _mesh_5_13_io_out_c_0) ^ ((fiEnable && (3152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_13_io_in_control_0_shift_b <=( _mesh_5_13_io_out_control_0_shift) ^ ((fiEnable && (3153 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_13_io_in_control_0_dataflow_b <=( _mesh_5_13_io_out_control_0_dataflow) ^ ((fiEnable && (3154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_13_io_in_control_0_propagate_b <=( _mesh_5_13_io_out_control_0_propagate) ^ ((fiEnable && (3155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_13_io_out_valid_0) begin
			b_423_0 <=( _mesh_6_13_io_out_b_0) ^ ((fiEnable && (3156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1447_0 <=( _mesh_6_13_io_out_c_0) ^ ((fiEnable && (3157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_13_io_in_control_0_shift_b <=( _mesh_6_13_io_out_control_0_shift) ^ ((fiEnable && (3158 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_13_io_in_control_0_dataflow_b <=( _mesh_6_13_io_out_control_0_dataflow) ^ ((fiEnable && (3159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_13_io_in_control_0_propagate_b <=( _mesh_6_13_io_out_control_0_propagate) ^ ((fiEnable && (3160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_13_io_out_valid_0) begin
			b_424_0 <=( _mesh_7_13_io_out_b_0) ^ ((fiEnable && (3161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1448_0 <=( _mesh_7_13_io_out_c_0) ^ ((fiEnable && (3162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_13_io_in_control_0_shift_b <=( _mesh_7_13_io_out_control_0_shift) ^ ((fiEnable && (3163 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_13_io_in_control_0_dataflow_b <=( _mesh_7_13_io_out_control_0_dataflow) ^ ((fiEnable && (3164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_13_io_in_control_0_propagate_b <=( _mesh_7_13_io_out_control_0_propagate) ^ ((fiEnable && (3165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_13_io_out_valid_0) begin
			b_425_0 <=( _mesh_8_13_io_out_b_0) ^ ((fiEnable && (3166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1449_0 <=( _mesh_8_13_io_out_c_0) ^ ((fiEnable && (3167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_13_io_in_control_0_shift_b <=( _mesh_8_13_io_out_control_0_shift) ^ ((fiEnable && (3168 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_13_io_in_control_0_dataflow_b <=( _mesh_8_13_io_out_control_0_dataflow) ^ ((fiEnable && (3169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_13_io_in_control_0_propagate_b <=( _mesh_8_13_io_out_control_0_propagate) ^ ((fiEnable && (3170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_13_io_out_valid_0) begin
			b_426_0 <=( _mesh_9_13_io_out_b_0) ^ ((fiEnable && (3171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1450_0 <=( _mesh_9_13_io_out_c_0) ^ ((fiEnable && (3172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_13_io_in_control_0_shift_b <=( _mesh_9_13_io_out_control_0_shift) ^ ((fiEnable && (3173 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_13_io_in_control_0_dataflow_b <=( _mesh_9_13_io_out_control_0_dataflow) ^ ((fiEnable && (3174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_13_io_in_control_0_propagate_b <=( _mesh_9_13_io_out_control_0_propagate) ^ ((fiEnable && (3175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_13_io_out_valid_0) begin
			b_427_0 <=( _mesh_10_13_io_out_b_0) ^ ((fiEnable && (3176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1451_0 <=( _mesh_10_13_io_out_c_0) ^ ((fiEnable && (3177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_13_io_in_control_0_shift_b <=( _mesh_10_13_io_out_control_0_shift) ^ ((fiEnable && (3178 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_13_io_in_control_0_dataflow_b <=( _mesh_10_13_io_out_control_0_dataflow) ^ ((fiEnable && (3179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_13_io_in_control_0_propagate_b <=( _mesh_10_13_io_out_control_0_propagate) ^ ((fiEnable && (3180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_13_io_out_valid_0) begin
			b_428_0 <=( _mesh_11_13_io_out_b_0) ^ ((fiEnable && (3181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1452_0 <=( _mesh_11_13_io_out_c_0) ^ ((fiEnable && (3182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_13_io_in_control_0_shift_b <=( _mesh_11_13_io_out_control_0_shift) ^ ((fiEnable && (3183 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_13_io_in_control_0_dataflow_b <=( _mesh_11_13_io_out_control_0_dataflow) ^ ((fiEnable && (3184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_13_io_in_control_0_propagate_b <=( _mesh_11_13_io_out_control_0_propagate) ^ ((fiEnable && (3185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_13_io_out_valid_0) begin
			b_429_0 <=( _mesh_12_13_io_out_b_0) ^ ((fiEnable && (3186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1453_0 <=( _mesh_12_13_io_out_c_0) ^ ((fiEnable && (3187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_13_io_in_control_0_shift_b <=( _mesh_12_13_io_out_control_0_shift) ^ ((fiEnable && (3188 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_13_io_in_control_0_dataflow_b <=( _mesh_12_13_io_out_control_0_dataflow) ^ ((fiEnable && (3189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_13_io_in_control_0_propagate_b <=( _mesh_12_13_io_out_control_0_propagate) ^ ((fiEnable && (3190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_13_io_out_valid_0) begin
			b_430_0 <=( _mesh_13_13_io_out_b_0) ^ ((fiEnable && (3191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1454_0 <=( _mesh_13_13_io_out_c_0) ^ ((fiEnable && (3192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_13_io_in_control_0_shift_b <=( _mesh_13_13_io_out_control_0_shift) ^ ((fiEnable && (3193 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_13_io_in_control_0_dataflow_b <=( _mesh_13_13_io_out_control_0_dataflow) ^ ((fiEnable && (3194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_13_io_in_control_0_propagate_b <=( _mesh_13_13_io_out_control_0_propagate) ^ ((fiEnable && (3195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_13_io_out_valid_0) begin
			b_431_0 <=( _mesh_14_13_io_out_b_0) ^ ((fiEnable && (3196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1455_0 <=( _mesh_14_13_io_out_c_0) ^ ((fiEnable && (3197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_13_io_in_control_0_shift_b <=( _mesh_14_13_io_out_control_0_shift) ^ ((fiEnable && (3198 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_13_io_in_control_0_dataflow_b <=( _mesh_14_13_io_out_control_0_dataflow) ^ ((fiEnable && (3199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_13_io_in_control_0_propagate_b <=( _mesh_14_13_io_out_control_0_propagate) ^ ((fiEnable && (3200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_13_io_out_valid_0) begin
			b_432_0 <=( _mesh_15_13_io_out_b_0) ^ ((fiEnable && (3201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1456_0 <=( _mesh_15_13_io_out_c_0) ^ ((fiEnable && (3202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_13_io_in_control_0_shift_b <=( _mesh_15_13_io_out_control_0_shift) ^ ((fiEnable && (3203 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_13_io_in_control_0_dataflow_b <=( _mesh_15_13_io_out_control_0_dataflow) ^ ((fiEnable && (3204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_13_io_in_control_0_propagate_b <=( _mesh_15_13_io_out_control_0_propagate) ^ ((fiEnable && (3205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_13_io_out_valid_0) begin
			b_433_0 <=( _mesh_16_13_io_out_b_0) ^ ((fiEnable && (3206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1457_0 <=( _mesh_16_13_io_out_c_0) ^ ((fiEnable && (3207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_13_io_in_control_0_shift_b <=( _mesh_16_13_io_out_control_0_shift) ^ ((fiEnable && (3208 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_13_io_in_control_0_dataflow_b <=( _mesh_16_13_io_out_control_0_dataflow) ^ ((fiEnable && (3209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_13_io_in_control_0_propagate_b <=( _mesh_16_13_io_out_control_0_propagate) ^ ((fiEnable && (3210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_13_io_out_valid_0) begin
			b_434_0 <=( _mesh_17_13_io_out_b_0) ^ ((fiEnable && (3211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1458_0 <=( _mesh_17_13_io_out_c_0) ^ ((fiEnable && (3212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_13_io_in_control_0_shift_b <=( _mesh_17_13_io_out_control_0_shift) ^ ((fiEnable && (3213 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_13_io_in_control_0_dataflow_b <=( _mesh_17_13_io_out_control_0_dataflow) ^ ((fiEnable && (3214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_13_io_in_control_0_propagate_b <=( _mesh_17_13_io_out_control_0_propagate) ^ ((fiEnable && (3215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_13_io_out_valid_0) begin
			b_435_0 <=( _mesh_18_13_io_out_b_0) ^ ((fiEnable && (3216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1459_0 <=( _mesh_18_13_io_out_c_0) ^ ((fiEnable && (3217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_13_io_in_control_0_shift_b <=( _mesh_18_13_io_out_control_0_shift) ^ ((fiEnable && (3218 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_13_io_in_control_0_dataflow_b <=( _mesh_18_13_io_out_control_0_dataflow) ^ ((fiEnable && (3219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_13_io_in_control_0_propagate_b <=( _mesh_18_13_io_out_control_0_propagate) ^ ((fiEnable && (3220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_13_io_out_valid_0) begin
			b_436_0 <=( _mesh_19_13_io_out_b_0) ^ ((fiEnable && (3221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1460_0 <=( _mesh_19_13_io_out_c_0) ^ ((fiEnable && (3222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_13_io_in_control_0_shift_b <=( _mesh_19_13_io_out_control_0_shift) ^ ((fiEnable && (3223 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_13_io_in_control_0_dataflow_b <=( _mesh_19_13_io_out_control_0_dataflow) ^ ((fiEnable && (3224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_13_io_in_control_0_propagate_b <=( _mesh_19_13_io_out_control_0_propagate) ^ ((fiEnable && (3225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_13_io_out_valid_0) begin
			b_437_0 <=( _mesh_20_13_io_out_b_0) ^ ((fiEnable && (3226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1461_0 <=( _mesh_20_13_io_out_c_0) ^ ((fiEnable && (3227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_13_io_in_control_0_shift_b <=( _mesh_20_13_io_out_control_0_shift) ^ ((fiEnable && (3228 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_13_io_in_control_0_dataflow_b <=( _mesh_20_13_io_out_control_0_dataflow) ^ ((fiEnable && (3229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_13_io_in_control_0_propagate_b <=( _mesh_20_13_io_out_control_0_propagate) ^ ((fiEnable && (3230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_13_io_out_valid_0) begin
			b_438_0 <=( _mesh_21_13_io_out_b_0) ^ ((fiEnable && (3231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1462_0 <=( _mesh_21_13_io_out_c_0) ^ ((fiEnable && (3232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_13_io_in_control_0_shift_b <=( _mesh_21_13_io_out_control_0_shift) ^ ((fiEnable && (3233 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_13_io_in_control_0_dataflow_b <=( _mesh_21_13_io_out_control_0_dataflow) ^ ((fiEnable && (3234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_13_io_in_control_0_propagate_b <=( _mesh_21_13_io_out_control_0_propagate) ^ ((fiEnable && (3235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_13_io_out_valid_0) begin
			b_439_0 <=( _mesh_22_13_io_out_b_0) ^ ((fiEnable && (3236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1463_0 <=( _mesh_22_13_io_out_c_0) ^ ((fiEnable && (3237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_13_io_in_control_0_shift_b <=( _mesh_22_13_io_out_control_0_shift) ^ ((fiEnable && (3238 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_13_io_in_control_0_dataflow_b <=( _mesh_22_13_io_out_control_0_dataflow) ^ ((fiEnable && (3239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_13_io_in_control_0_propagate_b <=( _mesh_22_13_io_out_control_0_propagate) ^ ((fiEnable && (3240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_13_io_out_valid_0) begin
			b_440_0 <=( _mesh_23_13_io_out_b_0) ^ ((fiEnable && (3241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1464_0 <=( _mesh_23_13_io_out_c_0) ^ ((fiEnable && (3242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_13_io_in_control_0_shift_b <=( _mesh_23_13_io_out_control_0_shift) ^ ((fiEnable && (3243 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_13_io_in_control_0_dataflow_b <=( _mesh_23_13_io_out_control_0_dataflow) ^ ((fiEnable && (3244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_13_io_in_control_0_propagate_b <=( _mesh_23_13_io_out_control_0_propagate) ^ ((fiEnable && (3245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_13_io_out_valid_0) begin
			b_441_0 <=( _mesh_24_13_io_out_b_0) ^ ((fiEnable && (3246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1465_0 <=( _mesh_24_13_io_out_c_0) ^ ((fiEnable && (3247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_13_io_in_control_0_shift_b <=( _mesh_24_13_io_out_control_0_shift) ^ ((fiEnable && (3248 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_13_io_in_control_0_dataflow_b <=( _mesh_24_13_io_out_control_0_dataflow) ^ ((fiEnable && (3249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_13_io_in_control_0_propagate_b <=( _mesh_24_13_io_out_control_0_propagate) ^ ((fiEnable && (3250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_13_io_out_valid_0) begin
			b_442_0 <=( _mesh_25_13_io_out_b_0) ^ ((fiEnable && (3251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1466_0 <=( _mesh_25_13_io_out_c_0) ^ ((fiEnable && (3252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_13_io_in_control_0_shift_b <=( _mesh_25_13_io_out_control_0_shift) ^ ((fiEnable && (3253 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_13_io_in_control_0_dataflow_b <=( _mesh_25_13_io_out_control_0_dataflow) ^ ((fiEnable && (3254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_13_io_in_control_0_propagate_b <=( _mesh_25_13_io_out_control_0_propagate) ^ ((fiEnable && (3255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_13_io_out_valid_0) begin
			b_443_0 <=( _mesh_26_13_io_out_b_0) ^ ((fiEnable && (3256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1467_0 <=( _mesh_26_13_io_out_c_0) ^ ((fiEnable && (3257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_13_io_in_control_0_shift_b <=( _mesh_26_13_io_out_control_0_shift) ^ ((fiEnable && (3258 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_13_io_in_control_0_dataflow_b <=( _mesh_26_13_io_out_control_0_dataflow) ^ ((fiEnable && (3259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_13_io_in_control_0_propagate_b <=( _mesh_26_13_io_out_control_0_propagate) ^ ((fiEnable && (3260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_13_io_out_valid_0) begin
			b_444_0 <=( _mesh_27_13_io_out_b_0) ^ ((fiEnable && (3261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1468_0 <=( _mesh_27_13_io_out_c_0) ^ ((fiEnable && (3262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_13_io_in_control_0_shift_b <=( _mesh_27_13_io_out_control_0_shift) ^ ((fiEnable && (3263 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_13_io_in_control_0_dataflow_b <=( _mesh_27_13_io_out_control_0_dataflow) ^ ((fiEnable && (3264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_13_io_in_control_0_propagate_b <=( _mesh_27_13_io_out_control_0_propagate) ^ ((fiEnable && (3265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_13_io_out_valid_0) begin
			b_445_0 <=( _mesh_28_13_io_out_b_0) ^ ((fiEnable && (3266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1469_0 <=( _mesh_28_13_io_out_c_0) ^ ((fiEnable && (3267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_13_io_in_control_0_shift_b <=( _mesh_28_13_io_out_control_0_shift) ^ ((fiEnable && (3268 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_13_io_in_control_0_dataflow_b <=( _mesh_28_13_io_out_control_0_dataflow) ^ ((fiEnable && (3269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_13_io_in_control_0_propagate_b <=( _mesh_28_13_io_out_control_0_propagate) ^ ((fiEnable && (3270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_13_io_out_valid_0) begin
			b_446_0 <=( _mesh_29_13_io_out_b_0) ^ ((fiEnable && (3271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1470_0 <=( _mesh_29_13_io_out_c_0) ^ ((fiEnable && (3272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_13_io_in_control_0_shift_b <=( _mesh_29_13_io_out_control_0_shift) ^ ((fiEnable && (3273 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_13_io_in_control_0_dataflow_b <=( _mesh_29_13_io_out_control_0_dataflow) ^ ((fiEnable && (3274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_13_io_in_control_0_propagate_b <=( _mesh_29_13_io_out_control_0_propagate) ^ ((fiEnable && (3275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_13_io_out_valid_0) begin
			b_447_0 <=( _mesh_30_13_io_out_b_0) ^ ((fiEnable && (3276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1471_0 <=( _mesh_30_13_io_out_c_0) ^ ((fiEnable && (3277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_13_io_in_control_0_shift_b <=( _mesh_30_13_io_out_control_0_shift) ^ ((fiEnable && (3278 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_13_io_in_control_0_dataflow_b <=( _mesh_30_13_io_out_control_0_dataflow) ^ ((fiEnable && (3279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_13_io_in_control_0_propagate_b <=( _mesh_30_13_io_out_control_0_propagate) ^ ((fiEnable && (3280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_14_0) begin
			b_448_0 <=( io_in_b_14_0) ^ ((fiEnable && (3281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1472_0 <=( io_in_d_14_0) ^ ((fiEnable && (3282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_14_io_in_control_0_shift_b <=( io_in_control_14_0_shift) ^ ((fiEnable && (3283 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_14_io_in_control_0_dataflow_b <=( io_in_control_14_0_dataflow) ^ ((fiEnable && (3284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_14_io_in_control_0_propagate_b <=( io_in_control_14_0_propagate) ^ ((fiEnable && (3285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_14_io_out_valid_0) begin
			b_449_0 <=( _mesh_0_14_io_out_b_0) ^ ((fiEnable && (3286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1473_0 <=( _mesh_0_14_io_out_c_0) ^ ((fiEnable && (3287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_14_io_in_control_0_shift_b <=( _mesh_0_14_io_out_control_0_shift) ^ ((fiEnable && (3288 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_14_io_in_control_0_dataflow_b <=( _mesh_0_14_io_out_control_0_dataflow) ^ ((fiEnable && (3289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_14_io_in_control_0_propagate_b <=( _mesh_0_14_io_out_control_0_propagate) ^ ((fiEnable && (3290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_14_io_out_valid_0) begin
			b_450_0 <=( _mesh_1_14_io_out_b_0) ^ ((fiEnable && (3291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1474_0 <=( _mesh_1_14_io_out_c_0) ^ ((fiEnable && (3292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_14_io_in_control_0_shift_b <=( _mesh_1_14_io_out_control_0_shift) ^ ((fiEnable && (3293 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_14_io_in_control_0_dataflow_b <=( _mesh_1_14_io_out_control_0_dataflow) ^ ((fiEnable && (3294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_14_io_in_control_0_propagate_b <=( _mesh_1_14_io_out_control_0_propagate) ^ ((fiEnable && (3295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_14_io_out_valid_0) begin
			b_451_0 <=( _mesh_2_14_io_out_b_0) ^ ((fiEnable && (3296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1475_0 <=( _mesh_2_14_io_out_c_0) ^ ((fiEnable && (3297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_14_io_in_control_0_shift_b <=( _mesh_2_14_io_out_control_0_shift) ^ ((fiEnable && (3298 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_14_io_in_control_0_dataflow_b <=( _mesh_2_14_io_out_control_0_dataflow) ^ ((fiEnable && (3299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_14_io_in_control_0_propagate_b <=( _mesh_2_14_io_out_control_0_propagate) ^ ((fiEnable && (3300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_14_io_out_valid_0) begin
			b_452_0 <=( _mesh_3_14_io_out_b_0) ^ ((fiEnable && (3301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1476_0 <=( _mesh_3_14_io_out_c_0) ^ ((fiEnable && (3302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_14_io_in_control_0_shift_b <=( _mesh_3_14_io_out_control_0_shift) ^ ((fiEnable && (3303 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_14_io_in_control_0_dataflow_b <=( _mesh_3_14_io_out_control_0_dataflow) ^ ((fiEnable && (3304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_14_io_in_control_0_propagate_b <=( _mesh_3_14_io_out_control_0_propagate) ^ ((fiEnable && (3305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_14_io_out_valid_0) begin
			b_453_0 <=( _mesh_4_14_io_out_b_0) ^ ((fiEnable && (3306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1477_0 <=( _mesh_4_14_io_out_c_0) ^ ((fiEnable && (3307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_14_io_in_control_0_shift_b <=( _mesh_4_14_io_out_control_0_shift) ^ ((fiEnable && (3308 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_14_io_in_control_0_dataflow_b <=( _mesh_4_14_io_out_control_0_dataflow) ^ ((fiEnable && (3309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_14_io_in_control_0_propagate_b <=( _mesh_4_14_io_out_control_0_propagate) ^ ((fiEnable && (3310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_14_io_out_valid_0) begin
			b_454_0 <=( _mesh_5_14_io_out_b_0) ^ ((fiEnable && (3311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1478_0 <=( _mesh_5_14_io_out_c_0) ^ ((fiEnable && (3312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_14_io_in_control_0_shift_b <=( _mesh_5_14_io_out_control_0_shift) ^ ((fiEnable && (3313 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_14_io_in_control_0_dataflow_b <=( _mesh_5_14_io_out_control_0_dataflow) ^ ((fiEnable && (3314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_14_io_in_control_0_propagate_b <=( _mesh_5_14_io_out_control_0_propagate) ^ ((fiEnable && (3315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_14_io_out_valid_0) begin
			b_455_0 <=( _mesh_6_14_io_out_b_0) ^ ((fiEnable && (3316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1479_0 <=( _mesh_6_14_io_out_c_0) ^ ((fiEnable && (3317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_14_io_in_control_0_shift_b <=( _mesh_6_14_io_out_control_0_shift) ^ ((fiEnable && (3318 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_14_io_in_control_0_dataflow_b <=( _mesh_6_14_io_out_control_0_dataflow) ^ ((fiEnable && (3319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_14_io_in_control_0_propagate_b <=( _mesh_6_14_io_out_control_0_propagate) ^ ((fiEnable && (3320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_14_io_out_valid_0) begin
			b_456_0 <=( _mesh_7_14_io_out_b_0) ^ ((fiEnable && (3321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1480_0 <=( _mesh_7_14_io_out_c_0) ^ ((fiEnable && (3322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_14_io_in_control_0_shift_b <=( _mesh_7_14_io_out_control_0_shift) ^ ((fiEnable && (3323 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_14_io_in_control_0_dataflow_b <=( _mesh_7_14_io_out_control_0_dataflow) ^ ((fiEnable && (3324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_14_io_in_control_0_propagate_b <=( _mesh_7_14_io_out_control_0_propagate) ^ ((fiEnable && (3325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_14_io_out_valid_0) begin
			b_457_0 <=( _mesh_8_14_io_out_b_0) ^ ((fiEnable && (3326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1481_0 <=( _mesh_8_14_io_out_c_0) ^ ((fiEnable && (3327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_14_io_in_control_0_shift_b <=( _mesh_8_14_io_out_control_0_shift) ^ ((fiEnable && (3328 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_14_io_in_control_0_dataflow_b <=( _mesh_8_14_io_out_control_0_dataflow) ^ ((fiEnable && (3329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_14_io_in_control_0_propagate_b <=( _mesh_8_14_io_out_control_0_propagate) ^ ((fiEnable && (3330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_14_io_out_valid_0) begin
			b_458_0 <=( _mesh_9_14_io_out_b_0) ^ ((fiEnable && (3331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1482_0 <=( _mesh_9_14_io_out_c_0) ^ ((fiEnable && (3332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_14_io_in_control_0_shift_b <=( _mesh_9_14_io_out_control_0_shift) ^ ((fiEnable && (3333 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_14_io_in_control_0_dataflow_b <=( _mesh_9_14_io_out_control_0_dataflow) ^ ((fiEnable && (3334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_14_io_in_control_0_propagate_b <=( _mesh_9_14_io_out_control_0_propagate) ^ ((fiEnable && (3335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_14_io_out_valid_0) begin
			b_459_0 <=( _mesh_10_14_io_out_b_0) ^ ((fiEnable && (3336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1483_0 <=( _mesh_10_14_io_out_c_0) ^ ((fiEnable && (3337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_14_io_in_control_0_shift_b <=( _mesh_10_14_io_out_control_0_shift) ^ ((fiEnable && (3338 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_14_io_in_control_0_dataflow_b <=( _mesh_10_14_io_out_control_0_dataflow) ^ ((fiEnable && (3339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_14_io_in_control_0_propagate_b <=( _mesh_10_14_io_out_control_0_propagate) ^ ((fiEnable && (3340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_14_io_out_valid_0) begin
			b_460_0 <=( _mesh_11_14_io_out_b_0) ^ ((fiEnable && (3341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1484_0 <=( _mesh_11_14_io_out_c_0) ^ ((fiEnable && (3342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_14_io_in_control_0_shift_b <=( _mesh_11_14_io_out_control_0_shift) ^ ((fiEnable && (3343 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_14_io_in_control_0_dataflow_b <=( _mesh_11_14_io_out_control_0_dataflow) ^ ((fiEnable && (3344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_14_io_in_control_0_propagate_b <=( _mesh_11_14_io_out_control_0_propagate) ^ ((fiEnable && (3345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_14_io_out_valid_0) begin
			b_461_0 <=( _mesh_12_14_io_out_b_0) ^ ((fiEnable && (3346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1485_0 <=( _mesh_12_14_io_out_c_0) ^ ((fiEnable && (3347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_14_io_in_control_0_shift_b <=( _mesh_12_14_io_out_control_0_shift) ^ ((fiEnable && (3348 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_14_io_in_control_0_dataflow_b <=( _mesh_12_14_io_out_control_0_dataflow) ^ ((fiEnable && (3349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_14_io_in_control_0_propagate_b <=( _mesh_12_14_io_out_control_0_propagate) ^ ((fiEnable && (3350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_14_io_out_valid_0) begin
			b_462_0 <=( _mesh_13_14_io_out_b_0) ^ ((fiEnable && (3351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1486_0 <=( _mesh_13_14_io_out_c_0) ^ ((fiEnable && (3352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_14_io_in_control_0_shift_b <=( _mesh_13_14_io_out_control_0_shift) ^ ((fiEnable && (3353 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_14_io_in_control_0_dataflow_b <=( _mesh_13_14_io_out_control_0_dataflow) ^ ((fiEnable && (3354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_14_io_in_control_0_propagate_b <=( _mesh_13_14_io_out_control_0_propagate) ^ ((fiEnable && (3355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_14_io_out_valid_0) begin
			b_463_0 <=( _mesh_14_14_io_out_b_0) ^ ((fiEnable && (3356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1487_0 <=( _mesh_14_14_io_out_c_0) ^ ((fiEnable && (3357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_14_io_in_control_0_shift_b <=( _mesh_14_14_io_out_control_0_shift) ^ ((fiEnable && (3358 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_14_io_in_control_0_dataflow_b <=( _mesh_14_14_io_out_control_0_dataflow) ^ ((fiEnable && (3359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_14_io_in_control_0_propagate_b <=( _mesh_14_14_io_out_control_0_propagate) ^ ((fiEnable && (3360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_14_io_out_valid_0) begin
			b_464_0 <=( _mesh_15_14_io_out_b_0) ^ ((fiEnable && (3361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1488_0 <=( _mesh_15_14_io_out_c_0) ^ ((fiEnable && (3362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_14_io_in_control_0_shift_b <=( _mesh_15_14_io_out_control_0_shift) ^ ((fiEnable && (3363 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_14_io_in_control_0_dataflow_b <=( _mesh_15_14_io_out_control_0_dataflow) ^ ((fiEnable && (3364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_14_io_in_control_0_propagate_b <=( _mesh_15_14_io_out_control_0_propagate) ^ ((fiEnable && (3365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_14_io_out_valid_0) begin
			b_465_0 <=( _mesh_16_14_io_out_b_0) ^ ((fiEnable && (3366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1489_0 <=( _mesh_16_14_io_out_c_0) ^ ((fiEnable && (3367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_14_io_in_control_0_shift_b <=( _mesh_16_14_io_out_control_0_shift) ^ ((fiEnable && (3368 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_14_io_in_control_0_dataflow_b <=( _mesh_16_14_io_out_control_0_dataflow) ^ ((fiEnable && (3369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_14_io_in_control_0_propagate_b <=( _mesh_16_14_io_out_control_0_propagate) ^ ((fiEnable && (3370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_14_io_out_valid_0) begin
			b_466_0 <=( _mesh_17_14_io_out_b_0) ^ ((fiEnable && (3371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1490_0 <=( _mesh_17_14_io_out_c_0) ^ ((fiEnable && (3372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_14_io_in_control_0_shift_b <=( _mesh_17_14_io_out_control_0_shift) ^ ((fiEnable && (3373 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_14_io_in_control_0_dataflow_b <=( _mesh_17_14_io_out_control_0_dataflow) ^ ((fiEnable && (3374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_14_io_in_control_0_propagate_b <=( _mesh_17_14_io_out_control_0_propagate) ^ ((fiEnable && (3375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_14_io_out_valid_0) begin
			b_467_0 <=( _mesh_18_14_io_out_b_0) ^ ((fiEnable && (3376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1491_0 <=( _mesh_18_14_io_out_c_0) ^ ((fiEnable && (3377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_14_io_in_control_0_shift_b <=( _mesh_18_14_io_out_control_0_shift) ^ ((fiEnable && (3378 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_14_io_in_control_0_dataflow_b <=( _mesh_18_14_io_out_control_0_dataflow) ^ ((fiEnable && (3379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_14_io_in_control_0_propagate_b <=( _mesh_18_14_io_out_control_0_propagate) ^ ((fiEnable && (3380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_14_io_out_valid_0) begin
			b_468_0 <=( _mesh_19_14_io_out_b_0) ^ ((fiEnable && (3381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1492_0 <=( _mesh_19_14_io_out_c_0) ^ ((fiEnable && (3382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_14_io_in_control_0_shift_b <=( _mesh_19_14_io_out_control_0_shift) ^ ((fiEnable && (3383 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_14_io_in_control_0_dataflow_b <=( _mesh_19_14_io_out_control_0_dataflow) ^ ((fiEnable && (3384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_14_io_in_control_0_propagate_b <=( _mesh_19_14_io_out_control_0_propagate) ^ ((fiEnable && (3385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_14_io_out_valid_0) begin
			b_469_0 <=( _mesh_20_14_io_out_b_0) ^ ((fiEnable && (3386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1493_0 <=( _mesh_20_14_io_out_c_0) ^ ((fiEnable && (3387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_14_io_in_control_0_shift_b <=( _mesh_20_14_io_out_control_0_shift) ^ ((fiEnable && (3388 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_14_io_in_control_0_dataflow_b <=( _mesh_20_14_io_out_control_0_dataflow) ^ ((fiEnable && (3389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_14_io_in_control_0_propagate_b <=( _mesh_20_14_io_out_control_0_propagate) ^ ((fiEnable && (3390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_14_io_out_valid_0) begin
			b_470_0 <=( _mesh_21_14_io_out_b_0) ^ ((fiEnable && (3391 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1494_0 <=( _mesh_21_14_io_out_c_0) ^ ((fiEnable && (3392 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_14_io_in_control_0_shift_b <=( _mesh_21_14_io_out_control_0_shift) ^ ((fiEnable && (3393 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_14_io_in_control_0_dataflow_b <=( _mesh_21_14_io_out_control_0_dataflow) ^ ((fiEnable && (3394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_14_io_in_control_0_propagate_b <=( _mesh_21_14_io_out_control_0_propagate) ^ ((fiEnable && (3395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_14_io_out_valid_0) begin
			b_471_0 <=( _mesh_22_14_io_out_b_0) ^ ((fiEnable && (3396 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1495_0 <=( _mesh_22_14_io_out_c_0) ^ ((fiEnable && (3397 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_14_io_in_control_0_shift_b <=( _mesh_22_14_io_out_control_0_shift) ^ ((fiEnable && (3398 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_14_io_in_control_0_dataflow_b <=( _mesh_22_14_io_out_control_0_dataflow) ^ ((fiEnable && (3399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_14_io_in_control_0_propagate_b <=( _mesh_22_14_io_out_control_0_propagate) ^ ((fiEnable && (3400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_14_io_out_valid_0) begin
			b_472_0 <=( _mesh_23_14_io_out_b_0) ^ ((fiEnable && (3401 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1496_0 <=( _mesh_23_14_io_out_c_0) ^ ((fiEnable && (3402 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_14_io_in_control_0_shift_b <=( _mesh_23_14_io_out_control_0_shift) ^ ((fiEnable && (3403 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_14_io_in_control_0_dataflow_b <=( _mesh_23_14_io_out_control_0_dataflow) ^ ((fiEnable && (3404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_14_io_in_control_0_propagate_b <=( _mesh_23_14_io_out_control_0_propagate) ^ ((fiEnable && (3405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_14_io_out_valid_0) begin
			b_473_0 <=( _mesh_24_14_io_out_b_0) ^ ((fiEnable && (3406 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1497_0 <=( _mesh_24_14_io_out_c_0) ^ ((fiEnable && (3407 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_14_io_in_control_0_shift_b <=( _mesh_24_14_io_out_control_0_shift) ^ ((fiEnable && (3408 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_14_io_in_control_0_dataflow_b <=( _mesh_24_14_io_out_control_0_dataflow) ^ ((fiEnable && (3409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_14_io_in_control_0_propagate_b <=( _mesh_24_14_io_out_control_0_propagate) ^ ((fiEnable && (3410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_14_io_out_valid_0) begin
			b_474_0 <=( _mesh_25_14_io_out_b_0) ^ ((fiEnable && (3411 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1498_0 <=( _mesh_25_14_io_out_c_0) ^ ((fiEnable && (3412 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_14_io_in_control_0_shift_b <=( _mesh_25_14_io_out_control_0_shift) ^ ((fiEnable && (3413 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_14_io_in_control_0_dataflow_b <=( _mesh_25_14_io_out_control_0_dataflow) ^ ((fiEnable && (3414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_14_io_in_control_0_propagate_b <=( _mesh_25_14_io_out_control_0_propagate) ^ ((fiEnable && (3415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_14_io_out_valid_0) begin
			b_475_0 <=( _mesh_26_14_io_out_b_0) ^ ((fiEnable && (3416 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1499_0 <=( _mesh_26_14_io_out_c_0) ^ ((fiEnable && (3417 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_14_io_in_control_0_shift_b <=( _mesh_26_14_io_out_control_0_shift) ^ ((fiEnable && (3418 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_14_io_in_control_0_dataflow_b <=( _mesh_26_14_io_out_control_0_dataflow) ^ ((fiEnable && (3419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_14_io_in_control_0_propagate_b <=( _mesh_26_14_io_out_control_0_propagate) ^ ((fiEnable && (3420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_14_io_out_valid_0) begin
			b_476_0 <=( _mesh_27_14_io_out_b_0) ^ ((fiEnable && (3421 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1500_0 <=( _mesh_27_14_io_out_c_0) ^ ((fiEnable && (3422 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_14_io_in_control_0_shift_b <=( _mesh_27_14_io_out_control_0_shift) ^ ((fiEnable && (3423 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_14_io_in_control_0_dataflow_b <=( _mesh_27_14_io_out_control_0_dataflow) ^ ((fiEnable && (3424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_14_io_in_control_0_propagate_b <=( _mesh_27_14_io_out_control_0_propagate) ^ ((fiEnable && (3425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_14_io_out_valid_0) begin
			b_477_0 <=( _mesh_28_14_io_out_b_0) ^ ((fiEnable && (3426 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1501_0 <=( _mesh_28_14_io_out_c_0) ^ ((fiEnable && (3427 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_14_io_in_control_0_shift_b <=( _mesh_28_14_io_out_control_0_shift) ^ ((fiEnable && (3428 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_14_io_in_control_0_dataflow_b <=( _mesh_28_14_io_out_control_0_dataflow) ^ ((fiEnable && (3429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_14_io_in_control_0_propagate_b <=( _mesh_28_14_io_out_control_0_propagate) ^ ((fiEnable && (3430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_14_io_out_valid_0) begin
			b_478_0 <=( _mesh_29_14_io_out_b_0) ^ ((fiEnable && (3431 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1502_0 <=( _mesh_29_14_io_out_c_0) ^ ((fiEnable && (3432 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_14_io_in_control_0_shift_b <=( _mesh_29_14_io_out_control_0_shift) ^ ((fiEnable && (3433 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_14_io_in_control_0_dataflow_b <=( _mesh_29_14_io_out_control_0_dataflow) ^ ((fiEnable && (3434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_14_io_in_control_0_propagate_b <=( _mesh_29_14_io_out_control_0_propagate) ^ ((fiEnable && (3435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_14_io_out_valid_0) begin
			b_479_0 <=( _mesh_30_14_io_out_b_0) ^ ((fiEnable && (3436 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1503_0 <=( _mesh_30_14_io_out_c_0) ^ ((fiEnable && (3437 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_14_io_in_control_0_shift_b <=( _mesh_30_14_io_out_control_0_shift) ^ ((fiEnable && (3438 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_14_io_in_control_0_dataflow_b <=( _mesh_30_14_io_out_control_0_dataflow) ^ ((fiEnable && (3439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_14_io_in_control_0_propagate_b <=( _mesh_30_14_io_out_control_0_propagate) ^ ((fiEnable && (3440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_15_0) begin
			b_480_0 <=( io_in_b_15_0) ^ ((fiEnable && (3441 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1504_0 <=( io_in_d_15_0) ^ ((fiEnable && (3442 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_15_io_in_control_0_shift_b <=( io_in_control_15_0_shift) ^ ((fiEnable && (3443 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_15_io_in_control_0_dataflow_b <=( io_in_control_15_0_dataflow) ^ ((fiEnable && (3444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_15_io_in_control_0_propagate_b <=( io_in_control_15_0_propagate) ^ ((fiEnable && (3445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_15_io_out_valid_0) begin
			b_481_0 <=( _mesh_0_15_io_out_b_0) ^ ((fiEnable && (3446 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1505_0 <=( _mesh_0_15_io_out_c_0) ^ ((fiEnable && (3447 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_15_io_in_control_0_shift_b <=( _mesh_0_15_io_out_control_0_shift) ^ ((fiEnable && (3448 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_15_io_in_control_0_dataflow_b <=( _mesh_0_15_io_out_control_0_dataflow) ^ ((fiEnable && (3449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_15_io_in_control_0_propagate_b <=( _mesh_0_15_io_out_control_0_propagate) ^ ((fiEnable && (3450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_15_io_out_valid_0) begin
			b_482_0 <=( _mesh_1_15_io_out_b_0) ^ ((fiEnable && (3451 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1506_0 <=( _mesh_1_15_io_out_c_0) ^ ((fiEnable && (3452 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_15_io_in_control_0_shift_b <=( _mesh_1_15_io_out_control_0_shift) ^ ((fiEnable && (3453 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_15_io_in_control_0_dataflow_b <=( _mesh_1_15_io_out_control_0_dataflow) ^ ((fiEnable && (3454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_15_io_in_control_0_propagate_b <=( _mesh_1_15_io_out_control_0_propagate) ^ ((fiEnable && (3455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_15_io_out_valid_0) begin
			b_483_0 <=( _mesh_2_15_io_out_b_0) ^ ((fiEnable && (3456 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1507_0 <=( _mesh_2_15_io_out_c_0) ^ ((fiEnable && (3457 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_15_io_in_control_0_shift_b <=( _mesh_2_15_io_out_control_0_shift) ^ ((fiEnable && (3458 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_15_io_in_control_0_dataflow_b <=( _mesh_2_15_io_out_control_0_dataflow) ^ ((fiEnable && (3459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_15_io_in_control_0_propagate_b <=( _mesh_2_15_io_out_control_0_propagate) ^ ((fiEnable && (3460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_15_io_out_valid_0) begin
			b_484_0 <=( _mesh_3_15_io_out_b_0) ^ ((fiEnable && (3461 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1508_0 <=( _mesh_3_15_io_out_c_0) ^ ((fiEnable && (3462 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_15_io_in_control_0_shift_b <=( _mesh_3_15_io_out_control_0_shift) ^ ((fiEnable && (3463 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_15_io_in_control_0_dataflow_b <=( _mesh_3_15_io_out_control_0_dataflow) ^ ((fiEnable && (3464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_15_io_in_control_0_propagate_b <=( _mesh_3_15_io_out_control_0_propagate) ^ ((fiEnable && (3465 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_15_io_out_valid_0) begin
			b_485_0 <=( _mesh_4_15_io_out_b_0) ^ ((fiEnable && (3466 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1509_0 <=( _mesh_4_15_io_out_c_0) ^ ((fiEnable && (3467 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_15_io_in_control_0_shift_b <=( _mesh_4_15_io_out_control_0_shift) ^ ((fiEnable && (3468 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_15_io_in_control_0_dataflow_b <=( _mesh_4_15_io_out_control_0_dataflow) ^ ((fiEnable && (3469 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_15_io_in_control_0_propagate_b <=( _mesh_4_15_io_out_control_0_propagate) ^ ((fiEnable && (3470 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_15_io_out_valid_0) begin
			b_486_0 <=( _mesh_5_15_io_out_b_0) ^ ((fiEnable && (3471 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1510_0 <=( _mesh_5_15_io_out_c_0) ^ ((fiEnable && (3472 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_15_io_in_control_0_shift_b <=( _mesh_5_15_io_out_control_0_shift) ^ ((fiEnable && (3473 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_15_io_in_control_0_dataflow_b <=( _mesh_5_15_io_out_control_0_dataflow) ^ ((fiEnable && (3474 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_15_io_in_control_0_propagate_b <=( _mesh_5_15_io_out_control_0_propagate) ^ ((fiEnable && (3475 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_15_io_out_valid_0) begin
			b_487_0 <=( _mesh_6_15_io_out_b_0) ^ ((fiEnable && (3476 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1511_0 <=( _mesh_6_15_io_out_c_0) ^ ((fiEnable && (3477 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_15_io_in_control_0_shift_b <=( _mesh_6_15_io_out_control_0_shift) ^ ((fiEnable && (3478 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_15_io_in_control_0_dataflow_b <=( _mesh_6_15_io_out_control_0_dataflow) ^ ((fiEnable && (3479 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_15_io_in_control_0_propagate_b <=( _mesh_6_15_io_out_control_0_propagate) ^ ((fiEnable && (3480 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_15_io_out_valid_0) begin
			b_488_0 <=( _mesh_7_15_io_out_b_0) ^ ((fiEnable && (3481 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1512_0 <=( _mesh_7_15_io_out_c_0) ^ ((fiEnable && (3482 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_15_io_in_control_0_shift_b <=( _mesh_7_15_io_out_control_0_shift) ^ ((fiEnable && (3483 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_15_io_in_control_0_dataflow_b <=( _mesh_7_15_io_out_control_0_dataflow) ^ ((fiEnable && (3484 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_15_io_in_control_0_propagate_b <=( _mesh_7_15_io_out_control_0_propagate) ^ ((fiEnable && (3485 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_15_io_out_valid_0) begin
			b_489_0 <=( _mesh_8_15_io_out_b_0) ^ ((fiEnable && (3486 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1513_0 <=( _mesh_8_15_io_out_c_0) ^ ((fiEnable && (3487 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_15_io_in_control_0_shift_b <=( _mesh_8_15_io_out_control_0_shift) ^ ((fiEnable && (3488 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_15_io_in_control_0_dataflow_b <=( _mesh_8_15_io_out_control_0_dataflow) ^ ((fiEnable && (3489 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_15_io_in_control_0_propagate_b <=( _mesh_8_15_io_out_control_0_propagate) ^ ((fiEnable && (3490 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_15_io_out_valid_0) begin
			b_490_0 <=( _mesh_9_15_io_out_b_0) ^ ((fiEnable && (3491 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1514_0 <=( _mesh_9_15_io_out_c_0) ^ ((fiEnable && (3492 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_15_io_in_control_0_shift_b <=( _mesh_9_15_io_out_control_0_shift) ^ ((fiEnable && (3493 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_15_io_in_control_0_dataflow_b <=( _mesh_9_15_io_out_control_0_dataflow) ^ ((fiEnable && (3494 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_15_io_in_control_0_propagate_b <=( _mesh_9_15_io_out_control_0_propagate) ^ ((fiEnable && (3495 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_15_io_out_valid_0) begin
			b_491_0 <=( _mesh_10_15_io_out_b_0) ^ ((fiEnable && (3496 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1515_0 <=( _mesh_10_15_io_out_c_0) ^ ((fiEnable && (3497 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_15_io_in_control_0_shift_b <=( _mesh_10_15_io_out_control_0_shift) ^ ((fiEnable && (3498 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_15_io_in_control_0_dataflow_b <=( _mesh_10_15_io_out_control_0_dataflow) ^ ((fiEnable && (3499 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_15_io_in_control_0_propagate_b <=( _mesh_10_15_io_out_control_0_propagate) ^ ((fiEnable && (3500 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_15_io_out_valid_0) begin
			b_492_0 <=( _mesh_11_15_io_out_b_0) ^ ((fiEnable && (3501 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1516_0 <=( _mesh_11_15_io_out_c_0) ^ ((fiEnable && (3502 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_15_io_in_control_0_shift_b <=( _mesh_11_15_io_out_control_0_shift) ^ ((fiEnable && (3503 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_15_io_in_control_0_dataflow_b <=( _mesh_11_15_io_out_control_0_dataflow) ^ ((fiEnable && (3504 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_15_io_in_control_0_propagate_b <=( _mesh_11_15_io_out_control_0_propagate) ^ ((fiEnable && (3505 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_15_io_out_valid_0) begin
			b_493_0 <=( _mesh_12_15_io_out_b_0) ^ ((fiEnable && (3506 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1517_0 <=( _mesh_12_15_io_out_c_0) ^ ((fiEnable && (3507 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_15_io_in_control_0_shift_b <=( _mesh_12_15_io_out_control_0_shift) ^ ((fiEnable && (3508 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_15_io_in_control_0_dataflow_b <=( _mesh_12_15_io_out_control_0_dataflow) ^ ((fiEnable && (3509 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_15_io_in_control_0_propagate_b <=( _mesh_12_15_io_out_control_0_propagate) ^ ((fiEnable && (3510 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_15_io_out_valid_0) begin
			b_494_0 <=( _mesh_13_15_io_out_b_0) ^ ((fiEnable && (3511 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1518_0 <=( _mesh_13_15_io_out_c_0) ^ ((fiEnable && (3512 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_15_io_in_control_0_shift_b <=( _mesh_13_15_io_out_control_0_shift) ^ ((fiEnable && (3513 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_15_io_in_control_0_dataflow_b <=( _mesh_13_15_io_out_control_0_dataflow) ^ ((fiEnable && (3514 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_15_io_in_control_0_propagate_b <=( _mesh_13_15_io_out_control_0_propagate) ^ ((fiEnable && (3515 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_15_io_out_valid_0) begin
			b_495_0 <=( _mesh_14_15_io_out_b_0) ^ ((fiEnable && (3516 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1519_0 <=( _mesh_14_15_io_out_c_0) ^ ((fiEnable && (3517 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_15_io_in_control_0_shift_b <=( _mesh_14_15_io_out_control_0_shift) ^ ((fiEnable && (3518 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_15_io_in_control_0_dataflow_b <=( _mesh_14_15_io_out_control_0_dataflow) ^ ((fiEnable && (3519 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_15_io_in_control_0_propagate_b <=( _mesh_14_15_io_out_control_0_propagate) ^ ((fiEnable && (3520 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_15_io_out_valid_0) begin
			b_496_0 <=( _mesh_15_15_io_out_b_0) ^ ((fiEnable && (3521 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1520_0 <=( _mesh_15_15_io_out_c_0) ^ ((fiEnable && (3522 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_15_io_in_control_0_shift_b <=( _mesh_15_15_io_out_control_0_shift) ^ ((fiEnable && (3523 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_15_io_in_control_0_dataflow_b <=( _mesh_15_15_io_out_control_0_dataflow) ^ ((fiEnable && (3524 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_15_io_in_control_0_propagate_b <=( _mesh_15_15_io_out_control_0_propagate) ^ ((fiEnable && (3525 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_15_io_out_valid_0) begin
			b_497_0 <=( _mesh_16_15_io_out_b_0) ^ ((fiEnable && (3526 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1521_0 <=( _mesh_16_15_io_out_c_0) ^ ((fiEnable && (3527 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_15_io_in_control_0_shift_b <=( _mesh_16_15_io_out_control_0_shift) ^ ((fiEnable && (3528 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_15_io_in_control_0_dataflow_b <=( _mesh_16_15_io_out_control_0_dataflow) ^ ((fiEnable && (3529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_15_io_in_control_0_propagate_b <=( _mesh_16_15_io_out_control_0_propagate) ^ ((fiEnable && (3530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_15_io_out_valid_0) begin
			b_498_0 <=( _mesh_17_15_io_out_b_0) ^ ((fiEnable && (3531 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1522_0 <=( _mesh_17_15_io_out_c_0) ^ ((fiEnable && (3532 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_15_io_in_control_0_shift_b <=( _mesh_17_15_io_out_control_0_shift) ^ ((fiEnable && (3533 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_15_io_in_control_0_dataflow_b <=( _mesh_17_15_io_out_control_0_dataflow) ^ ((fiEnable && (3534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_15_io_in_control_0_propagate_b <=( _mesh_17_15_io_out_control_0_propagate) ^ ((fiEnable && (3535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_15_io_out_valid_0) begin
			b_499_0 <=( _mesh_18_15_io_out_b_0) ^ ((fiEnable && (3536 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1523_0 <=( _mesh_18_15_io_out_c_0) ^ ((fiEnable && (3537 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_15_io_in_control_0_shift_b <=( _mesh_18_15_io_out_control_0_shift) ^ ((fiEnable && (3538 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_15_io_in_control_0_dataflow_b <=( _mesh_18_15_io_out_control_0_dataflow) ^ ((fiEnable && (3539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_15_io_in_control_0_propagate_b <=( _mesh_18_15_io_out_control_0_propagate) ^ ((fiEnable && (3540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_15_io_out_valid_0) begin
			b_500_0 <=( _mesh_19_15_io_out_b_0) ^ ((fiEnable && (3541 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1524_0 <=( _mesh_19_15_io_out_c_0) ^ ((fiEnable && (3542 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_15_io_in_control_0_shift_b <=( _mesh_19_15_io_out_control_0_shift) ^ ((fiEnable && (3543 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_15_io_in_control_0_dataflow_b <=( _mesh_19_15_io_out_control_0_dataflow) ^ ((fiEnable && (3544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_15_io_in_control_0_propagate_b <=( _mesh_19_15_io_out_control_0_propagate) ^ ((fiEnable && (3545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_15_io_out_valid_0) begin
			b_501_0 <=( _mesh_20_15_io_out_b_0) ^ ((fiEnable && (3546 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1525_0 <=( _mesh_20_15_io_out_c_0) ^ ((fiEnable && (3547 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_15_io_in_control_0_shift_b <=( _mesh_20_15_io_out_control_0_shift) ^ ((fiEnable && (3548 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_15_io_in_control_0_dataflow_b <=( _mesh_20_15_io_out_control_0_dataflow) ^ ((fiEnable && (3549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_15_io_in_control_0_propagate_b <=( _mesh_20_15_io_out_control_0_propagate) ^ ((fiEnable && (3550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_15_io_out_valid_0) begin
			b_502_0 <=( _mesh_21_15_io_out_b_0) ^ ((fiEnable && (3551 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1526_0 <=( _mesh_21_15_io_out_c_0) ^ ((fiEnable && (3552 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_15_io_in_control_0_shift_b <=( _mesh_21_15_io_out_control_0_shift) ^ ((fiEnable && (3553 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_15_io_in_control_0_dataflow_b <=( _mesh_21_15_io_out_control_0_dataflow) ^ ((fiEnable && (3554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_15_io_in_control_0_propagate_b <=( _mesh_21_15_io_out_control_0_propagate) ^ ((fiEnable && (3555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_15_io_out_valid_0) begin
			b_503_0 <=( _mesh_22_15_io_out_b_0) ^ ((fiEnable && (3556 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1527_0 <=( _mesh_22_15_io_out_c_0) ^ ((fiEnable && (3557 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_15_io_in_control_0_shift_b <=( _mesh_22_15_io_out_control_0_shift) ^ ((fiEnable && (3558 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_15_io_in_control_0_dataflow_b <=( _mesh_22_15_io_out_control_0_dataflow) ^ ((fiEnable && (3559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_15_io_in_control_0_propagate_b <=( _mesh_22_15_io_out_control_0_propagate) ^ ((fiEnable && (3560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_15_io_out_valid_0) begin
			b_504_0 <=( _mesh_23_15_io_out_b_0) ^ ((fiEnable && (3561 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1528_0 <=( _mesh_23_15_io_out_c_0) ^ ((fiEnable && (3562 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_15_io_in_control_0_shift_b <=( _mesh_23_15_io_out_control_0_shift) ^ ((fiEnable && (3563 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_15_io_in_control_0_dataflow_b <=( _mesh_23_15_io_out_control_0_dataflow) ^ ((fiEnable && (3564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_15_io_in_control_0_propagate_b <=( _mesh_23_15_io_out_control_0_propagate) ^ ((fiEnable && (3565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_15_io_out_valid_0) begin
			b_505_0 <=( _mesh_24_15_io_out_b_0) ^ ((fiEnable && (3566 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1529_0 <=( _mesh_24_15_io_out_c_0) ^ ((fiEnable && (3567 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_15_io_in_control_0_shift_b <=( _mesh_24_15_io_out_control_0_shift) ^ ((fiEnable && (3568 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_15_io_in_control_0_dataflow_b <=( _mesh_24_15_io_out_control_0_dataflow) ^ ((fiEnable && (3569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_15_io_in_control_0_propagate_b <=( _mesh_24_15_io_out_control_0_propagate) ^ ((fiEnable && (3570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_15_io_out_valid_0) begin
			b_506_0 <=( _mesh_25_15_io_out_b_0) ^ ((fiEnable && (3571 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1530_0 <=( _mesh_25_15_io_out_c_0) ^ ((fiEnable && (3572 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_15_io_in_control_0_shift_b <=( _mesh_25_15_io_out_control_0_shift) ^ ((fiEnable && (3573 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_15_io_in_control_0_dataflow_b <=( _mesh_25_15_io_out_control_0_dataflow) ^ ((fiEnable && (3574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_15_io_in_control_0_propagate_b <=( _mesh_25_15_io_out_control_0_propagate) ^ ((fiEnable && (3575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_15_io_out_valid_0) begin
			b_507_0 <=( _mesh_26_15_io_out_b_0) ^ ((fiEnable && (3576 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1531_0 <=( _mesh_26_15_io_out_c_0) ^ ((fiEnable && (3577 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_15_io_in_control_0_shift_b <=( _mesh_26_15_io_out_control_0_shift) ^ ((fiEnable && (3578 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_15_io_in_control_0_dataflow_b <=( _mesh_26_15_io_out_control_0_dataflow) ^ ((fiEnable && (3579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_15_io_in_control_0_propagate_b <=( _mesh_26_15_io_out_control_0_propagate) ^ ((fiEnable && (3580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_15_io_out_valid_0) begin
			b_508_0 <=( _mesh_27_15_io_out_b_0) ^ ((fiEnable && (3581 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1532_0 <=( _mesh_27_15_io_out_c_0) ^ ((fiEnable && (3582 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_15_io_in_control_0_shift_b <=( _mesh_27_15_io_out_control_0_shift) ^ ((fiEnable && (3583 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_15_io_in_control_0_dataflow_b <=( _mesh_27_15_io_out_control_0_dataflow) ^ ((fiEnable && (3584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_15_io_in_control_0_propagate_b <=( _mesh_27_15_io_out_control_0_propagate) ^ ((fiEnable && (3585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_15_io_out_valid_0) begin
			b_509_0 <=( _mesh_28_15_io_out_b_0) ^ ((fiEnable && (3586 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1533_0 <=( _mesh_28_15_io_out_c_0) ^ ((fiEnable && (3587 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_15_io_in_control_0_shift_b <=( _mesh_28_15_io_out_control_0_shift) ^ ((fiEnable && (3588 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_15_io_in_control_0_dataflow_b <=( _mesh_28_15_io_out_control_0_dataflow) ^ ((fiEnable && (3589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_15_io_in_control_0_propagate_b <=( _mesh_28_15_io_out_control_0_propagate) ^ ((fiEnable && (3590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_15_io_out_valid_0) begin
			b_510_0 <=( _mesh_29_15_io_out_b_0) ^ ((fiEnable && (3591 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1534_0 <=( _mesh_29_15_io_out_c_0) ^ ((fiEnable && (3592 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_15_io_in_control_0_shift_b <=( _mesh_29_15_io_out_control_0_shift) ^ ((fiEnable && (3593 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_15_io_in_control_0_dataflow_b <=( _mesh_29_15_io_out_control_0_dataflow) ^ ((fiEnable && (3594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_15_io_in_control_0_propagate_b <=( _mesh_29_15_io_out_control_0_propagate) ^ ((fiEnable && (3595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_15_io_out_valid_0) begin
			b_511_0 <=( _mesh_30_15_io_out_b_0) ^ ((fiEnable && (3596 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1535_0 <=( _mesh_30_15_io_out_c_0) ^ ((fiEnable && (3597 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_15_io_in_control_0_shift_b <=( _mesh_30_15_io_out_control_0_shift) ^ ((fiEnable && (3598 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_15_io_in_control_0_dataflow_b <=( _mesh_30_15_io_out_control_0_dataflow) ^ ((fiEnable && (3599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_15_io_in_control_0_propagate_b <=( _mesh_30_15_io_out_control_0_propagate) ^ ((fiEnable && (3600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_16_0) begin
			b_512_0 <=( io_in_b_16_0) ^ ((fiEnable && (3601 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1536_0 <=( io_in_d_16_0) ^ ((fiEnable && (3602 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_16_io_in_control_0_shift_b <=( io_in_control_16_0_shift) ^ ((fiEnable && (3603 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_16_io_in_control_0_dataflow_b <=( io_in_control_16_0_dataflow) ^ ((fiEnable && (3604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_16_io_in_control_0_propagate_b <=( io_in_control_16_0_propagate) ^ ((fiEnable && (3605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_16_io_out_valid_0) begin
			b_513_0 <=( _mesh_0_16_io_out_b_0) ^ ((fiEnable && (3606 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1537_0 <=( _mesh_0_16_io_out_c_0) ^ ((fiEnable && (3607 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_16_io_in_control_0_shift_b <=( _mesh_0_16_io_out_control_0_shift) ^ ((fiEnable && (3608 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_16_io_in_control_0_dataflow_b <=( _mesh_0_16_io_out_control_0_dataflow) ^ ((fiEnable && (3609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_16_io_in_control_0_propagate_b <=( _mesh_0_16_io_out_control_0_propagate) ^ ((fiEnable && (3610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_16_io_out_valid_0) begin
			b_514_0 <=( _mesh_1_16_io_out_b_0) ^ ((fiEnable && (3611 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1538_0 <=( _mesh_1_16_io_out_c_0) ^ ((fiEnable && (3612 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_16_io_in_control_0_shift_b <=( _mesh_1_16_io_out_control_0_shift) ^ ((fiEnable && (3613 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_16_io_in_control_0_dataflow_b <=( _mesh_1_16_io_out_control_0_dataflow) ^ ((fiEnable && (3614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_16_io_in_control_0_propagate_b <=( _mesh_1_16_io_out_control_0_propagate) ^ ((fiEnable && (3615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_16_io_out_valid_0) begin
			b_515_0 <=( _mesh_2_16_io_out_b_0) ^ ((fiEnable && (3616 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1539_0 <=( _mesh_2_16_io_out_c_0) ^ ((fiEnable && (3617 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_16_io_in_control_0_shift_b <=( _mesh_2_16_io_out_control_0_shift) ^ ((fiEnable && (3618 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_16_io_in_control_0_dataflow_b <=( _mesh_2_16_io_out_control_0_dataflow) ^ ((fiEnable && (3619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_16_io_in_control_0_propagate_b <=( _mesh_2_16_io_out_control_0_propagate) ^ ((fiEnable && (3620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_16_io_out_valid_0) begin
			b_516_0 <=( _mesh_3_16_io_out_b_0) ^ ((fiEnable && (3621 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1540_0 <=( _mesh_3_16_io_out_c_0) ^ ((fiEnable && (3622 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_16_io_in_control_0_shift_b <=( _mesh_3_16_io_out_control_0_shift) ^ ((fiEnable && (3623 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_16_io_in_control_0_dataflow_b <=( _mesh_3_16_io_out_control_0_dataflow) ^ ((fiEnable && (3624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_16_io_in_control_0_propagate_b <=( _mesh_3_16_io_out_control_0_propagate) ^ ((fiEnable && (3625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_16_io_out_valid_0) begin
			b_517_0 <=( _mesh_4_16_io_out_b_0) ^ ((fiEnable && (3626 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1541_0 <=( _mesh_4_16_io_out_c_0) ^ ((fiEnable && (3627 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_16_io_in_control_0_shift_b <=( _mesh_4_16_io_out_control_0_shift) ^ ((fiEnable && (3628 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_16_io_in_control_0_dataflow_b <=( _mesh_4_16_io_out_control_0_dataflow) ^ ((fiEnable && (3629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_16_io_in_control_0_propagate_b <=( _mesh_4_16_io_out_control_0_propagate) ^ ((fiEnable && (3630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_16_io_out_valid_0) begin
			b_518_0 <=( _mesh_5_16_io_out_b_0) ^ ((fiEnable && (3631 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1542_0 <=( _mesh_5_16_io_out_c_0) ^ ((fiEnable && (3632 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_16_io_in_control_0_shift_b <=( _mesh_5_16_io_out_control_0_shift) ^ ((fiEnable && (3633 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_16_io_in_control_0_dataflow_b <=( _mesh_5_16_io_out_control_0_dataflow) ^ ((fiEnable && (3634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_16_io_in_control_0_propagate_b <=( _mesh_5_16_io_out_control_0_propagate) ^ ((fiEnable && (3635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_16_io_out_valid_0) begin
			b_519_0 <=( _mesh_6_16_io_out_b_0) ^ ((fiEnable && (3636 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1543_0 <=( _mesh_6_16_io_out_c_0) ^ ((fiEnable && (3637 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_16_io_in_control_0_shift_b <=( _mesh_6_16_io_out_control_0_shift) ^ ((fiEnable && (3638 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_16_io_in_control_0_dataflow_b <=( _mesh_6_16_io_out_control_0_dataflow) ^ ((fiEnable && (3639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_16_io_in_control_0_propagate_b <=( _mesh_6_16_io_out_control_0_propagate) ^ ((fiEnable && (3640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_16_io_out_valid_0) begin
			b_520_0 <=( _mesh_7_16_io_out_b_0) ^ ((fiEnable && (3641 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1544_0 <=( _mesh_7_16_io_out_c_0) ^ ((fiEnable && (3642 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_16_io_in_control_0_shift_b <=( _mesh_7_16_io_out_control_0_shift) ^ ((fiEnable && (3643 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_16_io_in_control_0_dataflow_b <=( _mesh_7_16_io_out_control_0_dataflow) ^ ((fiEnable && (3644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_16_io_in_control_0_propagate_b <=( _mesh_7_16_io_out_control_0_propagate) ^ ((fiEnable && (3645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_16_io_out_valid_0) begin
			b_521_0 <=( _mesh_8_16_io_out_b_0) ^ ((fiEnable && (3646 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1545_0 <=( _mesh_8_16_io_out_c_0) ^ ((fiEnable && (3647 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_16_io_in_control_0_shift_b <=( _mesh_8_16_io_out_control_0_shift) ^ ((fiEnable && (3648 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_16_io_in_control_0_dataflow_b <=( _mesh_8_16_io_out_control_0_dataflow) ^ ((fiEnable && (3649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_16_io_in_control_0_propagate_b <=( _mesh_8_16_io_out_control_0_propagate) ^ ((fiEnable && (3650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_16_io_out_valid_0) begin
			b_522_0 <=( _mesh_9_16_io_out_b_0) ^ ((fiEnable && (3651 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1546_0 <=( _mesh_9_16_io_out_c_0) ^ ((fiEnable && (3652 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_16_io_in_control_0_shift_b <=( _mesh_9_16_io_out_control_0_shift) ^ ((fiEnable && (3653 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_16_io_in_control_0_dataflow_b <=( _mesh_9_16_io_out_control_0_dataflow) ^ ((fiEnable && (3654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_16_io_in_control_0_propagate_b <=( _mesh_9_16_io_out_control_0_propagate) ^ ((fiEnable && (3655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_16_io_out_valid_0) begin
			b_523_0 <=( _mesh_10_16_io_out_b_0) ^ ((fiEnable && (3656 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1547_0 <=( _mesh_10_16_io_out_c_0) ^ ((fiEnable && (3657 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_16_io_in_control_0_shift_b <=( _mesh_10_16_io_out_control_0_shift) ^ ((fiEnable && (3658 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_16_io_in_control_0_dataflow_b <=( _mesh_10_16_io_out_control_0_dataflow) ^ ((fiEnable && (3659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_16_io_in_control_0_propagate_b <=( _mesh_10_16_io_out_control_0_propagate) ^ ((fiEnable && (3660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_16_io_out_valid_0) begin
			b_524_0 <=( _mesh_11_16_io_out_b_0) ^ ((fiEnable && (3661 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1548_0 <=( _mesh_11_16_io_out_c_0) ^ ((fiEnable && (3662 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_16_io_in_control_0_shift_b <=( _mesh_11_16_io_out_control_0_shift) ^ ((fiEnable && (3663 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_16_io_in_control_0_dataflow_b <=( _mesh_11_16_io_out_control_0_dataflow) ^ ((fiEnable && (3664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_16_io_in_control_0_propagate_b <=( _mesh_11_16_io_out_control_0_propagate) ^ ((fiEnable && (3665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_16_io_out_valid_0) begin
			b_525_0 <=( _mesh_12_16_io_out_b_0) ^ ((fiEnable && (3666 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1549_0 <=( _mesh_12_16_io_out_c_0) ^ ((fiEnable && (3667 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_16_io_in_control_0_shift_b <=( _mesh_12_16_io_out_control_0_shift) ^ ((fiEnable && (3668 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_16_io_in_control_0_dataflow_b <=( _mesh_12_16_io_out_control_0_dataflow) ^ ((fiEnable && (3669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_16_io_in_control_0_propagate_b <=( _mesh_12_16_io_out_control_0_propagate) ^ ((fiEnable && (3670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_16_io_out_valid_0) begin
			b_526_0 <=( _mesh_13_16_io_out_b_0) ^ ((fiEnable && (3671 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1550_0 <=( _mesh_13_16_io_out_c_0) ^ ((fiEnable && (3672 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_16_io_in_control_0_shift_b <=( _mesh_13_16_io_out_control_0_shift) ^ ((fiEnable && (3673 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_16_io_in_control_0_dataflow_b <=( _mesh_13_16_io_out_control_0_dataflow) ^ ((fiEnable && (3674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_16_io_in_control_0_propagate_b <=( _mesh_13_16_io_out_control_0_propagate) ^ ((fiEnable && (3675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_16_io_out_valid_0) begin
			b_527_0 <=( _mesh_14_16_io_out_b_0) ^ ((fiEnable && (3676 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1551_0 <=( _mesh_14_16_io_out_c_0) ^ ((fiEnable && (3677 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_16_io_in_control_0_shift_b <=( _mesh_14_16_io_out_control_0_shift) ^ ((fiEnable && (3678 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_16_io_in_control_0_dataflow_b <=( _mesh_14_16_io_out_control_0_dataflow) ^ ((fiEnable && (3679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_16_io_in_control_0_propagate_b <=( _mesh_14_16_io_out_control_0_propagate) ^ ((fiEnable && (3680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_16_io_out_valid_0) begin
			b_528_0 <=( _mesh_15_16_io_out_b_0) ^ ((fiEnable && (3681 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1552_0 <=( _mesh_15_16_io_out_c_0) ^ ((fiEnable && (3682 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_16_io_in_control_0_shift_b <=( _mesh_15_16_io_out_control_0_shift) ^ ((fiEnable && (3683 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_16_io_in_control_0_dataflow_b <=( _mesh_15_16_io_out_control_0_dataflow) ^ ((fiEnable && (3684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_16_io_in_control_0_propagate_b <=( _mesh_15_16_io_out_control_0_propagate) ^ ((fiEnable && (3685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_16_io_out_valid_0) begin
			b_529_0 <=( _mesh_16_16_io_out_b_0) ^ ((fiEnable && (3686 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1553_0 <=( _mesh_16_16_io_out_c_0) ^ ((fiEnable && (3687 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_16_io_in_control_0_shift_b <=( _mesh_16_16_io_out_control_0_shift) ^ ((fiEnable && (3688 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_16_io_in_control_0_dataflow_b <=( _mesh_16_16_io_out_control_0_dataflow) ^ ((fiEnable && (3689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_16_io_in_control_0_propagate_b <=( _mesh_16_16_io_out_control_0_propagate) ^ ((fiEnable && (3690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_16_io_out_valid_0) begin
			b_530_0 <=( _mesh_17_16_io_out_b_0) ^ ((fiEnable && (3691 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1554_0 <=( _mesh_17_16_io_out_c_0) ^ ((fiEnable && (3692 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_16_io_in_control_0_shift_b <=( _mesh_17_16_io_out_control_0_shift) ^ ((fiEnable && (3693 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_16_io_in_control_0_dataflow_b <=( _mesh_17_16_io_out_control_0_dataflow) ^ ((fiEnable && (3694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_16_io_in_control_0_propagate_b <=( _mesh_17_16_io_out_control_0_propagate) ^ ((fiEnable && (3695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_16_io_out_valid_0) begin
			b_531_0 <=( _mesh_18_16_io_out_b_0) ^ ((fiEnable && (3696 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1555_0 <=( _mesh_18_16_io_out_c_0) ^ ((fiEnable && (3697 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_16_io_in_control_0_shift_b <=( _mesh_18_16_io_out_control_0_shift) ^ ((fiEnable && (3698 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_16_io_in_control_0_dataflow_b <=( _mesh_18_16_io_out_control_0_dataflow) ^ ((fiEnable && (3699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_16_io_in_control_0_propagate_b <=( _mesh_18_16_io_out_control_0_propagate) ^ ((fiEnable && (3700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_16_io_out_valid_0) begin
			b_532_0 <=( _mesh_19_16_io_out_b_0) ^ ((fiEnable && (3701 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1556_0 <=( _mesh_19_16_io_out_c_0) ^ ((fiEnable && (3702 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_16_io_in_control_0_shift_b <=( _mesh_19_16_io_out_control_0_shift) ^ ((fiEnable && (3703 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_16_io_in_control_0_dataflow_b <=( _mesh_19_16_io_out_control_0_dataflow) ^ ((fiEnable && (3704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_16_io_in_control_0_propagate_b <=( _mesh_19_16_io_out_control_0_propagate) ^ ((fiEnable && (3705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_16_io_out_valid_0) begin
			b_533_0 <=( _mesh_20_16_io_out_b_0) ^ ((fiEnable && (3706 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1557_0 <=( _mesh_20_16_io_out_c_0) ^ ((fiEnable && (3707 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_16_io_in_control_0_shift_b <=( _mesh_20_16_io_out_control_0_shift) ^ ((fiEnable && (3708 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_16_io_in_control_0_dataflow_b <=( _mesh_20_16_io_out_control_0_dataflow) ^ ((fiEnable && (3709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_16_io_in_control_0_propagate_b <=( _mesh_20_16_io_out_control_0_propagate) ^ ((fiEnable && (3710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_16_io_out_valid_0) begin
			b_534_0 <=( _mesh_21_16_io_out_b_0) ^ ((fiEnable && (3711 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1558_0 <=( _mesh_21_16_io_out_c_0) ^ ((fiEnable && (3712 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_16_io_in_control_0_shift_b <=( _mesh_21_16_io_out_control_0_shift) ^ ((fiEnable && (3713 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_16_io_in_control_0_dataflow_b <=( _mesh_21_16_io_out_control_0_dataflow) ^ ((fiEnable && (3714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_16_io_in_control_0_propagate_b <=( _mesh_21_16_io_out_control_0_propagate) ^ ((fiEnable && (3715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_16_io_out_valid_0) begin
			b_535_0 <=( _mesh_22_16_io_out_b_0) ^ ((fiEnable && (3716 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1559_0 <=( _mesh_22_16_io_out_c_0) ^ ((fiEnable && (3717 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_16_io_in_control_0_shift_b <=( _mesh_22_16_io_out_control_0_shift) ^ ((fiEnable && (3718 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_16_io_in_control_0_dataflow_b <=( _mesh_22_16_io_out_control_0_dataflow) ^ ((fiEnable && (3719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_16_io_in_control_0_propagate_b <=( _mesh_22_16_io_out_control_0_propagate) ^ ((fiEnable && (3720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_16_io_out_valid_0) begin
			b_536_0 <=( _mesh_23_16_io_out_b_0) ^ ((fiEnable && (3721 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1560_0 <=( _mesh_23_16_io_out_c_0) ^ ((fiEnable && (3722 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_16_io_in_control_0_shift_b <=( _mesh_23_16_io_out_control_0_shift) ^ ((fiEnable && (3723 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_16_io_in_control_0_dataflow_b <=( _mesh_23_16_io_out_control_0_dataflow) ^ ((fiEnable && (3724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_16_io_in_control_0_propagate_b <=( _mesh_23_16_io_out_control_0_propagate) ^ ((fiEnable && (3725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_16_io_out_valid_0) begin
			b_537_0 <=( _mesh_24_16_io_out_b_0) ^ ((fiEnable && (3726 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1561_0 <=( _mesh_24_16_io_out_c_0) ^ ((fiEnable && (3727 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_16_io_in_control_0_shift_b <=( _mesh_24_16_io_out_control_0_shift) ^ ((fiEnable && (3728 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_16_io_in_control_0_dataflow_b <=( _mesh_24_16_io_out_control_0_dataflow) ^ ((fiEnable && (3729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_16_io_in_control_0_propagate_b <=( _mesh_24_16_io_out_control_0_propagate) ^ ((fiEnable && (3730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_16_io_out_valid_0) begin
			b_538_0 <=( _mesh_25_16_io_out_b_0) ^ ((fiEnable && (3731 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1562_0 <=( _mesh_25_16_io_out_c_0) ^ ((fiEnable && (3732 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_16_io_in_control_0_shift_b <=( _mesh_25_16_io_out_control_0_shift) ^ ((fiEnable && (3733 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_16_io_in_control_0_dataflow_b <=( _mesh_25_16_io_out_control_0_dataflow) ^ ((fiEnable && (3734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_16_io_in_control_0_propagate_b <=( _mesh_25_16_io_out_control_0_propagate) ^ ((fiEnable && (3735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_16_io_out_valid_0) begin
			b_539_0 <=( _mesh_26_16_io_out_b_0) ^ ((fiEnable && (3736 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1563_0 <=( _mesh_26_16_io_out_c_0) ^ ((fiEnable && (3737 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_16_io_in_control_0_shift_b <=( _mesh_26_16_io_out_control_0_shift) ^ ((fiEnable && (3738 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_16_io_in_control_0_dataflow_b <=( _mesh_26_16_io_out_control_0_dataflow) ^ ((fiEnable && (3739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_16_io_in_control_0_propagate_b <=( _mesh_26_16_io_out_control_0_propagate) ^ ((fiEnable && (3740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_16_io_out_valid_0) begin
			b_540_0 <=( _mesh_27_16_io_out_b_0) ^ ((fiEnable && (3741 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1564_0 <=( _mesh_27_16_io_out_c_0) ^ ((fiEnable && (3742 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_16_io_in_control_0_shift_b <=( _mesh_27_16_io_out_control_0_shift) ^ ((fiEnable && (3743 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_16_io_in_control_0_dataflow_b <=( _mesh_27_16_io_out_control_0_dataflow) ^ ((fiEnable && (3744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_16_io_in_control_0_propagate_b <=( _mesh_27_16_io_out_control_0_propagate) ^ ((fiEnable && (3745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_16_io_out_valid_0) begin
			b_541_0 <=( _mesh_28_16_io_out_b_0) ^ ((fiEnable && (3746 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1565_0 <=( _mesh_28_16_io_out_c_0) ^ ((fiEnable && (3747 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_16_io_in_control_0_shift_b <=( _mesh_28_16_io_out_control_0_shift) ^ ((fiEnable && (3748 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_16_io_in_control_0_dataflow_b <=( _mesh_28_16_io_out_control_0_dataflow) ^ ((fiEnable && (3749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_16_io_in_control_0_propagate_b <=( _mesh_28_16_io_out_control_0_propagate) ^ ((fiEnable && (3750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_16_io_out_valid_0) begin
			b_542_0 <=( _mesh_29_16_io_out_b_0) ^ ((fiEnable && (3751 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1566_0 <=( _mesh_29_16_io_out_c_0) ^ ((fiEnable && (3752 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_16_io_in_control_0_shift_b <=( _mesh_29_16_io_out_control_0_shift) ^ ((fiEnable && (3753 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_16_io_in_control_0_dataflow_b <=( _mesh_29_16_io_out_control_0_dataflow) ^ ((fiEnable && (3754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_16_io_in_control_0_propagate_b <=( _mesh_29_16_io_out_control_0_propagate) ^ ((fiEnable && (3755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_16_io_out_valid_0) begin
			b_543_0 <=( _mesh_30_16_io_out_b_0) ^ ((fiEnable && (3756 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1567_0 <=( _mesh_30_16_io_out_c_0) ^ ((fiEnable && (3757 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_16_io_in_control_0_shift_b <=( _mesh_30_16_io_out_control_0_shift) ^ ((fiEnable && (3758 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_16_io_in_control_0_dataflow_b <=( _mesh_30_16_io_out_control_0_dataflow) ^ ((fiEnable && (3759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_16_io_in_control_0_propagate_b <=( _mesh_30_16_io_out_control_0_propagate) ^ ((fiEnable && (3760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_17_0) begin
			b_544_0 <=( io_in_b_17_0) ^ ((fiEnable && (3761 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1568_0 <=( io_in_d_17_0) ^ ((fiEnable && (3762 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_17_io_in_control_0_shift_b <=( io_in_control_17_0_shift) ^ ((fiEnable && (3763 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_17_io_in_control_0_dataflow_b <=( io_in_control_17_0_dataflow) ^ ((fiEnable && (3764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_17_io_in_control_0_propagate_b <=( io_in_control_17_0_propagate) ^ ((fiEnable && (3765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_17_io_out_valid_0) begin
			b_545_0 <=( _mesh_0_17_io_out_b_0) ^ ((fiEnable && (3766 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1569_0 <=( _mesh_0_17_io_out_c_0) ^ ((fiEnable && (3767 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_17_io_in_control_0_shift_b <=( _mesh_0_17_io_out_control_0_shift) ^ ((fiEnable && (3768 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_17_io_in_control_0_dataflow_b <=( _mesh_0_17_io_out_control_0_dataflow) ^ ((fiEnable && (3769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_17_io_in_control_0_propagate_b <=( _mesh_0_17_io_out_control_0_propagate) ^ ((fiEnable && (3770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_17_io_out_valid_0) begin
			b_546_0 <=( _mesh_1_17_io_out_b_0) ^ ((fiEnable && (3771 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1570_0 <=( _mesh_1_17_io_out_c_0) ^ ((fiEnable && (3772 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_17_io_in_control_0_shift_b <=( _mesh_1_17_io_out_control_0_shift) ^ ((fiEnable && (3773 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_17_io_in_control_0_dataflow_b <=( _mesh_1_17_io_out_control_0_dataflow) ^ ((fiEnable && (3774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_17_io_in_control_0_propagate_b <=( _mesh_1_17_io_out_control_0_propagate) ^ ((fiEnable && (3775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_17_io_out_valid_0) begin
			b_547_0 <=( _mesh_2_17_io_out_b_0) ^ ((fiEnable && (3776 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1571_0 <=( _mesh_2_17_io_out_c_0) ^ ((fiEnable && (3777 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_17_io_in_control_0_shift_b <=( _mesh_2_17_io_out_control_0_shift) ^ ((fiEnable && (3778 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_17_io_in_control_0_dataflow_b <=( _mesh_2_17_io_out_control_0_dataflow) ^ ((fiEnable && (3779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_17_io_in_control_0_propagate_b <=( _mesh_2_17_io_out_control_0_propagate) ^ ((fiEnable && (3780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_17_io_out_valid_0) begin
			b_548_0 <=( _mesh_3_17_io_out_b_0) ^ ((fiEnable && (3781 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1572_0 <=( _mesh_3_17_io_out_c_0) ^ ((fiEnable && (3782 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_17_io_in_control_0_shift_b <=( _mesh_3_17_io_out_control_0_shift) ^ ((fiEnable && (3783 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_17_io_in_control_0_dataflow_b <=( _mesh_3_17_io_out_control_0_dataflow) ^ ((fiEnable && (3784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_17_io_in_control_0_propagate_b <=( _mesh_3_17_io_out_control_0_propagate) ^ ((fiEnable && (3785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_17_io_out_valid_0) begin
			b_549_0 <=( _mesh_4_17_io_out_b_0) ^ ((fiEnable && (3786 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1573_0 <=( _mesh_4_17_io_out_c_0) ^ ((fiEnable && (3787 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_17_io_in_control_0_shift_b <=( _mesh_4_17_io_out_control_0_shift) ^ ((fiEnable && (3788 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_17_io_in_control_0_dataflow_b <=( _mesh_4_17_io_out_control_0_dataflow) ^ ((fiEnable && (3789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_17_io_in_control_0_propagate_b <=( _mesh_4_17_io_out_control_0_propagate) ^ ((fiEnable && (3790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_17_io_out_valid_0) begin
			b_550_0 <=( _mesh_5_17_io_out_b_0) ^ ((fiEnable && (3791 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1574_0 <=( _mesh_5_17_io_out_c_0) ^ ((fiEnable && (3792 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_17_io_in_control_0_shift_b <=( _mesh_5_17_io_out_control_0_shift) ^ ((fiEnable && (3793 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_17_io_in_control_0_dataflow_b <=( _mesh_5_17_io_out_control_0_dataflow) ^ ((fiEnable && (3794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_17_io_in_control_0_propagate_b <=( _mesh_5_17_io_out_control_0_propagate) ^ ((fiEnable && (3795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_17_io_out_valid_0) begin
			b_551_0 <=( _mesh_6_17_io_out_b_0) ^ ((fiEnable && (3796 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1575_0 <=( _mesh_6_17_io_out_c_0) ^ ((fiEnable && (3797 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_17_io_in_control_0_shift_b <=( _mesh_6_17_io_out_control_0_shift) ^ ((fiEnable && (3798 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_17_io_in_control_0_dataflow_b <=( _mesh_6_17_io_out_control_0_dataflow) ^ ((fiEnable && (3799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_17_io_in_control_0_propagate_b <=( _mesh_6_17_io_out_control_0_propagate) ^ ((fiEnable && (3800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_17_io_out_valid_0) begin
			b_552_0 <=( _mesh_7_17_io_out_b_0) ^ ((fiEnable && (3801 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1576_0 <=( _mesh_7_17_io_out_c_0) ^ ((fiEnable && (3802 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_17_io_in_control_0_shift_b <=( _mesh_7_17_io_out_control_0_shift) ^ ((fiEnable && (3803 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_17_io_in_control_0_dataflow_b <=( _mesh_7_17_io_out_control_0_dataflow) ^ ((fiEnable && (3804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_17_io_in_control_0_propagate_b <=( _mesh_7_17_io_out_control_0_propagate) ^ ((fiEnable && (3805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_17_io_out_valid_0) begin
			b_553_0 <=( _mesh_8_17_io_out_b_0) ^ ((fiEnable && (3806 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1577_0 <=( _mesh_8_17_io_out_c_0) ^ ((fiEnable && (3807 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_17_io_in_control_0_shift_b <=( _mesh_8_17_io_out_control_0_shift) ^ ((fiEnable && (3808 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_17_io_in_control_0_dataflow_b <=( _mesh_8_17_io_out_control_0_dataflow) ^ ((fiEnable && (3809 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_17_io_in_control_0_propagate_b <=( _mesh_8_17_io_out_control_0_propagate) ^ ((fiEnable && (3810 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_17_io_out_valid_0) begin
			b_554_0 <=( _mesh_9_17_io_out_b_0) ^ ((fiEnable && (3811 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1578_0 <=( _mesh_9_17_io_out_c_0) ^ ((fiEnable && (3812 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_17_io_in_control_0_shift_b <=( _mesh_9_17_io_out_control_0_shift) ^ ((fiEnable && (3813 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_17_io_in_control_0_dataflow_b <=( _mesh_9_17_io_out_control_0_dataflow) ^ ((fiEnable && (3814 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_17_io_in_control_0_propagate_b <=( _mesh_9_17_io_out_control_0_propagate) ^ ((fiEnable && (3815 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_17_io_out_valid_0) begin
			b_555_0 <=( _mesh_10_17_io_out_b_0) ^ ((fiEnable && (3816 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1579_0 <=( _mesh_10_17_io_out_c_0) ^ ((fiEnable && (3817 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_17_io_in_control_0_shift_b <=( _mesh_10_17_io_out_control_0_shift) ^ ((fiEnable && (3818 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_17_io_in_control_0_dataflow_b <=( _mesh_10_17_io_out_control_0_dataflow) ^ ((fiEnable && (3819 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_17_io_in_control_0_propagate_b <=( _mesh_10_17_io_out_control_0_propagate) ^ ((fiEnable && (3820 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_17_io_out_valid_0) begin
			b_556_0 <=( _mesh_11_17_io_out_b_0) ^ ((fiEnable && (3821 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1580_0 <=( _mesh_11_17_io_out_c_0) ^ ((fiEnable && (3822 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_17_io_in_control_0_shift_b <=( _mesh_11_17_io_out_control_0_shift) ^ ((fiEnable && (3823 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_17_io_in_control_0_dataflow_b <=( _mesh_11_17_io_out_control_0_dataflow) ^ ((fiEnable && (3824 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_17_io_in_control_0_propagate_b <=( _mesh_11_17_io_out_control_0_propagate) ^ ((fiEnable && (3825 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_17_io_out_valid_0) begin
			b_557_0 <=( _mesh_12_17_io_out_b_0) ^ ((fiEnable && (3826 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1581_0 <=( _mesh_12_17_io_out_c_0) ^ ((fiEnable && (3827 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_17_io_in_control_0_shift_b <=( _mesh_12_17_io_out_control_0_shift) ^ ((fiEnable && (3828 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_17_io_in_control_0_dataflow_b <=( _mesh_12_17_io_out_control_0_dataflow) ^ ((fiEnable && (3829 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_17_io_in_control_0_propagate_b <=( _mesh_12_17_io_out_control_0_propagate) ^ ((fiEnable && (3830 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_17_io_out_valid_0) begin
			b_558_0 <=( _mesh_13_17_io_out_b_0) ^ ((fiEnable && (3831 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1582_0 <=( _mesh_13_17_io_out_c_0) ^ ((fiEnable && (3832 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_17_io_in_control_0_shift_b <=( _mesh_13_17_io_out_control_0_shift) ^ ((fiEnable && (3833 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_17_io_in_control_0_dataflow_b <=( _mesh_13_17_io_out_control_0_dataflow) ^ ((fiEnable && (3834 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_17_io_in_control_0_propagate_b <=( _mesh_13_17_io_out_control_0_propagate) ^ ((fiEnable && (3835 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_17_io_out_valid_0) begin
			b_559_0 <=( _mesh_14_17_io_out_b_0) ^ ((fiEnable && (3836 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1583_0 <=( _mesh_14_17_io_out_c_0) ^ ((fiEnable && (3837 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_17_io_in_control_0_shift_b <=( _mesh_14_17_io_out_control_0_shift) ^ ((fiEnable && (3838 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_17_io_in_control_0_dataflow_b <=( _mesh_14_17_io_out_control_0_dataflow) ^ ((fiEnable && (3839 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_17_io_in_control_0_propagate_b <=( _mesh_14_17_io_out_control_0_propagate) ^ ((fiEnable && (3840 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_17_io_out_valid_0) begin
			b_560_0 <=( _mesh_15_17_io_out_b_0) ^ ((fiEnable && (3841 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1584_0 <=( _mesh_15_17_io_out_c_0) ^ ((fiEnable && (3842 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_17_io_in_control_0_shift_b <=( _mesh_15_17_io_out_control_0_shift) ^ ((fiEnable && (3843 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_17_io_in_control_0_dataflow_b <=( _mesh_15_17_io_out_control_0_dataflow) ^ ((fiEnable && (3844 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_17_io_in_control_0_propagate_b <=( _mesh_15_17_io_out_control_0_propagate) ^ ((fiEnable && (3845 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_17_io_out_valid_0) begin
			b_561_0 <=( _mesh_16_17_io_out_b_0) ^ ((fiEnable && (3846 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1585_0 <=( _mesh_16_17_io_out_c_0) ^ ((fiEnable && (3847 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_17_io_in_control_0_shift_b <=( _mesh_16_17_io_out_control_0_shift) ^ ((fiEnable && (3848 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_17_io_in_control_0_dataflow_b <=( _mesh_16_17_io_out_control_0_dataflow) ^ ((fiEnable && (3849 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_17_io_in_control_0_propagate_b <=( _mesh_16_17_io_out_control_0_propagate) ^ ((fiEnable && (3850 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_17_io_out_valid_0) begin
			b_562_0 <=( _mesh_17_17_io_out_b_0) ^ ((fiEnable && (3851 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1586_0 <=( _mesh_17_17_io_out_c_0) ^ ((fiEnable && (3852 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_17_io_in_control_0_shift_b <=( _mesh_17_17_io_out_control_0_shift) ^ ((fiEnable && (3853 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_17_io_in_control_0_dataflow_b <=( _mesh_17_17_io_out_control_0_dataflow) ^ ((fiEnable && (3854 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_17_io_in_control_0_propagate_b <=( _mesh_17_17_io_out_control_0_propagate) ^ ((fiEnable && (3855 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_17_io_out_valid_0) begin
			b_563_0 <=( _mesh_18_17_io_out_b_0) ^ ((fiEnable && (3856 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1587_0 <=( _mesh_18_17_io_out_c_0) ^ ((fiEnable && (3857 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_17_io_in_control_0_shift_b <=( _mesh_18_17_io_out_control_0_shift) ^ ((fiEnable && (3858 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_17_io_in_control_0_dataflow_b <=( _mesh_18_17_io_out_control_0_dataflow) ^ ((fiEnable && (3859 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_17_io_in_control_0_propagate_b <=( _mesh_18_17_io_out_control_0_propagate) ^ ((fiEnable && (3860 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_17_io_out_valid_0) begin
			b_564_0 <=( _mesh_19_17_io_out_b_0) ^ ((fiEnable && (3861 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1588_0 <=( _mesh_19_17_io_out_c_0) ^ ((fiEnable && (3862 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_17_io_in_control_0_shift_b <=( _mesh_19_17_io_out_control_0_shift) ^ ((fiEnable && (3863 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_17_io_in_control_0_dataflow_b <=( _mesh_19_17_io_out_control_0_dataflow) ^ ((fiEnable && (3864 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_17_io_in_control_0_propagate_b <=( _mesh_19_17_io_out_control_0_propagate) ^ ((fiEnable && (3865 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_17_io_out_valid_0) begin
			b_565_0 <=( _mesh_20_17_io_out_b_0) ^ ((fiEnable && (3866 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1589_0 <=( _mesh_20_17_io_out_c_0) ^ ((fiEnable && (3867 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_17_io_in_control_0_shift_b <=( _mesh_20_17_io_out_control_0_shift) ^ ((fiEnable && (3868 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_17_io_in_control_0_dataflow_b <=( _mesh_20_17_io_out_control_0_dataflow) ^ ((fiEnable && (3869 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_17_io_in_control_0_propagate_b <=( _mesh_20_17_io_out_control_0_propagate) ^ ((fiEnable && (3870 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_17_io_out_valid_0) begin
			b_566_0 <=( _mesh_21_17_io_out_b_0) ^ ((fiEnable && (3871 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1590_0 <=( _mesh_21_17_io_out_c_0) ^ ((fiEnable && (3872 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_17_io_in_control_0_shift_b <=( _mesh_21_17_io_out_control_0_shift) ^ ((fiEnable && (3873 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_17_io_in_control_0_dataflow_b <=( _mesh_21_17_io_out_control_0_dataflow) ^ ((fiEnable && (3874 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_17_io_in_control_0_propagate_b <=( _mesh_21_17_io_out_control_0_propagate) ^ ((fiEnable && (3875 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_17_io_out_valid_0) begin
			b_567_0 <=( _mesh_22_17_io_out_b_0) ^ ((fiEnable && (3876 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1591_0 <=( _mesh_22_17_io_out_c_0) ^ ((fiEnable && (3877 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_17_io_in_control_0_shift_b <=( _mesh_22_17_io_out_control_0_shift) ^ ((fiEnable && (3878 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_17_io_in_control_0_dataflow_b <=( _mesh_22_17_io_out_control_0_dataflow) ^ ((fiEnable && (3879 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_17_io_in_control_0_propagate_b <=( _mesh_22_17_io_out_control_0_propagate) ^ ((fiEnable && (3880 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_17_io_out_valid_0) begin
			b_568_0 <=( _mesh_23_17_io_out_b_0) ^ ((fiEnable && (3881 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1592_0 <=( _mesh_23_17_io_out_c_0) ^ ((fiEnable && (3882 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_17_io_in_control_0_shift_b <=( _mesh_23_17_io_out_control_0_shift) ^ ((fiEnable && (3883 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_17_io_in_control_0_dataflow_b <=( _mesh_23_17_io_out_control_0_dataflow) ^ ((fiEnable && (3884 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_17_io_in_control_0_propagate_b <=( _mesh_23_17_io_out_control_0_propagate) ^ ((fiEnable && (3885 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_17_io_out_valid_0) begin
			b_569_0 <=( _mesh_24_17_io_out_b_0) ^ ((fiEnable && (3886 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1593_0 <=( _mesh_24_17_io_out_c_0) ^ ((fiEnable && (3887 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_17_io_in_control_0_shift_b <=( _mesh_24_17_io_out_control_0_shift) ^ ((fiEnable && (3888 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_17_io_in_control_0_dataflow_b <=( _mesh_24_17_io_out_control_0_dataflow) ^ ((fiEnable && (3889 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_17_io_in_control_0_propagate_b <=( _mesh_24_17_io_out_control_0_propagate) ^ ((fiEnable && (3890 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_17_io_out_valid_0) begin
			b_570_0 <=( _mesh_25_17_io_out_b_0) ^ ((fiEnable && (3891 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1594_0 <=( _mesh_25_17_io_out_c_0) ^ ((fiEnable && (3892 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_17_io_in_control_0_shift_b <=( _mesh_25_17_io_out_control_0_shift) ^ ((fiEnable && (3893 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_17_io_in_control_0_dataflow_b <=( _mesh_25_17_io_out_control_0_dataflow) ^ ((fiEnable && (3894 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_17_io_in_control_0_propagate_b <=( _mesh_25_17_io_out_control_0_propagate) ^ ((fiEnable && (3895 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_17_io_out_valid_0) begin
			b_571_0 <=( _mesh_26_17_io_out_b_0) ^ ((fiEnable && (3896 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1595_0 <=( _mesh_26_17_io_out_c_0) ^ ((fiEnable && (3897 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_17_io_in_control_0_shift_b <=( _mesh_26_17_io_out_control_0_shift) ^ ((fiEnable && (3898 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_17_io_in_control_0_dataflow_b <=( _mesh_26_17_io_out_control_0_dataflow) ^ ((fiEnable && (3899 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_17_io_in_control_0_propagate_b <=( _mesh_26_17_io_out_control_0_propagate) ^ ((fiEnable && (3900 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_17_io_out_valid_0) begin
			b_572_0 <=( _mesh_27_17_io_out_b_0) ^ ((fiEnable && (3901 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1596_0 <=( _mesh_27_17_io_out_c_0) ^ ((fiEnable && (3902 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_17_io_in_control_0_shift_b <=( _mesh_27_17_io_out_control_0_shift) ^ ((fiEnable && (3903 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_17_io_in_control_0_dataflow_b <=( _mesh_27_17_io_out_control_0_dataflow) ^ ((fiEnable && (3904 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_17_io_in_control_0_propagate_b <=( _mesh_27_17_io_out_control_0_propagate) ^ ((fiEnable && (3905 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_17_io_out_valid_0) begin
			b_573_0 <=( _mesh_28_17_io_out_b_0) ^ ((fiEnable && (3906 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1597_0 <=( _mesh_28_17_io_out_c_0) ^ ((fiEnable && (3907 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_17_io_in_control_0_shift_b <=( _mesh_28_17_io_out_control_0_shift) ^ ((fiEnable && (3908 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_17_io_in_control_0_dataflow_b <=( _mesh_28_17_io_out_control_0_dataflow) ^ ((fiEnable && (3909 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_17_io_in_control_0_propagate_b <=( _mesh_28_17_io_out_control_0_propagate) ^ ((fiEnable && (3910 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_17_io_out_valid_0) begin
			b_574_0 <=( _mesh_29_17_io_out_b_0) ^ ((fiEnable && (3911 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1598_0 <=( _mesh_29_17_io_out_c_0) ^ ((fiEnable && (3912 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_17_io_in_control_0_shift_b <=( _mesh_29_17_io_out_control_0_shift) ^ ((fiEnable && (3913 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_17_io_in_control_0_dataflow_b <=( _mesh_29_17_io_out_control_0_dataflow) ^ ((fiEnable && (3914 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_17_io_in_control_0_propagate_b <=( _mesh_29_17_io_out_control_0_propagate) ^ ((fiEnable && (3915 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_17_io_out_valid_0) begin
			b_575_0 <=( _mesh_30_17_io_out_b_0) ^ ((fiEnable && (3916 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1599_0 <=( _mesh_30_17_io_out_c_0) ^ ((fiEnable && (3917 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_17_io_in_control_0_shift_b <=( _mesh_30_17_io_out_control_0_shift) ^ ((fiEnable && (3918 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_17_io_in_control_0_dataflow_b <=( _mesh_30_17_io_out_control_0_dataflow) ^ ((fiEnable && (3919 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_17_io_in_control_0_propagate_b <=( _mesh_30_17_io_out_control_0_propagate) ^ ((fiEnable && (3920 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_18_0) begin
			b_576_0 <=( io_in_b_18_0) ^ ((fiEnable && (3921 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1600_0 <=( io_in_d_18_0) ^ ((fiEnable && (3922 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_18_io_in_control_0_shift_b <=( io_in_control_18_0_shift) ^ ((fiEnable && (3923 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_18_io_in_control_0_dataflow_b <=( io_in_control_18_0_dataflow) ^ ((fiEnable && (3924 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_18_io_in_control_0_propagate_b <=( io_in_control_18_0_propagate) ^ ((fiEnable && (3925 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_18_io_out_valid_0) begin
			b_577_0 <=( _mesh_0_18_io_out_b_0) ^ ((fiEnable && (3926 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1601_0 <=( _mesh_0_18_io_out_c_0) ^ ((fiEnable && (3927 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_18_io_in_control_0_shift_b <=( _mesh_0_18_io_out_control_0_shift) ^ ((fiEnable && (3928 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_18_io_in_control_0_dataflow_b <=( _mesh_0_18_io_out_control_0_dataflow) ^ ((fiEnable && (3929 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_18_io_in_control_0_propagate_b <=( _mesh_0_18_io_out_control_0_propagate) ^ ((fiEnable && (3930 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_18_io_out_valid_0) begin
			b_578_0 <=( _mesh_1_18_io_out_b_0) ^ ((fiEnable && (3931 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1602_0 <=( _mesh_1_18_io_out_c_0) ^ ((fiEnable && (3932 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_18_io_in_control_0_shift_b <=( _mesh_1_18_io_out_control_0_shift) ^ ((fiEnable && (3933 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_18_io_in_control_0_dataflow_b <=( _mesh_1_18_io_out_control_0_dataflow) ^ ((fiEnable && (3934 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_18_io_in_control_0_propagate_b <=( _mesh_1_18_io_out_control_0_propagate) ^ ((fiEnable && (3935 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_18_io_out_valid_0) begin
			b_579_0 <=( _mesh_2_18_io_out_b_0) ^ ((fiEnable && (3936 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1603_0 <=( _mesh_2_18_io_out_c_0) ^ ((fiEnable && (3937 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_18_io_in_control_0_shift_b <=( _mesh_2_18_io_out_control_0_shift) ^ ((fiEnable && (3938 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_18_io_in_control_0_dataflow_b <=( _mesh_2_18_io_out_control_0_dataflow) ^ ((fiEnable && (3939 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_18_io_in_control_0_propagate_b <=( _mesh_2_18_io_out_control_0_propagate) ^ ((fiEnable && (3940 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_18_io_out_valid_0) begin
			b_580_0 <=( _mesh_3_18_io_out_b_0) ^ ((fiEnable && (3941 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1604_0 <=( _mesh_3_18_io_out_c_0) ^ ((fiEnable && (3942 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_18_io_in_control_0_shift_b <=( _mesh_3_18_io_out_control_0_shift) ^ ((fiEnable && (3943 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_18_io_in_control_0_dataflow_b <=( _mesh_3_18_io_out_control_0_dataflow) ^ ((fiEnable && (3944 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_18_io_in_control_0_propagate_b <=( _mesh_3_18_io_out_control_0_propagate) ^ ((fiEnable && (3945 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_18_io_out_valid_0) begin
			b_581_0 <=( _mesh_4_18_io_out_b_0) ^ ((fiEnable && (3946 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1605_0 <=( _mesh_4_18_io_out_c_0) ^ ((fiEnable && (3947 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_18_io_in_control_0_shift_b <=( _mesh_4_18_io_out_control_0_shift) ^ ((fiEnable && (3948 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_18_io_in_control_0_dataflow_b <=( _mesh_4_18_io_out_control_0_dataflow) ^ ((fiEnable && (3949 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_18_io_in_control_0_propagate_b <=( _mesh_4_18_io_out_control_0_propagate) ^ ((fiEnable && (3950 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_18_io_out_valid_0) begin
			b_582_0 <=( _mesh_5_18_io_out_b_0) ^ ((fiEnable && (3951 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1606_0 <=( _mesh_5_18_io_out_c_0) ^ ((fiEnable && (3952 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_18_io_in_control_0_shift_b <=( _mesh_5_18_io_out_control_0_shift) ^ ((fiEnable && (3953 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_18_io_in_control_0_dataflow_b <=( _mesh_5_18_io_out_control_0_dataflow) ^ ((fiEnable && (3954 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_18_io_in_control_0_propagate_b <=( _mesh_5_18_io_out_control_0_propagate) ^ ((fiEnable && (3955 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_18_io_out_valid_0) begin
			b_583_0 <=( _mesh_6_18_io_out_b_0) ^ ((fiEnable && (3956 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1607_0 <=( _mesh_6_18_io_out_c_0) ^ ((fiEnable && (3957 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_18_io_in_control_0_shift_b <=( _mesh_6_18_io_out_control_0_shift) ^ ((fiEnable && (3958 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_18_io_in_control_0_dataflow_b <=( _mesh_6_18_io_out_control_0_dataflow) ^ ((fiEnable && (3959 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_18_io_in_control_0_propagate_b <=( _mesh_6_18_io_out_control_0_propagate) ^ ((fiEnable && (3960 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_18_io_out_valid_0) begin
			b_584_0 <=( _mesh_7_18_io_out_b_0) ^ ((fiEnable && (3961 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1608_0 <=( _mesh_7_18_io_out_c_0) ^ ((fiEnable && (3962 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_18_io_in_control_0_shift_b <=( _mesh_7_18_io_out_control_0_shift) ^ ((fiEnable && (3963 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_18_io_in_control_0_dataflow_b <=( _mesh_7_18_io_out_control_0_dataflow) ^ ((fiEnable && (3964 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_18_io_in_control_0_propagate_b <=( _mesh_7_18_io_out_control_0_propagate) ^ ((fiEnable && (3965 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_18_io_out_valid_0) begin
			b_585_0 <=( _mesh_8_18_io_out_b_0) ^ ((fiEnable && (3966 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1609_0 <=( _mesh_8_18_io_out_c_0) ^ ((fiEnable && (3967 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_18_io_in_control_0_shift_b <=( _mesh_8_18_io_out_control_0_shift) ^ ((fiEnable && (3968 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_18_io_in_control_0_dataflow_b <=( _mesh_8_18_io_out_control_0_dataflow) ^ ((fiEnable && (3969 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_18_io_in_control_0_propagate_b <=( _mesh_8_18_io_out_control_0_propagate) ^ ((fiEnable && (3970 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_18_io_out_valid_0) begin
			b_586_0 <=( _mesh_9_18_io_out_b_0) ^ ((fiEnable && (3971 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1610_0 <=( _mesh_9_18_io_out_c_0) ^ ((fiEnable && (3972 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_18_io_in_control_0_shift_b <=( _mesh_9_18_io_out_control_0_shift) ^ ((fiEnable && (3973 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_18_io_in_control_0_dataflow_b <=( _mesh_9_18_io_out_control_0_dataflow) ^ ((fiEnable && (3974 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_18_io_in_control_0_propagate_b <=( _mesh_9_18_io_out_control_0_propagate) ^ ((fiEnable && (3975 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_18_io_out_valid_0) begin
			b_587_0 <=( _mesh_10_18_io_out_b_0) ^ ((fiEnable && (3976 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1611_0 <=( _mesh_10_18_io_out_c_0) ^ ((fiEnable && (3977 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_18_io_in_control_0_shift_b <=( _mesh_10_18_io_out_control_0_shift) ^ ((fiEnable && (3978 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_18_io_in_control_0_dataflow_b <=( _mesh_10_18_io_out_control_0_dataflow) ^ ((fiEnable && (3979 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_18_io_in_control_0_propagate_b <=( _mesh_10_18_io_out_control_0_propagate) ^ ((fiEnable && (3980 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_18_io_out_valid_0) begin
			b_588_0 <=( _mesh_11_18_io_out_b_0) ^ ((fiEnable && (3981 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1612_0 <=( _mesh_11_18_io_out_c_0) ^ ((fiEnable && (3982 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_18_io_in_control_0_shift_b <=( _mesh_11_18_io_out_control_0_shift) ^ ((fiEnable && (3983 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_18_io_in_control_0_dataflow_b <=( _mesh_11_18_io_out_control_0_dataflow) ^ ((fiEnable && (3984 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_18_io_in_control_0_propagate_b <=( _mesh_11_18_io_out_control_0_propagate) ^ ((fiEnable && (3985 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_18_io_out_valid_0) begin
			b_589_0 <=( _mesh_12_18_io_out_b_0) ^ ((fiEnable && (3986 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1613_0 <=( _mesh_12_18_io_out_c_0) ^ ((fiEnable && (3987 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_18_io_in_control_0_shift_b <=( _mesh_12_18_io_out_control_0_shift) ^ ((fiEnable && (3988 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_18_io_in_control_0_dataflow_b <=( _mesh_12_18_io_out_control_0_dataflow) ^ ((fiEnable && (3989 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_18_io_in_control_0_propagate_b <=( _mesh_12_18_io_out_control_0_propagate) ^ ((fiEnable && (3990 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_18_io_out_valid_0) begin
			b_590_0 <=( _mesh_13_18_io_out_b_0) ^ ((fiEnable && (3991 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1614_0 <=( _mesh_13_18_io_out_c_0) ^ ((fiEnable && (3992 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_18_io_in_control_0_shift_b <=( _mesh_13_18_io_out_control_0_shift) ^ ((fiEnable && (3993 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_18_io_in_control_0_dataflow_b <=( _mesh_13_18_io_out_control_0_dataflow) ^ ((fiEnable && (3994 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_18_io_in_control_0_propagate_b <=( _mesh_13_18_io_out_control_0_propagate) ^ ((fiEnable && (3995 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_18_io_out_valid_0) begin
			b_591_0 <=( _mesh_14_18_io_out_b_0) ^ ((fiEnable && (3996 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1615_0 <=( _mesh_14_18_io_out_c_0) ^ ((fiEnable && (3997 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_18_io_in_control_0_shift_b <=( _mesh_14_18_io_out_control_0_shift) ^ ((fiEnable && (3998 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_18_io_in_control_0_dataflow_b <=( _mesh_14_18_io_out_control_0_dataflow) ^ ((fiEnable && (3999 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_18_io_in_control_0_propagate_b <=( _mesh_14_18_io_out_control_0_propagate) ^ ((fiEnable && (4000 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_18_io_out_valid_0) begin
			b_592_0 <=( _mesh_15_18_io_out_b_0) ^ ((fiEnable && (4001 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1616_0 <=( _mesh_15_18_io_out_c_0) ^ ((fiEnable && (4002 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_18_io_in_control_0_shift_b <=( _mesh_15_18_io_out_control_0_shift) ^ ((fiEnable && (4003 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_18_io_in_control_0_dataflow_b <=( _mesh_15_18_io_out_control_0_dataflow) ^ ((fiEnable && (4004 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_18_io_in_control_0_propagate_b <=( _mesh_15_18_io_out_control_0_propagate) ^ ((fiEnable && (4005 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_18_io_out_valid_0) begin
			b_593_0 <=( _mesh_16_18_io_out_b_0) ^ ((fiEnable && (4006 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1617_0 <=( _mesh_16_18_io_out_c_0) ^ ((fiEnable && (4007 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_18_io_in_control_0_shift_b <=( _mesh_16_18_io_out_control_0_shift) ^ ((fiEnable && (4008 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_18_io_in_control_0_dataflow_b <=( _mesh_16_18_io_out_control_0_dataflow) ^ ((fiEnable && (4009 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_18_io_in_control_0_propagate_b <=( _mesh_16_18_io_out_control_0_propagate) ^ ((fiEnable && (4010 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_18_io_out_valid_0) begin
			b_594_0 <=( _mesh_17_18_io_out_b_0) ^ ((fiEnable && (4011 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1618_0 <=( _mesh_17_18_io_out_c_0) ^ ((fiEnable && (4012 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_18_io_in_control_0_shift_b <=( _mesh_17_18_io_out_control_0_shift) ^ ((fiEnable && (4013 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_18_io_in_control_0_dataflow_b <=( _mesh_17_18_io_out_control_0_dataflow) ^ ((fiEnable && (4014 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_18_io_in_control_0_propagate_b <=( _mesh_17_18_io_out_control_0_propagate) ^ ((fiEnable && (4015 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_18_io_out_valid_0) begin
			b_595_0 <=( _mesh_18_18_io_out_b_0) ^ ((fiEnable && (4016 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1619_0 <=( _mesh_18_18_io_out_c_0) ^ ((fiEnable && (4017 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_18_io_in_control_0_shift_b <=( _mesh_18_18_io_out_control_0_shift) ^ ((fiEnable && (4018 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_18_io_in_control_0_dataflow_b <=( _mesh_18_18_io_out_control_0_dataflow) ^ ((fiEnable && (4019 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_18_io_in_control_0_propagate_b <=( _mesh_18_18_io_out_control_0_propagate) ^ ((fiEnable && (4020 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_18_io_out_valid_0) begin
			b_596_0 <=( _mesh_19_18_io_out_b_0) ^ ((fiEnable && (4021 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1620_0 <=( _mesh_19_18_io_out_c_0) ^ ((fiEnable && (4022 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_18_io_in_control_0_shift_b <=( _mesh_19_18_io_out_control_0_shift) ^ ((fiEnable && (4023 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_18_io_in_control_0_dataflow_b <=( _mesh_19_18_io_out_control_0_dataflow) ^ ((fiEnable && (4024 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_18_io_in_control_0_propagate_b <=( _mesh_19_18_io_out_control_0_propagate) ^ ((fiEnable && (4025 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_18_io_out_valid_0) begin
			b_597_0 <=( _mesh_20_18_io_out_b_0) ^ ((fiEnable && (4026 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1621_0 <=( _mesh_20_18_io_out_c_0) ^ ((fiEnable && (4027 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_18_io_in_control_0_shift_b <=( _mesh_20_18_io_out_control_0_shift) ^ ((fiEnable && (4028 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_18_io_in_control_0_dataflow_b <=( _mesh_20_18_io_out_control_0_dataflow) ^ ((fiEnable && (4029 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_18_io_in_control_0_propagate_b <=( _mesh_20_18_io_out_control_0_propagate) ^ ((fiEnable && (4030 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_18_io_out_valid_0) begin
			b_598_0 <=( _mesh_21_18_io_out_b_0) ^ ((fiEnable && (4031 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1622_0 <=( _mesh_21_18_io_out_c_0) ^ ((fiEnable && (4032 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_18_io_in_control_0_shift_b <=( _mesh_21_18_io_out_control_0_shift) ^ ((fiEnable && (4033 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_18_io_in_control_0_dataflow_b <=( _mesh_21_18_io_out_control_0_dataflow) ^ ((fiEnable && (4034 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_18_io_in_control_0_propagate_b <=( _mesh_21_18_io_out_control_0_propagate) ^ ((fiEnable && (4035 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_18_io_out_valid_0) begin
			b_599_0 <=( _mesh_22_18_io_out_b_0) ^ ((fiEnable && (4036 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1623_0 <=( _mesh_22_18_io_out_c_0) ^ ((fiEnable && (4037 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_18_io_in_control_0_shift_b <=( _mesh_22_18_io_out_control_0_shift) ^ ((fiEnable && (4038 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_18_io_in_control_0_dataflow_b <=( _mesh_22_18_io_out_control_0_dataflow) ^ ((fiEnable && (4039 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_18_io_in_control_0_propagate_b <=( _mesh_22_18_io_out_control_0_propagate) ^ ((fiEnable && (4040 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_18_io_out_valid_0) begin
			b_600_0 <=( _mesh_23_18_io_out_b_0) ^ ((fiEnable && (4041 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1624_0 <=( _mesh_23_18_io_out_c_0) ^ ((fiEnable && (4042 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_18_io_in_control_0_shift_b <=( _mesh_23_18_io_out_control_0_shift) ^ ((fiEnable && (4043 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_18_io_in_control_0_dataflow_b <=( _mesh_23_18_io_out_control_0_dataflow) ^ ((fiEnable && (4044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_18_io_in_control_0_propagate_b <=( _mesh_23_18_io_out_control_0_propagate) ^ ((fiEnable && (4045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_18_io_out_valid_0) begin
			b_601_0 <=( _mesh_24_18_io_out_b_0) ^ ((fiEnable && (4046 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1625_0 <=( _mesh_24_18_io_out_c_0) ^ ((fiEnable && (4047 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_18_io_in_control_0_shift_b <=( _mesh_24_18_io_out_control_0_shift) ^ ((fiEnable && (4048 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_18_io_in_control_0_dataflow_b <=( _mesh_24_18_io_out_control_0_dataflow) ^ ((fiEnable && (4049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_18_io_in_control_0_propagate_b <=( _mesh_24_18_io_out_control_0_propagate) ^ ((fiEnable && (4050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_18_io_out_valid_0) begin
			b_602_0 <=( _mesh_25_18_io_out_b_0) ^ ((fiEnable && (4051 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1626_0 <=( _mesh_25_18_io_out_c_0) ^ ((fiEnable && (4052 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_18_io_in_control_0_shift_b <=( _mesh_25_18_io_out_control_0_shift) ^ ((fiEnable && (4053 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_18_io_in_control_0_dataflow_b <=( _mesh_25_18_io_out_control_0_dataflow) ^ ((fiEnable && (4054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_18_io_in_control_0_propagate_b <=( _mesh_25_18_io_out_control_0_propagate) ^ ((fiEnable && (4055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_18_io_out_valid_0) begin
			b_603_0 <=( _mesh_26_18_io_out_b_0) ^ ((fiEnable && (4056 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1627_0 <=( _mesh_26_18_io_out_c_0) ^ ((fiEnable && (4057 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_18_io_in_control_0_shift_b <=( _mesh_26_18_io_out_control_0_shift) ^ ((fiEnable && (4058 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_18_io_in_control_0_dataflow_b <=( _mesh_26_18_io_out_control_0_dataflow) ^ ((fiEnable && (4059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_18_io_in_control_0_propagate_b <=( _mesh_26_18_io_out_control_0_propagate) ^ ((fiEnable && (4060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_18_io_out_valid_0) begin
			b_604_0 <=( _mesh_27_18_io_out_b_0) ^ ((fiEnable && (4061 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1628_0 <=( _mesh_27_18_io_out_c_0) ^ ((fiEnable && (4062 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_18_io_in_control_0_shift_b <=( _mesh_27_18_io_out_control_0_shift) ^ ((fiEnable && (4063 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_18_io_in_control_0_dataflow_b <=( _mesh_27_18_io_out_control_0_dataflow) ^ ((fiEnable && (4064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_18_io_in_control_0_propagate_b <=( _mesh_27_18_io_out_control_0_propagate) ^ ((fiEnable && (4065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_18_io_out_valid_0) begin
			b_605_0 <=( _mesh_28_18_io_out_b_0) ^ ((fiEnable && (4066 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1629_0 <=( _mesh_28_18_io_out_c_0) ^ ((fiEnable && (4067 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_18_io_in_control_0_shift_b <=( _mesh_28_18_io_out_control_0_shift) ^ ((fiEnable && (4068 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_18_io_in_control_0_dataflow_b <=( _mesh_28_18_io_out_control_0_dataflow) ^ ((fiEnable && (4069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_18_io_in_control_0_propagate_b <=( _mesh_28_18_io_out_control_0_propagate) ^ ((fiEnable && (4070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_18_io_out_valid_0) begin
			b_606_0 <=( _mesh_29_18_io_out_b_0) ^ ((fiEnable && (4071 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1630_0 <=( _mesh_29_18_io_out_c_0) ^ ((fiEnable && (4072 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_18_io_in_control_0_shift_b <=( _mesh_29_18_io_out_control_0_shift) ^ ((fiEnable && (4073 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_18_io_in_control_0_dataflow_b <=( _mesh_29_18_io_out_control_0_dataflow) ^ ((fiEnable && (4074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_18_io_in_control_0_propagate_b <=( _mesh_29_18_io_out_control_0_propagate) ^ ((fiEnable && (4075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_18_io_out_valid_0) begin
			b_607_0 <=( _mesh_30_18_io_out_b_0) ^ ((fiEnable && (4076 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1631_0 <=( _mesh_30_18_io_out_c_0) ^ ((fiEnable && (4077 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_18_io_in_control_0_shift_b <=( _mesh_30_18_io_out_control_0_shift) ^ ((fiEnable && (4078 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_18_io_in_control_0_dataflow_b <=( _mesh_30_18_io_out_control_0_dataflow) ^ ((fiEnable && (4079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_18_io_in_control_0_propagate_b <=( _mesh_30_18_io_out_control_0_propagate) ^ ((fiEnable && (4080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_19_0) begin
			b_608_0 <=( io_in_b_19_0) ^ ((fiEnable && (4081 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1632_0 <=( io_in_d_19_0) ^ ((fiEnable && (4082 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_19_io_in_control_0_shift_b <=( io_in_control_19_0_shift) ^ ((fiEnable && (4083 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_19_io_in_control_0_dataflow_b <=( io_in_control_19_0_dataflow) ^ ((fiEnable && (4084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_19_io_in_control_0_propagate_b <=( io_in_control_19_0_propagate) ^ ((fiEnable && (4085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_19_io_out_valid_0) begin
			b_609_0 <=( _mesh_0_19_io_out_b_0) ^ ((fiEnable && (4086 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1633_0 <=( _mesh_0_19_io_out_c_0) ^ ((fiEnable && (4087 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_19_io_in_control_0_shift_b <=( _mesh_0_19_io_out_control_0_shift) ^ ((fiEnable && (4088 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_19_io_in_control_0_dataflow_b <=( _mesh_0_19_io_out_control_0_dataflow) ^ ((fiEnable && (4089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_19_io_in_control_0_propagate_b <=( _mesh_0_19_io_out_control_0_propagate) ^ ((fiEnable && (4090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_19_io_out_valid_0) begin
			b_610_0 <=( _mesh_1_19_io_out_b_0) ^ ((fiEnable && (4091 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1634_0 <=( _mesh_1_19_io_out_c_0) ^ ((fiEnable && (4092 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_19_io_in_control_0_shift_b <=( _mesh_1_19_io_out_control_0_shift) ^ ((fiEnable && (4093 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_19_io_in_control_0_dataflow_b <=( _mesh_1_19_io_out_control_0_dataflow) ^ ((fiEnable && (4094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_19_io_in_control_0_propagate_b <=( _mesh_1_19_io_out_control_0_propagate) ^ ((fiEnable && (4095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_19_io_out_valid_0) begin
			b_611_0 <=( _mesh_2_19_io_out_b_0) ^ ((fiEnable && (4096 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1635_0 <=( _mesh_2_19_io_out_c_0) ^ ((fiEnable && (4097 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_19_io_in_control_0_shift_b <=( _mesh_2_19_io_out_control_0_shift) ^ ((fiEnable && (4098 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_19_io_in_control_0_dataflow_b <=( _mesh_2_19_io_out_control_0_dataflow) ^ ((fiEnable && (4099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_19_io_in_control_0_propagate_b <=( _mesh_2_19_io_out_control_0_propagate) ^ ((fiEnable && (4100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_19_io_out_valid_0) begin
			b_612_0 <=( _mesh_3_19_io_out_b_0) ^ ((fiEnable && (4101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1636_0 <=( _mesh_3_19_io_out_c_0) ^ ((fiEnable && (4102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_19_io_in_control_0_shift_b <=( _mesh_3_19_io_out_control_0_shift) ^ ((fiEnable && (4103 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_19_io_in_control_0_dataflow_b <=( _mesh_3_19_io_out_control_0_dataflow) ^ ((fiEnable && (4104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_19_io_in_control_0_propagate_b <=( _mesh_3_19_io_out_control_0_propagate) ^ ((fiEnable && (4105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_19_io_out_valid_0) begin
			b_613_0 <=( _mesh_4_19_io_out_b_0) ^ ((fiEnable && (4106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1637_0 <=( _mesh_4_19_io_out_c_0) ^ ((fiEnable && (4107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_19_io_in_control_0_shift_b <=( _mesh_4_19_io_out_control_0_shift) ^ ((fiEnable && (4108 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_19_io_in_control_0_dataflow_b <=( _mesh_4_19_io_out_control_0_dataflow) ^ ((fiEnable && (4109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_19_io_in_control_0_propagate_b <=( _mesh_4_19_io_out_control_0_propagate) ^ ((fiEnable && (4110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_19_io_out_valid_0) begin
			b_614_0 <=( _mesh_5_19_io_out_b_0) ^ ((fiEnable && (4111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1638_0 <=( _mesh_5_19_io_out_c_0) ^ ((fiEnable && (4112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_19_io_in_control_0_shift_b <=( _mesh_5_19_io_out_control_0_shift) ^ ((fiEnable && (4113 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_19_io_in_control_0_dataflow_b <=( _mesh_5_19_io_out_control_0_dataflow) ^ ((fiEnable && (4114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_19_io_in_control_0_propagate_b <=( _mesh_5_19_io_out_control_0_propagate) ^ ((fiEnable && (4115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_19_io_out_valid_0) begin
			b_615_0 <=( _mesh_6_19_io_out_b_0) ^ ((fiEnable && (4116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1639_0 <=( _mesh_6_19_io_out_c_0) ^ ((fiEnable && (4117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_19_io_in_control_0_shift_b <=( _mesh_6_19_io_out_control_0_shift) ^ ((fiEnable && (4118 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_19_io_in_control_0_dataflow_b <=( _mesh_6_19_io_out_control_0_dataflow) ^ ((fiEnable && (4119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_19_io_in_control_0_propagate_b <=( _mesh_6_19_io_out_control_0_propagate) ^ ((fiEnable && (4120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_19_io_out_valid_0) begin
			b_616_0 <=( _mesh_7_19_io_out_b_0) ^ ((fiEnable && (4121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1640_0 <=( _mesh_7_19_io_out_c_0) ^ ((fiEnable && (4122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_19_io_in_control_0_shift_b <=( _mesh_7_19_io_out_control_0_shift) ^ ((fiEnable && (4123 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_19_io_in_control_0_dataflow_b <=( _mesh_7_19_io_out_control_0_dataflow) ^ ((fiEnable && (4124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_19_io_in_control_0_propagate_b <=( _mesh_7_19_io_out_control_0_propagate) ^ ((fiEnable && (4125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_19_io_out_valid_0) begin
			b_617_0 <=( _mesh_8_19_io_out_b_0) ^ ((fiEnable && (4126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1641_0 <=( _mesh_8_19_io_out_c_0) ^ ((fiEnable && (4127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_19_io_in_control_0_shift_b <=( _mesh_8_19_io_out_control_0_shift) ^ ((fiEnable && (4128 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_19_io_in_control_0_dataflow_b <=( _mesh_8_19_io_out_control_0_dataflow) ^ ((fiEnable && (4129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_19_io_in_control_0_propagate_b <=( _mesh_8_19_io_out_control_0_propagate) ^ ((fiEnable && (4130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_19_io_out_valid_0) begin
			b_618_0 <=( _mesh_9_19_io_out_b_0) ^ ((fiEnable && (4131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1642_0 <=( _mesh_9_19_io_out_c_0) ^ ((fiEnable && (4132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_19_io_in_control_0_shift_b <=( _mesh_9_19_io_out_control_0_shift) ^ ((fiEnable && (4133 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_19_io_in_control_0_dataflow_b <=( _mesh_9_19_io_out_control_0_dataflow) ^ ((fiEnable && (4134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_19_io_in_control_0_propagate_b <=( _mesh_9_19_io_out_control_0_propagate) ^ ((fiEnable && (4135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_19_io_out_valid_0) begin
			b_619_0 <=( _mesh_10_19_io_out_b_0) ^ ((fiEnable && (4136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1643_0 <=( _mesh_10_19_io_out_c_0) ^ ((fiEnable && (4137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_19_io_in_control_0_shift_b <=( _mesh_10_19_io_out_control_0_shift) ^ ((fiEnable && (4138 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_19_io_in_control_0_dataflow_b <=( _mesh_10_19_io_out_control_0_dataflow) ^ ((fiEnable && (4139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_19_io_in_control_0_propagate_b <=( _mesh_10_19_io_out_control_0_propagate) ^ ((fiEnable && (4140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_19_io_out_valid_0) begin
			b_620_0 <=( _mesh_11_19_io_out_b_0) ^ ((fiEnable && (4141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1644_0 <=( _mesh_11_19_io_out_c_0) ^ ((fiEnable && (4142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_19_io_in_control_0_shift_b <=( _mesh_11_19_io_out_control_0_shift) ^ ((fiEnable && (4143 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_19_io_in_control_0_dataflow_b <=( _mesh_11_19_io_out_control_0_dataflow) ^ ((fiEnable && (4144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_19_io_in_control_0_propagate_b <=( _mesh_11_19_io_out_control_0_propagate) ^ ((fiEnable && (4145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_19_io_out_valid_0) begin
			b_621_0 <=( _mesh_12_19_io_out_b_0) ^ ((fiEnable && (4146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1645_0 <=( _mesh_12_19_io_out_c_0) ^ ((fiEnable && (4147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_19_io_in_control_0_shift_b <=( _mesh_12_19_io_out_control_0_shift) ^ ((fiEnable && (4148 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_19_io_in_control_0_dataflow_b <=( _mesh_12_19_io_out_control_0_dataflow) ^ ((fiEnable && (4149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_19_io_in_control_0_propagate_b <=( _mesh_12_19_io_out_control_0_propagate) ^ ((fiEnable && (4150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_19_io_out_valid_0) begin
			b_622_0 <=( _mesh_13_19_io_out_b_0) ^ ((fiEnable && (4151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1646_0 <=( _mesh_13_19_io_out_c_0) ^ ((fiEnable && (4152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_19_io_in_control_0_shift_b <=( _mesh_13_19_io_out_control_0_shift) ^ ((fiEnable && (4153 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_19_io_in_control_0_dataflow_b <=( _mesh_13_19_io_out_control_0_dataflow) ^ ((fiEnable && (4154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_19_io_in_control_0_propagate_b <=( _mesh_13_19_io_out_control_0_propagate) ^ ((fiEnable && (4155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_19_io_out_valid_0) begin
			b_623_0 <=( _mesh_14_19_io_out_b_0) ^ ((fiEnable && (4156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1647_0 <=( _mesh_14_19_io_out_c_0) ^ ((fiEnable && (4157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_19_io_in_control_0_shift_b <=( _mesh_14_19_io_out_control_0_shift) ^ ((fiEnable && (4158 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_19_io_in_control_0_dataflow_b <=( _mesh_14_19_io_out_control_0_dataflow) ^ ((fiEnable && (4159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_19_io_in_control_0_propagate_b <=( _mesh_14_19_io_out_control_0_propagate) ^ ((fiEnable && (4160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_19_io_out_valid_0) begin
			b_624_0 <=( _mesh_15_19_io_out_b_0) ^ ((fiEnable && (4161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1648_0 <=( _mesh_15_19_io_out_c_0) ^ ((fiEnable && (4162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_19_io_in_control_0_shift_b <=( _mesh_15_19_io_out_control_0_shift) ^ ((fiEnable && (4163 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_19_io_in_control_0_dataflow_b <=( _mesh_15_19_io_out_control_0_dataflow) ^ ((fiEnable && (4164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_19_io_in_control_0_propagate_b <=( _mesh_15_19_io_out_control_0_propagate) ^ ((fiEnable && (4165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_19_io_out_valid_0) begin
			b_625_0 <=( _mesh_16_19_io_out_b_0) ^ ((fiEnable && (4166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1649_0 <=( _mesh_16_19_io_out_c_0) ^ ((fiEnable && (4167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_19_io_in_control_0_shift_b <=( _mesh_16_19_io_out_control_0_shift) ^ ((fiEnable && (4168 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_19_io_in_control_0_dataflow_b <=( _mesh_16_19_io_out_control_0_dataflow) ^ ((fiEnable && (4169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_19_io_in_control_0_propagate_b <=( _mesh_16_19_io_out_control_0_propagate) ^ ((fiEnable && (4170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_19_io_out_valid_0) begin
			b_626_0 <=( _mesh_17_19_io_out_b_0) ^ ((fiEnable && (4171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1650_0 <=( _mesh_17_19_io_out_c_0) ^ ((fiEnable && (4172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_19_io_in_control_0_shift_b <=( _mesh_17_19_io_out_control_0_shift) ^ ((fiEnable && (4173 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_19_io_in_control_0_dataflow_b <=( _mesh_17_19_io_out_control_0_dataflow) ^ ((fiEnable && (4174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_19_io_in_control_0_propagate_b <=( _mesh_17_19_io_out_control_0_propagate) ^ ((fiEnable && (4175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_19_io_out_valid_0) begin
			b_627_0 <=( _mesh_18_19_io_out_b_0) ^ ((fiEnable && (4176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1651_0 <=( _mesh_18_19_io_out_c_0) ^ ((fiEnable && (4177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_19_io_in_control_0_shift_b <=( _mesh_18_19_io_out_control_0_shift) ^ ((fiEnable && (4178 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_19_io_in_control_0_dataflow_b <=( _mesh_18_19_io_out_control_0_dataflow) ^ ((fiEnable && (4179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_19_io_in_control_0_propagate_b <=( _mesh_18_19_io_out_control_0_propagate) ^ ((fiEnable && (4180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_19_io_out_valid_0) begin
			b_628_0 <=( _mesh_19_19_io_out_b_0) ^ ((fiEnable && (4181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1652_0 <=( _mesh_19_19_io_out_c_0) ^ ((fiEnable && (4182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_19_io_in_control_0_shift_b <=( _mesh_19_19_io_out_control_0_shift) ^ ((fiEnable && (4183 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_19_io_in_control_0_dataflow_b <=( _mesh_19_19_io_out_control_0_dataflow) ^ ((fiEnable && (4184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_19_io_in_control_0_propagate_b <=( _mesh_19_19_io_out_control_0_propagate) ^ ((fiEnable && (4185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_19_io_out_valid_0) begin
			b_629_0 <=( _mesh_20_19_io_out_b_0) ^ ((fiEnable && (4186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1653_0 <=( _mesh_20_19_io_out_c_0) ^ ((fiEnable && (4187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_19_io_in_control_0_shift_b <=( _mesh_20_19_io_out_control_0_shift) ^ ((fiEnable && (4188 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_19_io_in_control_0_dataflow_b <=( _mesh_20_19_io_out_control_0_dataflow) ^ ((fiEnable && (4189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_19_io_in_control_0_propagate_b <=( _mesh_20_19_io_out_control_0_propagate) ^ ((fiEnable && (4190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_19_io_out_valid_0) begin
			b_630_0 <=( _mesh_21_19_io_out_b_0) ^ ((fiEnable && (4191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1654_0 <=( _mesh_21_19_io_out_c_0) ^ ((fiEnable && (4192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_19_io_in_control_0_shift_b <=( _mesh_21_19_io_out_control_0_shift) ^ ((fiEnable && (4193 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_19_io_in_control_0_dataflow_b <=( _mesh_21_19_io_out_control_0_dataflow) ^ ((fiEnable && (4194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_19_io_in_control_0_propagate_b <=( _mesh_21_19_io_out_control_0_propagate) ^ ((fiEnable && (4195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_19_io_out_valid_0) begin
			b_631_0 <=( _mesh_22_19_io_out_b_0) ^ ((fiEnable && (4196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1655_0 <=( _mesh_22_19_io_out_c_0) ^ ((fiEnable && (4197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_19_io_in_control_0_shift_b <=( _mesh_22_19_io_out_control_0_shift) ^ ((fiEnable && (4198 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_19_io_in_control_0_dataflow_b <=( _mesh_22_19_io_out_control_0_dataflow) ^ ((fiEnable && (4199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_19_io_in_control_0_propagate_b <=( _mesh_22_19_io_out_control_0_propagate) ^ ((fiEnable && (4200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_19_io_out_valid_0) begin
			b_632_0 <=( _mesh_23_19_io_out_b_0) ^ ((fiEnable && (4201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1656_0 <=( _mesh_23_19_io_out_c_0) ^ ((fiEnable && (4202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_19_io_in_control_0_shift_b <=( _mesh_23_19_io_out_control_0_shift) ^ ((fiEnable && (4203 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_19_io_in_control_0_dataflow_b <=( _mesh_23_19_io_out_control_0_dataflow) ^ ((fiEnable && (4204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_19_io_in_control_0_propagate_b <=( _mesh_23_19_io_out_control_0_propagate) ^ ((fiEnable && (4205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_19_io_out_valid_0) begin
			b_633_0 <=( _mesh_24_19_io_out_b_0) ^ ((fiEnable && (4206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1657_0 <=( _mesh_24_19_io_out_c_0) ^ ((fiEnable && (4207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_19_io_in_control_0_shift_b <=( _mesh_24_19_io_out_control_0_shift) ^ ((fiEnable && (4208 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_19_io_in_control_0_dataflow_b <=( _mesh_24_19_io_out_control_0_dataflow) ^ ((fiEnable && (4209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_19_io_in_control_0_propagate_b <=( _mesh_24_19_io_out_control_0_propagate) ^ ((fiEnable && (4210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_19_io_out_valid_0) begin
			b_634_0 <=( _mesh_25_19_io_out_b_0) ^ ((fiEnable && (4211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1658_0 <=( _mesh_25_19_io_out_c_0) ^ ((fiEnable && (4212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_19_io_in_control_0_shift_b <=( _mesh_25_19_io_out_control_0_shift) ^ ((fiEnable && (4213 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_19_io_in_control_0_dataflow_b <=( _mesh_25_19_io_out_control_0_dataflow) ^ ((fiEnable && (4214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_19_io_in_control_0_propagate_b <=( _mesh_25_19_io_out_control_0_propagate) ^ ((fiEnable && (4215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_19_io_out_valid_0) begin
			b_635_0 <=( _mesh_26_19_io_out_b_0) ^ ((fiEnable && (4216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1659_0 <=( _mesh_26_19_io_out_c_0) ^ ((fiEnable && (4217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_19_io_in_control_0_shift_b <=( _mesh_26_19_io_out_control_0_shift) ^ ((fiEnable && (4218 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_19_io_in_control_0_dataflow_b <=( _mesh_26_19_io_out_control_0_dataflow) ^ ((fiEnable && (4219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_19_io_in_control_0_propagate_b <=( _mesh_26_19_io_out_control_0_propagate) ^ ((fiEnable && (4220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_19_io_out_valid_0) begin
			b_636_0 <=( _mesh_27_19_io_out_b_0) ^ ((fiEnable && (4221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1660_0 <=( _mesh_27_19_io_out_c_0) ^ ((fiEnable && (4222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_19_io_in_control_0_shift_b <=( _mesh_27_19_io_out_control_0_shift) ^ ((fiEnable && (4223 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_19_io_in_control_0_dataflow_b <=( _mesh_27_19_io_out_control_0_dataflow) ^ ((fiEnable && (4224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_19_io_in_control_0_propagate_b <=( _mesh_27_19_io_out_control_0_propagate) ^ ((fiEnable && (4225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_19_io_out_valid_0) begin
			b_637_0 <=( _mesh_28_19_io_out_b_0) ^ ((fiEnable && (4226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1661_0 <=( _mesh_28_19_io_out_c_0) ^ ((fiEnable && (4227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_19_io_in_control_0_shift_b <=( _mesh_28_19_io_out_control_0_shift) ^ ((fiEnable && (4228 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_19_io_in_control_0_dataflow_b <=( _mesh_28_19_io_out_control_0_dataflow) ^ ((fiEnable && (4229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_19_io_in_control_0_propagate_b <=( _mesh_28_19_io_out_control_0_propagate) ^ ((fiEnable && (4230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_19_io_out_valid_0) begin
			b_638_0 <=( _mesh_29_19_io_out_b_0) ^ ((fiEnable && (4231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1662_0 <=( _mesh_29_19_io_out_c_0) ^ ((fiEnable && (4232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_19_io_in_control_0_shift_b <=( _mesh_29_19_io_out_control_0_shift) ^ ((fiEnable && (4233 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_19_io_in_control_0_dataflow_b <=( _mesh_29_19_io_out_control_0_dataflow) ^ ((fiEnable && (4234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_19_io_in_control_0_propagate_b <=( _mesh_29_19_io_out_control_0_propagate) ^ ((fiEnable && (4235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_19_io_out_valid_0) begin
			b_639_0 <=( _mesh_30_19_io_out_b_0) ^ ((fiEnable && (4236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1663_0 <=( _mesh_30_19_io_out_c_0) ^ ((fiEnable && (4237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_19_io_in_control_0_shift_b <=( _mesh_30_19_io_out_control_0_shift) ^ ((fiEnable && (4238 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_19_io_in_control_0_dataflow_b <=( _mesh_30_19_io_out_control_0_dataflow) ^ ((fiEnable && (4239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_19_io_in_control_0_propagate_b <=( _mesh_30_19_io_out_control_0_propagate) ^ ((fiEnable && (4240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_20_0) begin
			b_640_0 <=( io_in_b_20_0) ^ ((fiEnable && (4241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1664_0 <=( io_in_d_20_0) ^ ((fiEnable && (4242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_20_io_in_control_0_shift_b <=( io_in_control_20_0_shift) ^ ((fiEnable && (4243 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_20_io_in_control_0_dataflow_b <=( io_in_control_20_0_dataflow) ^ ((fiEnable && (4244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_20_io_in_control_0_propagate_b <=( io_in_control_20_0_propagate) ^ ((fiEnable && (4245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_20_io_out_valid_0) begin
			b_641_0 <=( _mesh_0_20_io_out_b_0) ^ ((fiEnable && (4246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1665_0 <=( _mesh_0_20_io_out_c_0) ^ ((fiEnable && (4247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_20_io_in_control_0_shift_b <=( _mesh_0_20_io_out_control_0_shift) ^ ((fiEnable && (4248 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_20_io_in_control_0_dataflow_b <=( _mesh_0_20_io_out_control_0_dataflow) ^ ((fiEnable && (4249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_20_io_in_control_0_propagate_b <=( _mesh_0_20_io_out_control_0_propagate) ^ ((fiEnable && (4250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_20_io_out_valid_0) begin
			b_642_0 <=( _mesh_1_20_io_out_b_0) ^ ((fiEnable && (4251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1666_0 <=( _mesh_1_20_io_out_c_0) ^ ((fiEnable && (4252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_20_io_in_control_0_shift_b <=( _mesh_1_20_io_out_control_0_shift) ^ ((fiEnable && (4253 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_20_io_in_control_0_dataflow_b <=( _mesh_1_20_io_out_control_0_dataflow) ^ ((fiEnable && (4254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_20_io_in_control_0_propagate_b <=( _mesh_1_20_io_out_control_0_propagate) ^ ((fiEnable && (4255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_20_io_out_valid_0) begin
			b_643_0 <=( _mesh_2_20_io_out_b_0) ^ ((fiEnable && (4256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1667_0 <=( _mesh_2_20_io_out_c_0) ^ ((fiEnable && (4257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_20_io_in_control_0_shift_b <=( _mesh_2_20_io_out_control_0_shift) ^ ((fiEnable && (4258 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_20_io_in_control_0_dataflow_b <=( _mesh_2_20_io_out_control_0_dataflow) ^ ((fiEnable && (4259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_20_io_in_control_0_propagate_b <=( _mesh_2_20_io_out_control_0_propagate) ^ ((fiEnable && (4260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_20_io_out_valid_0) begin
			b_644_0 <=( _mesh_3_20_io_out_b_0) ^ ((fiEnable && (4261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1668_0 <=( _mesh_3_20_io_out_c_0) ^ ((fiEnable && (4262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_20_io_in_control_0_shift_b <=( _mesh_3_20_io_out_control_0_shift) ^ ((fiEnable && (4263 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_20_io_in_control_0_dataflow_b <=( _mesh_3_20_io_out_control_0_dataflow) ^ ((fiEnable && (4264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_20_io_in_control_0_propagate_b <=( _mesh_3_20_io_out_control_0_propagate) ^ ((fiEnable && (4265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_20_io_out_valid_0) begin
			b_645_0 <=( _mesh_4_20_io_out_b_0) ^ ((fiEnable && (4266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1669_0 <=( _mesh_4_20_io_out_c_0) ^ ((fiEnable && (4267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_20_io_in_control_0_shift_b <=( _mesh_4_20_io_out_control_0_shift) ^ ((fiEnable && (4268 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_20_io_in_control_0_dataflow_b <=( _mesh_4_20_io_out_control_0_dataflow) ^ ((fiEnable && (4269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_20_io_in_control_0_propagate_b <=( _mesh_4_20_io_out_control_0_propagate) ^ ((fiEnable && (4270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_20_io_out_valid_0) begin
			b_646_0 <=( _mesh_5_20_io_out_b_0) ^ ((fiEnable && (4271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1670_0 <=( _mesh_5_20_io_out_c_0) ^ ((fiEnable && (4272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_20_io_in_control_0_shift_b <=( _mesh_5_20_io_out_control_0_shift) ^ ((fiEnable && (4273 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_20_io_in_control_0_dataflow_b <=( _mesh_5_20_io_out_control_0_dataflow) ^ ((fiEnable && (4274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_20_io_in_control_0_propagate_b <=( _mesh_5_20_io_out_control_0_propagate) ^ ((fiEnable && (4275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_20_io_out_valid_0) begin
			b_647_0 <=( _mesh_6_20_io_out_b_0) ^ ((fiEnable && (4276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1671_0 <=( _mesh_6_20_io_out_c_0) ^ ((fiEnable && (4277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_20_io_in_control_0_shift_b <=( _mesh_6_20_io_out_control_0_shift) ^ ((fiEnable && (4278 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_20_io_in_control_0_dataflow_b <=( _mesh_6_20_io_out_control_0_dataflow) ^ ((fiEnable && (4279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_20_io_in_control_0_propagate_b <=( _mesh_6_20_io_out_control_0_propagate) ^ ((fiEnable && (4280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_20_io_out_valid_0) begin
			b_648_0 <=( _mesh_7_20_io_out_b_0) ^ ((fiEnable && (4281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1672_0 <=( _mesh_7_20_io_out_c_0) ^ ((fiEnable && (4282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_20_io_in_control_0_shift_b <=( _mesh_7_20_io_out_control_0_shift) ^ ((fiEnable && (4283 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_20_io_in_control_0_dataflow_b <=( _mesh_7_20_io_out_control_0_dataflow) ^ ((fiEnable && (4284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_20_io_in_control_0_propagate_b <=( _mesh_7_20_io_out_control_0_propagate) ^ ((fiEnable && (4285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_20_io_out_valid_0) begin
			b_649_0 <=( _mesh_8_20_io_out_b_0) ^ ((fiEnable && (4286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1673_0 <=( _mesh_8_20_io_out_c_0) ^ ((fiEnable && (4287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_20_io_in_control_0_shift_b <=( _mesh_8_20_io_out_control_0_shift) ^ ((fiEnable && (4288 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_20_io_in_control_0_dataflow_b <=( _mesh_8_20_io_out_control_0_dataflow) ^ ((fiEnable && (4289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_20_io_in_control_0_propagate_b <=( _mesh_8_20_io_out_control_0_propagate) ^ ((fiEnable && (4290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_20_io_out_valid_0) begin
			b_650_0 <=( _mesh_9_20_io_out_b_0) ^ ((fiEnable && (4291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1674_0 <=( _mesh_9_20_io_out_c_0) ^ ((fiEnable && (4292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_20_io_in_control_0_shift_b <=( _mesh_9_20_io_out_control_0_shift) ^ ((fiEnable && (4293 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_20_io_in_control_0_dataflow_b <=( _mesh_9_20_io_out_control_0_dataflow) ^ ((fiEnable && (4294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_20_io_in_control_0_propagate_b <=( _mesh_9_20_io_out_control_0_propagate) ^ ((fiEnable && (4295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_20_io_out_valid_0) begin
			b_651_0 <=( _mesh_10_20_io_out_b_0) ^ ((fiEnable && (4296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1675_0 <=( _mesh_10_20_io_out_c_0) ^ ((fiEnable && (4297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_20_io_in_control_0_shift_b <=( _mesh_10_20_io_out_control_0_shift) ^ ((fiEnable && (4298 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_20_io_in_control_0_dataflow_b <=( _mesh_10_20_io_out_control_0_dataflow) ^ ((fiEnable && (4299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_20_io_in_control_0_propagate_b <=( _mesh_10_20_io_out_control_0_propagate) ^ ((fiEnable && (4300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_20_io_out_valid_0) begin
			b_652_0 <=( _mesh_11_20_io_out_b_0) ^ ((fiEnable && (4301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1676_0 <=( _mesh_11_20_io_out_c_0) ^ ((fiEnable && (4302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_20_io_in_control_0_shift_b <=( _mesh_11_20_io_out_control_0_shift) ^ ((fiEnable && (4303 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_20_io_in_control_0_dataflow_b <=( _mesh_11_20_io_out_control_0_dataflow) ^ ((fiEnable && (4304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_20_io_in_control_0_propagate_b <=( _mesh_11_20_io_out_control_0_propagate) ^ ((fiEnable && (4305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_20_io_out_valid_0) begin
			b_653_0 <=( _mesh_12_20_io_out_b_0) ^ ((fiEnable && (4306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1677_0 <=( _mesh_12_20_io_out_c_0) ^ ((fiEnable && (4307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_20_io_in_control_0_shift_b <=( _mesh_12_20_io_out_control_0_shift) ^ ((fiEnable && (4308 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_20_io_in_control_0_dataflow_b <=( _mesh_12_20_io_out_control_0_dataflow) ^ ((fiEnable && (4309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_20_io_in_control_0_propagate_b <=( _mesh_12_20_io_out_control_0_propagate) ^ ((fiEnable && (4310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_20_io_out_valid_0) begin
			b_654_0 <=( _mesh_13_20_io_out_b_0) ^ ((fiEnable && (4311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1678_0 <=( _mesh_13_20_io_out_c_0) ^ ((fiEnable && (4312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_20_io_in_control_0_shift_b <=( _mesh_13_20_io_out_control_0_shift) ^ ((fiEnable && (4313 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_20_io_in_control_0_dataflow_b <=( _mesh_13_20_io_out_control_0_dataflow) ^ ((fiEnable && (4314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_20_io_in_control_0_propagate_b <=( _mesh_13_20_io_out_control_0_propagate) ^ ((fiEnable && (4315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_20_io_out_valid_0) begin
			b_655_0 <=( _mesh_14_20_io_out_b_0) ^ ((fiEnable && (4316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1679_0 <=( _mesh_14_20_io_out_c_0) ^ ((fiEnable && (4317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_20_io_in_control_0_shift_b <=( _mesh_14_20_io_out_control_0_shift) ^ ((fiEnable && (4318 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_20_io_in_control_0_dataflow_b <=( _mesh_14_20_io_out_control_0_dataflow) ^ ((fiEnable && (4319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_20_io_in_control_0_propagate_b <=( _mesh_14_20_io_out_control_0_propagate) ^ ((fiEnable && (4320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_20_io_out_valid_0) begin
			b_656_0 <=( _mesh_15_20_io_out_b_0) ^ ((fiEnable && (4321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1680_0 <=( _mesh_15_20_io_out_c_0) ^ ((fiEnable && (4322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_20_io_in_control_0_shift_b <=( _mesh_15_20_io_out_control_0_shift) ^ ((fiEnable && (4323 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_20_io_in_control_0_dataflow_b <=( _mesh_15_20_io_out_control_0_dataflow) ^ ((fiEnable && (4324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_20_io_in_control_0_propagate_b <=( _mesh_15_20_io_out_control_0_propagate) ^ ((fiEnable && (4325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_20_io_out_valid_0) begin
			b_657_0 <=( _mesh_16_20_io_out_b_0) ^ ((fiEnable && (4326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1681_0 <=( _mesh_16_20_io_out_c_0) ^ ((fiEnable && (4327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_20_io_in_control_0_shift_b <=( _mesh_16_20_io_out_control_0_shift) ^ ((fiEnable && (4328 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_20_io_in_control_0_dataflow_b <=( _mesh_16_20_io_out_control_0_dataflow) ^ ((fiEnable && (4329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_20_io_in_control_0_propagate_b <=( _mesh_16_20_io_out_control_0_propagate) ^ ((fiEnable && (4330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_20_io_out_valid_0) begin
			b_658_0 <=( _mesh_17_20_io_out_b_0) ^ ((fiEnable && (4331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1682_0 <=( _mesh_17_20_io_out_c_0) ^ ((fiEnable && (4332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_20_io_in_control_0_shift_b <=( _mesh_17_20_io_out_control_0_shift) ^ ((fiEnable && (4333 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_20_io_in_control_0_dataflow_b <=( _mesh_17_20_io_out_control_0_dataflow) ^ ((fiEnable && (4334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_20_io_in_control_0_propagate_b <=( _mesh_17_20_io_out_control_0_propagate) ^ ((fiEnable && (4335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_20_io_out_valid_0) begin
			b_659_0 <=( _mesh_18_20_io_out_b_0) ^ ((fiEnable && (4336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1683_0 <=( _mesh_18_20_io_out_c_0) ^ ((fiEnable && (4337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_20_io_in_control_0_shift_b <=( _mesh_18_20_io_out_control_0_shift) ^ ((fiEnable && (4338 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_20_io_in_control_0_dataflow_b <=( _mesh_18_20_io_out_control_0_dataflow) ^ ((fiEnable && (4339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_20_io_in_control_0_propagate_b <=( _mesh_18_20_io_out_control_0_propagate) ^ ((fiEnable && (4340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_20_io_out_valid_0) begin
			b_660_0 <=( _mesh_19_20_io_out_b_0) ^ ((fiEnable && (4341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1684_0 <=( _mesh_19_20_io_out_c_0) ^ ((fiEnable && (4342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_20_io_in_control_0_shift_b <=( _mesh_19_20_io_out_control_0_shift) ^ ((fiEnable && (4343 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_20_io_in_control_0_dataflow_b <=( _mesh_19_20_io_out_control_0_dataflow) ^ ((fiEnable && (4344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_20_io_in_control_0_propagate_b <=( _mesh_19_20_io_out_control_0_propagate) ^ ((fiEnable && (4345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_20_io_out_valid_0) begin
			b_661_0 <=( _mesh_20_20_io_out_b_0) ^ ((fiEnable && (4346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1685_0 <=( _mesh_20_20_io_out_c_0) ^ ((fiEnable && (4347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_20_io_in_control_0_shift_b <=( _mesh_20_20_io_out_control_0_shift) ^ ((fiEnable && (4348 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_20_io_in_control_0_dataflow_b <=( _mesh_20_20_io_out_control_0_dataflow) ^ ((fiEnable && (4349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_20_io_in_control_0_propagate_b <=( _mesh_20_20_io_out_control_0_propagate) ^ ((fiEnable && (4350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_20_io_out_valid_0) begin
			b_662_0 <=( _mesh_21_20_io_out_b_0) ^ ((fiEnable && (4351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1686_0 <=( _mesh_21_20_io_out_c_0) ^ ((fiEnable && (4352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_20_io_in_control_0_shift_b <=( _mesh_21_20_io_out_control_0_shift) ^ ((fiEnable && (4353 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_20_io_in_control_0_dataflow_b <=( _mesh_21_20_io_out_control_0_dataflow) ^ ((fiEnable && (4354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_20_io_in_control_0_propagate_b <=( _mesh_21_20_io_out_control_0_propagate) ^ ((fiEnable && (4355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_20_io_out_valid_0) begin
			b_663_0 <=( _mesh_22_20_io_out_b_0) ^ ((fiEnable && (4356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1687_0 <=( _mesh_22_20_io_out_c_0) ^ ((fiEnable && (4357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_20_io_in_control_0_shift_b <=( _mesh_22_20_io_out_control_0_shift) ^ ((fiEnable && (4358 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_20_io_in_control_0_dataflow_b <=( _mesh_22_20_io_out_control_0_dataflow) ^ ((fiEnable && (4359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_20_io_in_control_0_propagate_b <=( _mesh_22_20_io_out_control_0_propagate) ^ ((fiEnable && (4360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_20_io_out_valid_0) begin
			b_664_0 <=( _mesh_23_20_io_out_b_0) ^ ((fiEnable && (4361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1688_0 <=( _mesh_23_20_io_out_c_0) ^ ((fiEnable && (4362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_20_io_in_control_0_shift_b <=( _mesh_23_20_io_out_control_0_shift) ^ ((fiEnable && (4363 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_20_io_in_control_0_dataflow_b <=( _mesh_23_20_io_out_control_0_dataflow) ^ ((fiEnable && (4364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_20_io_in_control_0_propagate_b <=( _mesh_23_20_io_out_control_0_propagate) ^ ((fiEnable && (4365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_20_io_out_valid_0) begin
			b_665_0 <=( _mesh_24_20_io_out_b_0) ^ ((fiEnable && (4366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1689_0 <=( _mesh_24_20_io_out_c_0) ^ ((fiEnable && (4367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_20_io_in_control_0_shift_b <=( _mesh_24_20_io_out_control_0_shift) ^ ((fiEnable && (4368 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_20_io_in_control_0_dataflow_b <=( _mesh_24_20_io_out_control_0_dataflow) ^ ((fiEnable && (4369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_20_io_in_control_0_propagate_b <=( _mesh_24_20_io_out_control_0_propagate) ^ ((fiEnable && (4370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_20_io_out_valid_0) begin
			b_666_0 <=( _mesh_25_20_io_out_b_0) ^ ((fiEnable && (4371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1690_0 <=( _mesh_25_20_io_out_c_0) ^ ((fiEnable && (4372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_20_io_in_control_0_shift_b <=( _mesh_25_20_io_out_control_0_shift) ^ ((fiEnable && (4373 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_20_io_in_control_0_dataflow_b <=( _mesh_25_20_io_out_control_0_dataflow) ^ ((fiEnable && (4374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_20_io_in_control_0_propagate_b <=( _mesh_25_20_io_out_control_0_propagate) ^ ((fiEnable && (4375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_20_io_out_valid_0) begin
			b_667_0 <=( _mesh_26_20_io_out_b_0) ^ ((fiEnable && (4376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1691_0 <=( _mesh_26_20_io_out_c_0) ^ ((fiEnable && (4377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_20_io_in_control_0_shift_b <=( _mesh_26_20_io_out_control_0_shift) ^ ((fiEnable && (4378 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_20_io_in_control_0_dataflow_b <=( _mesh_26_20_io_out_control_0_dataflow) ^ ((fiEnable && (4379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_20_io_in_control_0_propagate_b <=( _mesh_26_20_io_out_control_0_propagate) ^ ((fiEnable && (4380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_20_io_out_valid_0) begin
			b_668_0 <=( _mesh_27_20_io_out_b_0) ^ ((fiEnable && (4381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1692_0 <=( _mesh_27_20_io_out_c_0) ^ ((fiEnable && (4382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_20_io_in_control_0_shift_b <=( _mesh_27_20_io_out_control_0_shift) ^ ((fiEnable && (4383 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_20_io_in_control_0_dataflow_b <=( _mesh_27_20_io_out_control_0_dataflow) ^ ((fiEnable && (4384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_20_io_in_control_0_propagate_b <=( _mesh_27_20_io_out_control_0_propagate) ^ ((fiEnable && (4385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_20_io_out_valid_0) begin
			b_669_0 <=( _mesh_28_20_io_out_b_0) ^ ((fiEnable && (4386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1693_0 <=( _mesh_28_20_io_out_c_0) ^ ((fiEnable && (4387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_20_io_in_control_0_shift_b <=( _mesh_28_20_io_out_control_0_shift) ^ ((fiEnable && (4388 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_20_io_in_control_0_dataflow_b <=( _mesh_28_20_io_out_control_0_dataflow) ^ ((fiEnable && (4389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_20_io_in_control_0_propagate_b <=( _mesh_28_20_io_out_control_0_propagate) ^ ((fiEnable && (4390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_20_io_out_valid_0) begin
			b_670_0 <=( _mesh_29_20_io_out_b_0) ^ ((fiEnable && (4391 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1694_0 <=( _mesh_29_20_io_out_c_0) ^ ((fiEnable && (4392 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_20_io_in_control_0_shift_b <=( _mesh_29_20_io_out_control_0_shift) ^ ((fiEnable && (4393 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_20_io_in_control_0_dataflow_b <=( _mesh_29_20_io_out_control_0_dataflow) ^ ((fiEnable && (4394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_20_io_in_control_0_propagate_b <=( _mesh_29_20_io_out_control_0_propagate) ^ ((fiEnable && (4395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_20_io_out_valid_0) begin
			b_671_0 <=( _mesh_30_20_io_out_b_0) ^ ((fiEnable && (4396 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1695_0 <=( _mesh_30_20_io_out_c_0) ^ ((fiEnable && (4397 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_20_io_in_control_0_shift_b <=( _mesh_30_20_io_out_control_0_shift) ^ ((fiEnable && (4398 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_20_io_in_control_0_dataflow_b <=( _mesh_30_20_io_out_control_0_dataflow) ^ ((fiEnable && (4399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_20_io_in_control_0_propagate_b <=( _mesh_30_20_io_out_control_0_propagate) ^ ((fiEnable && (4400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_21_0) begin
			b_672_0 <=( io_in_b_21_0) ^ ((fiEnable && (4401 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1696_0 <=( io_in_d_21_0) ^ ((fiEnable && (4402 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_21_io_in_control_0_shift_b <=( io_in_control_21_0_shift) ^ ((fiEnable && (4403 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_21_io_in_control_0_dataflow_b <=( io_in_control_21_0_dataflow) ^ ((fiEnable && (4404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_21_io_in_control_0_propagate_b <=( io_in_control_21_0_propagate) ^ ((fiEnable && (4405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_21_io_out_valid_0) begin
			b_673_0 <=( _mesh_0_21_io_out_b_0) ^ ((fiEnable && (4406 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1697_0 <=( _mesh_0_21_io_out_c_0) ^ ((fiEnable && (4407 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_21_io_in_control_0_shift_b <=( _mesh_0_21_io_out_control_0_shift) ^ ((fiEnable && (4408 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_21_io_in_control_0_dataflow_b <=( _mesh_0_21_io_out_control_0_dataflow) ^ ((fiEnable && (4409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_21_io_in_control_0_propagate_b <=( _mesh_0_21_io_out_control_0_propagate) ^ ((fiEnable && (4410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_21_io_out_valid_0) begin
			b_674_0 <=( _mesh_1_21_io_out_b_0) ^ ((fiEnable && (4411 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1698_0 <=( _mesh_1_21_io_out_c_0) ^ ((fiEnable && (4412 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_21_io_in_control_0_shift_b <=( _mesh_1_21_io_out_control_0_shift) ^ ((fiEnable && (4413 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_21_io_in_control_0_dataflow_b <=( _mesh_1_21_io_out_control_0_dataflow) ^ ((fiEnable && (4414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_21_io_in_control_0_propagate_b <=( _mesh_1_21_io_out_control_0_propagate) ^ ((fiEnable && (4415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_21_io_out_valid_0) begin
			b_675_0 <=( _mesh_2_21_io_out_b_0) ^ ((fiEnable && (4416 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1699_0 <=( _mesh_2_21_io_out_c_0) ^ ((fiEnable && (4417 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_21_io_in_control_0_shift_b <=( _mesh_2_21_io_out_control_0_shift) ^ ((fiEnable && (4418 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_21_io_in_control_0_dataflow_b <=( _mesh_2_21_io_out_control_0_dataflow) ^ ((fiEnable && (4419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_21_io_in_control_0_propagate_b <=( _mesh_2_21_io_out_control_0_propagate) ^ ((fiEnable && (4420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_21_io_out_valid_0) begin
			b_676_0 <=( _mesh_3_21_io_out_b_0) ^ ((fiEnable && (4421 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1700_0 <=( _mesh_3_21_io_out_c_0) ^ ((fiEnable && (4422 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_21_io_in_control_0_shift_b <=( _mesh_3_21_io_out_control_0_shift) ^ ((fiEnable && (4423 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_21_io_in_control_0_dataflow_b <=( _mesh_3_21_io_out_control_0_dataflow) ^ ((fiEnable && (4424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_21_io_in_control_0_propagate_b <=( _mesh_3_21_io_out_control_0_propagate) ^ ((fiEnable && (4425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_21_io_out_valid_0) begin
			b_677_0 <=( _mesh_4_21_io_out_b_0) ^ ((fiEnable && (4426 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1701_0 <=( _mesh_4_21_io_out_c_0) ^ ((fiEnable && (4427 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_21_io_in_control_0_shift_b <=( _mesh_4_21_io_out_control_0_shift) ^ ((fiEnable && (4428 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_21_io_in_control_0_dataflow_b <=( _mesh_4_21_io_out_control_0_dataflow) ^ ((fiEnable && (4429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_21_io_in_control_0_propagate_b <=( _mesh_4_21_io_out_control_0_propagate) ^ ((fiEnable && (4430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_21_io_out_valid_0) begin
			b_678_0 <=( _mesh_5_21_io_out_b_0) ^ ((fiEnable && (4431 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1702_0 <=( _mesh_5_21_io_out_c_0) ^ ((fiEnable && (4432 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_21_io_in_control_0_shift_b <=( _mesh_5_21_io_out_control_0_shift) ^ ((fiEnable && (4433 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_21_io_in_control_0_dataflow_b <=( _mesh_5_21_io_out_control_0_dataflow) ^ ((fiEnable && (4434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_21_io_in_control_0_propagate_b <=( _mesh_5_21_io_out_control_0_propagate) ^ ((fiEnable && (4435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_21_io_out_valid_0) begin
			b_679_0 <=( _mesh_6_21_io_out_b_0) ^ ((fiEnable && (4436 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1703_0 <=( _mesh_6_21_io_out_c_0) ^ ((fiEnable && (4437 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_21_io_in_control_0_shift_b <=( _mesh_6_21_io_out_control_0_shift) ^ ((fiEnable && (4438 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_21_io_in_control_0_dataflow_b <=( _mesh_6_21_io_out_control_0_dataflow) ^ ((fiEnable && (4439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_21_io_in_control_0_propagate_b <=( _mesh_6_21_io_out_control_0_propagate) ^ ((fiEnable && (4440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_21_io_out_valid_0) begin
			b_680_0 <=( _mesh_7_21_io_out_b_0) ^ ((fiEnable && (4441 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1704_0 <=( _mesh_7_21_io_out_c_0) ^ ((fiEnable && (4442 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_21_io_in_control_0_shift_b <=( _mesh_7_21_io_out_control_0_shift) ^ ((fiEnable && (4443 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_21_io_in_control_0_dataflow_b <=( _mesh_7_21_io_out_control_0_dataflow) ^ ((fiEnable && (4444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_21_io_in_control_0_propagate_b <=( _mesh_7_21_io_out_control_0_propagate) ^ ((fiEnable && (4445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_21_io_out_valid_0) begin
			b_681_0 <=( _mesh_8_21_io_out_b_0) ^ ((fiEnable && (4446 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1705_0 <=( _mesh_8_21_io_out_c_0) ^ ((fiEnable && (4447 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_21_io_in_control_0_shift_b <=( _mesh_8_21_io_out_control_0_shift) ^ ((fiEnable && (4448 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_21_io_in_control_0_dataflow_b <=( _mesh_8_21_io_out_control_0_dataflow) ^ ((fiEnable && (4449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_21_io_in_control_0_propagate_b <=( _mesh_8_21_io_out_control_0_propagate) ^ ((fiEnable && (4450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_21_io_out_valid_0) begin
			b_682_0 <=( _mesh_9_21_io_out_b_0) ^ ((fiEnable && (4451 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1706_0 <=( _mesh_9_21_io_out_c_0) ^ ((fiEnable && (4452 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_21_io_in_control_0_shift_b <=( _mesh_9_21_io_out_control_0_shift) ^ ((fiEnable && (4453 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_21_io_in_control_0_dataflow_b <=( _mesh_9_21_io_out_control_0_dataflow) ^ ((fiEnable && (4454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_21_io_in_control_0_propagate_b <=( _mesh_9_21_io_out_control_0_propagate) ^ ((fiEnable && (4455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_21_io_out_valid_0) begin
			b_683_0 <=( _mesh_10_21_io_out_b_0) ^ ((fiEnable && (4456 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1707_0 <=( _mesh_10_21_io_out_c_0) ^ ((fiEnable && (4457 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_21_io_in_control_0_shift_b <=( _mesh_10_21_io_out_control_0_shift) ^ ((fiEnable && (4458 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_21_io_in_control_0_dataflow_b <=( _mesh_10_21_io_out_control_0_dataflow) ^ ((fiEnable && (4459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_21_io_in_control_0_propagate_b <=( _mesh_10_21_io_out_control_0_propagate) ^ ((fiEnable && (4460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_21_io_out_valid_0) begin
			b_684_0 <=( _mesh_11_21_io_out_b_0) ^ ((fiEnable && (4461 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1708_0 <=( _mesh_11_21_io_out_c_0) ^ ((fiEnable && (4462 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_21_io_in_control_0_shift_b <=( _mesh_11_21_io_out_control_0_shift) ^ ((fiEnable && (4463 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_21_io_in_control_0_dataflow_b <=( _mesh_11_21_io_out_control_0_dataflow) ^ ((fiEnable && (4464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_21_io_in_control_0_propagate_b <=( _mesh_11_21_io_out_control_0_propagate) ^ ((fiEnable && (4465 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_21_io_out_valid_0) begin
			b_685_0 <=( _mesh_12_21_io_out_b_0) ^ ((fiEnable && (4466 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1709_0 <=( _mesh_12_21_io_out_c_0) ^ ((fiEnable && (4467 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_21_io_in_control_0_shift_b <=( _mesh_12_21_io_out_control_0_shift) ^ ((fiEnable && (4468 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_21_io_in_control_0_dataflow_b <=( _mesh_12_21_io_out_control_0_dataflow) ^ ((fiEnable && (4469 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_21_io_in_control_0_propagate_b <=( _mesh_12_21_io_out_control_0_propagate) ^ ((fiEnable && (4470 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_21_io_out_valid_0) begin
			b_686_0 <=( _mesh_13_21_io_out_b_0) ^ ((fiEnable && (4471 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1710_0 <=( _mesh_13_21_io_out_c_0) ^ ((fiEnable && (4472 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_21_io_in_control_0_shift_b <=( _mesh_13_21_io_out_control_0_shift) ^ ((fiEnable && (4473 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_21_io_in_control_0_dataflow_b <=( _mesh_13_21_io_out_control_0_dataflow) ^ ((fiEnable && (4474 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_21_io_in_control_0_propagate_b <=( _mesh_13_21_io_out_control_0_propagate) ^ ((fiEnable && (4475 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_21_io_out_valid_0) begin
			b_687_0 <=( _mesh_14_21_io_out_b_0) ^ ((fiEnable && (4476 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1711_0 <=( _mesh_14_21_io_out_c_0) ^ ((fiEnable && (4477 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_21_io_in_control_0_shift_b <=( _mesh_14_21_io_out_control_0_shift) ^ ((fiEnable && (4478 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_21_io_in_control_0_dataflow_b <=( _mesh_14_21_io_out_control_0_dataflow) ^ ((fiEnable && (4479 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_21_io_in_control_0_propagate_b <=( _mesh_14_21_io_out_control_0_propagate) ^ ((fiEnable && (4480 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_21_io_out_valid_0) begin
			b_688_0 <=( _mesh_15_21_io_out_b_0) ^ ((fiEnable && (4481 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1712_0 <=( _mesh_15_21_io_out_c_0) ^ ((fiEnable && (4482 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_21_io_in_control_0_shift_b <=( _mesh_15_21_io_out_control_0_shift) ^ ((fiEnable && (4483 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_21_io_in_control_0_dataflow_b <=( _mesh_15_21_io_out_control_0_dataflow) ^ ((fiEnable && (4484 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_21_io_in_control_0_propagate_b <=( _mesh_15_21_io_out_control_0_propagate) ^ ((fiEnable && (4485 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_21_io_out_valid_0) begin
			b_689_0 <=( _mesh_16_21_io_out_b_0) ^ ((fiEnable && (4486 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1713_0 <=( _mesh_16_21_io_out_c_0) ^ ((fiEnable && (4487 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_21_io_in_control_0_shift_b <=( _mesh_16_21_io_out_control_0_shift) ^ ((fiEnable && (4488 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_21_io_in_control_0_dataflow_b <=( _mesh_16_21_io_out_control_0_dataflow) ^ ((fiEnable && (4489 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_21_io_in_control_0_propagate_b <=( _mesh_16_21_io_out_control_0_propagate) ^ ((fiEnable && (4490 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_21_io_out_valid_0) begin
			b_690_0 <=( _mesh_17_21_io_out_b_0) ^ ((fiEnable && (4491 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1714_0 <=( _mesh_17_21_io_out_c_0) ^ ((fiEnable && (4492 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_21_io_in_control_0_shift_b <=( _mesh_17_21_io_out_control_0_shift) ^ ((fiEnable && (4493 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_21_io_in_control_0_dataflow_b <=( _mesh_17_21_io_out_control_0_dataflow) ^ ((fiEnable && (4494 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_21_io_in_control_0_propagate_b <=( _mesh_17_21_io_out_control_0_propagate) ^ ((fiEnable && (4495 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_21_io_out_valid_0) begin
			b_691_0 <=( _mesh_18_21_io_out_b_0) ^ ((fiEnable && (4496 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1715_0 <=( _mesh_18_21_io_out_c_0) ^ ((fiEnable && (4497 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_21_io_in_control_0_shift_b <=( _mesh_18_21_io_out_control_0_shift) ^ ((fiEnable && (4498 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_21_io_in_control_0_dataflow_b <=( _mesh_18_21_io_out_control_0_dataflow) ^ ((fiEnable && (4499 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_21_io_in_control_0_propagate_b <=( _mesh_18_21_io_out_control_0_propagate) ^ ((fiEnable && (4500 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_21_io_out_valid_0) begin
			b_692_0 <=( _mesh_19_21_io_out_b_0) ^ ((fiEnable && (4501 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1716_0 <=( _mesh_19_21_io_out_c_0) ^ ((fiEnable && (4502 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_21_io_in_control_0_shift_b <=( _mesh_19_21_io_out_control_0_shift) ^ ((fiEnable && (4503 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_21_io_in_control_0_dataflow_b <=( _mesh_19_21_io_out_control_0_dataflow) ^ ((fiEnable && (4504 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_21_io_in_control_0_propagate_b <=( _mesh_19_21_io_out_control_0_propagate) ^ ((fiEnable && (4505 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_21_io_out_valid_0) begin
			b_693_0 <=( _mesh_20_21_io_out_b_0) ^ ((fiEnable && (4506 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1717_0 <=( _mesh_20_21_io_out_c_0) ^ ((fiEnable && (4507 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_21_io_in_control_0_shift_b <=( _mesh_20_21_io_out_control_0_shift) ^ ((fiEnable && (4508 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_21_io_in_control_0_dataflow_b <=( _mesh_20_21_io_out_control_0_dataflow) ^ ((fiEnable && (4509 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_21_io_in_control_0_propagate_b <=( _mesh_20_21_io_out_control_0_propagate) ^ ((fiEnable && (4510 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_21_io_out_valid_0) begin
			b_694_0 <=( _mesh_21_21_io_out_b_0) ^ ((fiEnable && (4511 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1718_0 <=( _mesh_21_21_io_out_c_0) ^ ((fiEnable && (4512 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_21_io_in_control_0_shift_b <=( _mesh_21_21_io_out_control_0_shift) ^ ((fiEnable && (4513 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_21_io_in_control_0_dataflow_b <=( _mesh_21_21_io_out_control_0_dataflow) ^ ((fiEnable && (4514 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_21_io_in_control_0_propagate_b <=( _mesh_21_21_io_out_control_0_propagate) ^ ((fiEnable && (4515 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_21_io_out_valid_0) begin
			b_695_0 <=( _mesh_22_21_io_out_b_0) ^ ((fiEnable && (4516 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1719_0 <=( _mesh_22_21_io_out_c_0) ^ ((fiEnable && (4517 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_21_io_in_control_0_shift_b <=( _mesh_22_21_io_out_control_0_shift) ^ ((fiEnable && (4518 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_21_io_in_control_0_dataflow_b <=( _mesh_22_21_io_out_control_0_dataflow) ^ ((fiEnable && (4519 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_21_io_in_control_0_propagate_b <=( _mesh_22_21_io_out_control_0_propagate) ^ ((fiEnable && (4520 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_21_io_out_valid_0) begin
			b_696_0 <=( _mesh_23_21_io_out_b_0) ^ ((fiEnable && (4521 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1720_0 <=( _mesh_23_21_io_out_c_0) ^ ((fiEnable && (4522 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_21_io_in_control_0_shift_b <=( _mesh_23_21_io_out_control_0_shift) ^ ((fiEnable && (4523 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_21_io_in_control_0_dataflow_b <=( _mesh_23_21_io_out_control_0_dataflow) ^ ((fiEnable && (4524 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_21_io_in_control_0_propagate_b <=( _mesh_23_21_io_out_control_0_propagate) ^ ((fiEnable && (4525 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_21_io_out_valid_0) begin
			b_697_0 <=( _mesh_24_21_io_out_b_0) ^ ((fiEnable && (4526 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1721_0 <=( _mesh_24_21_io_out_c_0) ^ ((fiEnable && (4527 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_21_io_in_control_0_shift_b <=( _mesh_24_21_io_out_control_0_shift) ^ ((fiEnable && (4528 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_21_io_in_control_0_dataflow_b <=( _mesh_24_21_io_out_control_0_dataflow) ^ ((fiEnable && (4529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_21_io_in_control_0_propagate_b <=( _mesh_24_21_io_out_control_0_propagate) ^ ((fiEnable && (4530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_21_io_out_valid_0) begin
			b_698_0 <=( _mesh_25_21_io_out_b_0) ^ ((fiEnable && (4531 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1722_0 <=( _mesh_25_21_io_out_c_0) ^ ((fiEnable && (4532 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_21_io_in_control_0_shift_b <=( _mesh_25_21_io_out_control_0_shift) ^ ((fiEnable && (4533 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_21_io_in_control_0_dataflow_b <=( _mesh_25_21_io_out_control_0_dataflow) ^ ((fiEnable && (4534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_21_io_in_control_0_propagate_b <=( _mesh_25_21_io_out_control_0_propagate) ^ ((fiEnable && (4535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_21_io_out_valid_0) begin
			b_699_0 <=( _mesh_26_21_io_out_b_0) ^ ((fiEnable && (4536 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1723_0 <=( _mesh_26_21_io_out_c_0) ^ ((fiEnable && (4537 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_21_io_in_control_0_shift_b <=( _mesh_26_21_io_out_control_0_shift) ^ ((fiEnable && (4538 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_21_io_in_control_0_dataflow_b <=( _mesh_26_21_io_out_control_0_dataflow) ^ ((fiEnable && (4539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_21_io_in_control_0_propagate_b <=( _mesh_26_21_io_out_control_0_propagate) ^ ((fiEnable && (4540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_21_io_out_valid_0) begin
			b_700_0 <=( _mesh_27_21_io_out_b_0) ^ ((fiEnable && (4541 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1724_0 <=( _mesh_27_21_io_out_c_0) ^ ((fiEnable && (4542 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_21_io_in_control_0_shift_b <=( _mesh_27_21_io_out_control_0_shift) ^ ((fiEnable && (4543 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_21_io_in_control_0_dataflow_b <=( _mesh_27_21_io_out_control_0_dataflow) ^ ((fiEnable && (4544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_21_io_in_control_0_propagate_b <=( _mesh_27_21_io_out_control_0_propagate) ^ ((fiEnable && (4545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_21_io_out_valid_0) begin
			b_701_0 <=( _mesh_28_21_io_out_b_0) ^ ((fiEnable && (4546 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1725_0 <=( _mesh_28_21_io_out_c_0) ^ ((fiEnable && (4547 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_21_io_in_control_0_shift_b <=( _mesh_28_21_io_out_control_0_shift) ^ ((fiEnable && (4548 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_21_io_in_control_0_dataflow_b <=( _mesh_28_21_io_out_control_0_dataflow) ^ ((fiEnable && (4549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_21_io_in_control_0_propagate_b <=( _mesh_28_21_io_out_control_0_propagate) ^ ((fiEnable && (4550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_21_io_out_valid_0) begin
			b_702_0 <=( _mesh_29_21_io_out_b_0) ^ ((fiEnable && (4551 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1726_0 <=( _mesh_29_21_io_out_c_0) ^ ((fiEnable && (4552 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_21_io_in_control_0_shift_b <=( _mesh_29_21_io_out_control_0_shift) ^ ((fiEnable && (4553 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_21_io_in_control_0_dataflow_b <=( _mesh_29_21_io_out_control_0_dataflow) ^ ((fiEnable && (4554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_21_io_in_control_0_propagate_b <=( _mesh_29_21_io_out_control_0_propagate) ^ ((fiEnable && (4555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_21_io_out_valid_0) begin
			b_703_0 <=( _mesh_30_21_io_out_b_0) ^ ((fiEnable && (4556 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1727_0 <=( _mesh_30_21_io_out_c_0) ^ ((fiEnable && (4557 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_21_io_in_control_0_shift_b <=( _mesh_30_21_io_out_control_0_shift) ^ ((fiEnable && (4558 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_21_io_in_control_0_dataflow_b <=( _mesh_30_21_io_out_control_0_dataflow) ^ ((fiEnable && (4559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_21_io_in_control_0_propagate_b <=( _mesh_30_21_io_out_control_0_propagate) ^ ((fiEnable && (4560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_22_0) begin
			b_704_0 <=( io_in_b_22_0) ^ ((fiEnable && (4561 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1728_0 <=( io_in_d_22_0) ^ ((fiEnable && (4562 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_22_io_in_control_0_shift_b <=( io_in_control_22_0_shift) ^ ((fiEnable && (4563 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_22_io_in_control_0_dataflow_b <=( io_in_control_22_0_dataflow) ^ ((fiEnable && (4564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_22_io_in_control_0_propagate_b <=( io_in_control_22_0_propagate) ^ ((fiEnable && (4565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_22_io_out_valid_0) begin
			b_705_0 <=( _mesh_0_22_io_out_b_0) ^ ((fiEnable && (4566 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1729_0 <=( _mesh_0_22_io_out_c_0) ^ ((fiEnable && (4567 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_22_io_in_control_0_shift_b <=( _mesh_0_22_io_out_control_0_shift) ^ ((fiEnable && (4568 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_22_io_in_control_0_dataflow_b <=( _mesh_0_22_io_out_control_0_dataflow) ^ ((fiEnable && (4569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_22_io_in_control_0_propagate_b <=( _mesh_0_22_io_out_control_0_propagate) ^ ((fiEnable && (4570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_22_io_out_valid_0) begin
			b_706_0 <=( _mesh_1_22_io_out_b_0) ^ ((fiEnable && (4571 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1730_0 <=( _mesh_1_22_io_out_c_0) ^ ((fiEnable && (4572 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_22_io_in_control_0_shift_b <=( _mesh_1_22_io_out_control_0_shift) ^ ((fiEnable && (4573 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_22_io_in_control_0_dataflow_b <=( _mesh_1_22_io_out_control_0_dataflow) ^ ((fiEnable && (4574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_22_io_in_control_0_propagate_b <=( _mesh_1_22_io_out_control_0_propagate) ^ ((fiEnable && (4575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_22_io_out_valid_0) begin
			b_707_0 <=( _mesh_2_22_io_out_b_0) ^ ((fiEnable && (4576 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1731_0 <=( _mesh_2_22_io_out_c_0) ^ ((fiEnable && (4577 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_22_io_in_control_0_shift_b <=( _mesh_2_22_io_out_control_0_shift) ^ ((fiEnable && (4578 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_22_io_in_control_0_dataflow_b <=( _mesh_2_22_io_out_control_0_dataflow) ^ ((fiEnable && (4579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_22_io_in_control_0_propagate_b <=( _mesh_2_22_io_out_control_0_propagate) ^ ((fiEnable && (4580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_22_io_out_valid_0) begin
			b_708_0 <=( _mesh_3_22_io_out_b_0) ^ ((fiEnable && (4581 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1732_0 <=( _mesh_3_22_io_out_c_0) ^ ((fiEnable && (4582 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_22_io_in_control_0_shift_b <=( _mesh_3_22_io_out_control_0_shift) ^ ((fiEnable && (4583 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_22_io_in_control_0_dataflow_b <=( _mesh_3_22_io_out_control_0_dataflow) ^ ((fiEnable && (4584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_22_io_in_control_0_propagate_b <=( _mesh_3_22_io_out_control_0_propagate) ^ ((fiEnable && (4585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_22_io_out_valid_0) begin
			b_709_0 <=( _mesh_4_22_io_out_b_0) ^ ((fiEnable && (4586 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1733_0 <=( _mesh_4_22_io_out_c_0) ^ ((fiEnable && (4587 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_22_io_in_control_0_shift_b <=( _mesh_4_22_io_out_control_0_shift) ^ ((fiEnable && (4588 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_22_io_in_control_0_dataflow_b <=( _mesh_4_22_io_out_control_0_dataflow) ^ ((fiEnable && (4589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_22_io_in_control_0_propagate_b <=( _mesh_4_22_io_out_control_0_propagate) ^ ((fiEnable && (4590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_22_io_out_valid_0) begin
			b_710_0 <=( _mesh_5_22_io_out_b_0) ^ ((fiEnable && (4591 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1734_0 <=( _mesh_5_22_io_out_c_0) ^ ((fiEnable && (4592 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_22_io_in_control_0_shift_b <=( _mesh_5_22_io_out_control_0_shift) ^ ((fiEnable && (4593 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_22_io_in_control_0_dataflow_b <=( _mesh_5_22_io_out_control_0_dataflow) ^ ((fiEnable && (4594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_22_io_in_control_0_propagate_b <=( _mesh_5_22_io_out_control_0_propagate) ^ ((fiEnable && (4595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_22_io_out_valid_0) begin
			b_711_0 <=( _mesh_6_22_io_out_b_0) ^ ((fiEnable && (4596 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1735_0 <=( _mesh_6_22_io_out_c_0) ^ ((fiEnable && (4597 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_22_io_in_control_0_shift_b <=( _mesh_6_22_io_out_control_0_shift) ^ ((fiEnable && (4598 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_22_io_in_control_0_dataflow_b <=( _mesh_6_22_io_out_control_0_dataflow) ^ ((fiEnable && (4599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_22_io_in_control_0_propagate_b <=( _mesh_6_22_io_out_control_0_propagate) ^ ((fiEnable && (4600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_22_io_out_valid_0) begin
			b_712_0 <=( _mesh_7_22_io_out_b_0) ^ ((fiEnable && (4601 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1736_0 <=( _mesh_7_22_io_out_c_0) ^ ((fiEnable && (4602 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_22_io_in_control_0_shift_b <=( _mesh_7_22_io_out_control_0_shift) ^ ((fiEnable && (4603 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_22_io_in_control_0_dataflow_b <=( _mesh_7_22_io_out_control_0_dataflow) ^ ((fiEnable && (4604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_22_io_in_control_0_propagate_b <=( _mesh_7_22_io_out_control_0_propagate) ^ ((fiEnable && (4605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_22_io_out_valid_0) begin
			b_713_0 <=( _mesh_8_22_io_out_b_0) ^ ((fiEnable && (4606 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1737_0 <=( _mesh_8_22_io_out_c_0) ^ ((fiEnable && (4607 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_22_io_in_control_0_shift_b <=( _mesh_8_22_io_out_control_0_shift) ^ ((fiEnable && (4608 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_22_io_in_control_0_dataflow_b <=( _mesh_8_22_io_out_control_0_dataflow) ^ ((fiEnable && (4609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_22_io_in_control_0_propagate_b <=( _mesh_8_22_io_out_control_0_propagate) ^ ((fiEnable && (4610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_22_io_out_valid_0) begin
			b_714_0 <=( _mesh_9_22_io_out_b_0) ^ ((fiEnable && (4611 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1738_0 <=( _mesh_9_22_io_out_c_0) ^ ((fiEnable && (4612 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_22_io_in_control_0_shift_b <=( _mesh_9_22_io_out_control_0_shift) ^ ((fiEnable && (4613 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_22_io_in_control_0_dataflow_b <=( _mesh_9_22_io_out_control_0_dataflow) ^ ((fiEnable && (4614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_22_io_in_control_0_propagate_b <=( _mesh_9_22_io_out_control_0_propagate) ^ ((fiEnable && (4615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_22_io_out_valid_0) begin
			b_715_0 <=( _mesh_10_22_io_out_b_0) ^ ((fiEnable && (4616 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1739_0 <=( _mesh_10_22_io_out_c_0) ^ ((fiEnable && (4617 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_22_io_in_control_0_shift_b <=( _mesh_10_22_io_out_control_0_shift) ^ ((fiEnable && (4618 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_22_io_in_control_0_dataflow_b <=( _mesh_10_22_io_out_control_0_dataflow) ^ ((fiEnable && (4619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_22_io_in_control_0_propagate_b <=( _mesh_10_22_io_out_control_0_propagate) ^ ((fiEnable && (4620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_22_io_out_valid_0) begin
			b_716_0 <=( _mesh_11_22_io_out_b_0) ^ ((fiEnable && (4621 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1740_0 <=( _mesh_11_22_io_out_c_0) ^ ((fiEnable && (4622 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_22_io_in_control_0_shift_b <=( _mesh_11_22_io_out_control_0_shift) ^ ((fiEnable && (4623 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_22_io_in_control_0_dataflow_b <=( _mesh_11_22_io_out_control_0_dataflow) ^ ((fiEnable && (4624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_22_io_in_control_0_propagate_b <=( _mesh_11_22_io_out_control_0_propagate) ^ ((fiEnable && (4625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_22_io_out_valid_0) begin
			b_717_0 <=( _mesh_12_22_io_out_b_0) ^ ((fiEnable && (4626 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1741_0 <=( _mesh_12_22_io_out_c_0) ^ ((fiEnable && (4627 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_22_io_in_control_0_shift_b <=( _mesh_12_22_io_out_control_0_shift) ^ ((fiEnable && (4628 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_22_io_in_control_0_dataflow_b <=( _mesh_12_22_io_out_control_0_dataflow) ^ ((fiEnable && (4629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_22_io_in_control_0_propagate_b <=( _mesh_12_22_io_out_control_0_propagate) ^ ((fiEnable && (4630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_22_io_out_valid_0) begin
			b_718_0 <=( _mesh_13_22_io_out_b_0) ^ ((fiEnable && (4631 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1742_0 <=( _mesh_13_22_io_out_c_0) ^ ((fiEnable && (4632 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_22_io_in_control_0_shift_b <=( _mesh_13_22_io_out_control_0_shift) ^ ((fiEnable && (4633 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_22_io_in_control_0_dataflow_b <=( _mesh_13_22_io_out_control_0_dataflow) ^ ((fiEnable && (4634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_22_io_in_control_0_propagate_b <=( _mesh_13_22_io_out_control_0_propagate) ^ ((fiEnable && (4635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_22_io_out_valid_0) begin
			b_719_0 <=( _mesh_14_22_io_out_b_0) ^ ((fiEnable && (4636 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1743_0 <=( _mesh_14_22_io_out_c_0) ^ ((fiEnable && (4637 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_22_io_in_control_0_shift_b <=( _mesh_14_22_io_out_control_0_shift) ^ ((fiEnable && (4638 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_22_io_in_control_0_dataflow_b <=( _mesh_14_22_io_out_control_0_dataflow) ^ ((fiEnable && (4639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_22_io_in_control_0_propagate_b <=( _mesh_14_22_io_out_control_0_propagate) ^ ((fiEnable && (4640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_22_io_out_valid_0) begin
			b_720_0 <=( _mesh_15_22_io_out_b_0) ^ ((fiEnable && (4641 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1744_0 <=( _mesh_15_22_io_out_c_0) ^ ((fiEnable && (4642 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_22_io_in_control_0_shift_b <=( _mesh_15_22_io_out_control_0_shift) ^ ((fiEnable && (4643 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_22_io_in_control_0_dataflow_b <=( _mesh_15_22_io_out_control_0_dataflow) ^ ((fiEnable && (4644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_22_io_in_control_0_propagate_b <=( _mesh_15_22_io_out_control_0_propagate) ^ ((fiEnable && (4645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_22_io_out_valid_0) begin
			b_721_0 <=( _mesh_16_22_io_out_b_0) ^ ((fiEnable && (4646 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1745_0 <=( _mesh_16_22_io_out_c_0) ^ ((fiEnable && (4647 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_22_io_in_control_0_shift_b <=( _mesh_16_22_io_out_control_0_shift) ^ ((fiEnable && (4648 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_22_io_in_control_0_dataflow_b <=( _mesh_16_22_io_out_control_0_dataflow) ^ ((fiEnable && (4649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_22_io_in_control_0_propagate_b <=( _mesh_16_22_io_out_control_0_propagate) ^ ((fiEnable && (4650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_22_io_out_valid_0) begin
			b_722_0 <=( _mesh_17_22_io_out_b_0) ^ ((fiEnable && (4651 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1746_0 <=( _mesh_17_22_io_out_c_0) ^ ((fiEnable && (4652 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_22_io_in_control_0_shift_b <=( _mesh_17_22_io_out_control_0_shift) ^ ((fiEnable && (4653 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_22_io_in_control_0_dataflow_b <=( _mesh_17_22_io_out_control_0_dataflow) ^ ((fiEnable && (4654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_22_io_in_control_0_propagate_b <=( _mesh_17_22_io_out_control_0_propagate) ^ ((fiEnable && (4655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_22_io_out_valid_0) begin
			b_723_0 <=( _mesh_18_22_io_out_b_0) ^ ((fiEnable && (4656 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1747_0 <=( _mesh_18_22_io_out_c_0) ^ ((fiEnable && (4657 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_22_io_in_control_0_shift_b <=( _mesh_18_22_io_out_control_0_shift) ^ ((fiEnable && (4658 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_22_io_in_control_0_dataflow_b <=( _mesh_18_22_io_out_control_0_dataflow) ^ ((fiEnable && (4659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_22_io_in_control_0_propagate_b <=( _mesh_18_22_io_out_control_0_propagate) ^ ((fiEnable && (4660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_22_io_out_valid_0) begin
			b_724_0 <=( _mesh_19_22_io_out_b_0) ^ ((fiEnable && (4661 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1748_0 <=( _mesh_19_22_io_out_c_0) ^ ((fiEnable && (4662 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_22_io_in_control_0_shift_b <=( _mesh_19_22_io_out_control_0_shift) ^ ((fiEnable && (4663 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_22_io_in_control_0_dataflow_b <=( _mesh_19_22_io_out_control_0_dataflow) ^ ((fiEnable && (4664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_22_io_in_control_0_propagate_b <=( _mesh_19_22_io_out_control_0_propagate) ^ ((fiEnable && (4665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_22_io_out_valid_0) begin
			b_725_0 <=( _mesh_20_22_io_out_b_0) ^ ((fiEnable && (4666 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1749_0 <=( _mesh_20_22_io_out_c_0) ^ ((fiEnable && (4667 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_22_io_in_control_0_shift_b <=( _mesh_20_22_io_out_control_0_shift) ^ ((fiEnable && (4668 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_22_io_in_control_0_dataflow_b <=( _mesh_20_22_io_out_control_0_dataflow) ^ ((fiEnable && (4669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_22_io_in_control_0_propagate_b <=( _mesh_20_22_io_out_control_0_propagate) ^ ((fiEnable && (4670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_22_io_out_valid_0) begin
			b_726_0 <=( _mesh_21_22_io_out_b_0) ^ ((fiEnable && (4671 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1750_0 <=( _mesh_21_22_io_out_c_0) ^ ((fiEnable && (4672 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_22_io_in_control_0_shift_b <=( _mesh_21_22_io_out_control_0_shift) ^ ((fiEnable && (4673 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_22_io_in_control_0_dataflow_b <=( _mesh_21_22_io_out_control_0_dataflow) ^ ((fiEnable && (4674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_22_io_in_control_0_propagate_b <=( _mesh_21_22_io_out_control_0_propagate) ^ ((fiEnable && (4675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_22_io_out_valid_0) begin
			b_727_0 <=( _mesh_22_22_io_out_b_0) ^ ((fiEnable && (4676 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1751_0 <=( _mesh_22_22_io_out_c_0) ^ ((fiEnable && (4677 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_22_io_in_control_0_shift_b <=( _mesh_22_22_io_out_control_0_shift) ^ ((fiEnable && (4678 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_22_io_in_control_0_dataflow_b <=( _mesh_22_22_io_out_control_0_dataflow) ^ ((fiEnable && (4679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_22_io_in_control_0_propagate_b <=( _mesh_22_22_io_out_control_0_propagate) ^ ((fiEnable && (4680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_22_io_out_valid_0) begin
			b_728_0 <=( _mesh_23_22_io_out_b_0) ^ ((fiEnable && (4681 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1752_0 <=( _mesh_23_22_io_out_c_0) ^ ((fiEnable && (4682 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_22_io_in_control_0_shift_b <=( _mesh_23_22_io_out_control_0_shift) ^ ((fiEnable && (4683 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_22_io_in_control_0_dataflow_b <=( _mesh_23_22_io_out_control_0_dataflow) ^ ((fiEnable && (4684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_22_io_in_control_0_propagate_b <=( _mesh_23_22_io_out_control_0_propagate) ^ ((fiEnable && (4685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_22_io_out_valid_0) begin
			b_729_0 <=( _mesh_24_22_io_out_b_0) ^ ((fiEnable && (4686 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1753_0 <=( _mesh_24_22_io_out_c_0) ^ ((fiEnable && (4687 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_22_io_in_control_0_shift_b <=( _mesh_24_22_io_out_control_0_shift) ^ ((fiEnable && (4688 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_22_io_in_control_0_dataflow_b <=( _mesh_24_22_io_out_control_0_dataflow) ^ ((fiEnable && (4689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_22_io_in_control_0_propagate_b <=( _mesh_24_22_io_out_control_0_propagate) ^ ((fiEnable && (4690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_22_io_out_valid_0) begin
			b_730_0 <=( _mesh_25_22_io_out_b_0) ^ ((fiEnable && (4691 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1754_0 <=( _mesh_25_22_io_out_c_0) ^ ((fiEnable && (4692 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_22_io_in_control_0_shift_b <=( _mesh_25_22_io_out_control_0_shift) ^ ((fiEnable && (4693 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_22_io_in_control_0_dataflow_b <=( _mesh_25_22_io_out_control_0_dataflow) ^ ((fiEnable && (4694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_22_io_in_control_0_propagate_b <=( _mesh_25_22_io_out_control_0_propagate) ^ ((fiEnable && (4695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_22_io_out_valid_0) begin
			b_731_0 <=( _mesh_26_22_io_out_b_0) ^ ((fiEnable && (4696 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1755_0 <=( _mesh_26_22_io_out_c_0) ^ ((fiEnable && (4697 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_22_io_in_control_0_shift_b <=( _mesh_26_22_io_out_control_0_shift) ^ ((fiEnable && (4698 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_22_io_in_control_0_dataflow_b <=( _mesh_26_22_io_out_control_0_dataflow) ^ ((fiEnable && (4699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_22_io_in_control_0_propagate_b <=( _mesh_26_22_io_out_control_0_propagate) ^ ((fiEnable && (4700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_22_io_out_valid_0) begin
			b_732_0 <=( _mesh_27_22_io_out_b_0) ^ ((fiEnable && (4701 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1756_0 <=( _mesh_27_22_io_out_c_0) ^ ((fiEnable && (4702 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_22_io_in_control_0_shift_b <=( _mesh_27_22_io_out_control_0_shift) ^ ((fiEnable && (4703 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_22_io_in_control_0_dataflow_b <=( _mesh_27_22_io_out_control_0_dataflow) ^ ((fiEnable && (4704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_22_io_in_control_0_propagate_b <=( _mesh_27_22_io_out_control_0_propagate) ^ ((fiEnable && (4705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_22_io_out_valid_0) begin
			b_733_0 <=( _mesh_28_22_io_out_b_0) ^ ((fiEnable && (4706 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1757_0 <=( _mesh_28_22_io_out_c_0) ^ ((fiEnable && (4707 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_22_io_in_control_0_shift_b <=( _mesh_28_22_io_out_control_0_shift) ^ ((fiEnable && (4708 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_22_io_in_control_0_dataflow_b <=( _mesh_28_22_io_out_control_0_dataflow) ^ ((fiEnable && (4709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_22_io_in_control_0_propagate_b <=( _mesh_28_22_io_out_control_0_propagate) ^ ((fiEnable && (4710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_22_io_out_valid_0) begin
			b_734_0 <=( _mesh_29_22_io_out_b_0) ^ ((fiEnable && (4711 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1758_0 <=( _mesh_29_22_io_out_c_0) ^ ((fiEnable && (4712 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_22_io_in_control_0_shift_b <=( _mesh_29_22_io_out_control_0_shift) ^ ((fiEnable && (4713 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_22_io_in_control_0_dataflow_b <=( _mesh_29_22_io_out_control_0_dataflow) ^ ((fiEnable && (4714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_22_io_in_control_0_propagate_b <=( _mesh_29_22_io_out_control_0_propagate) ^ ((fiEnable && (4715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_22_io_out_valid_0) begin
			b_735_0 <=( _mesh_30_22_io_out_b_0) ^ ((fiEnable && (4716 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1759_0 <=( _mesh_30_22_io_out_c_0) ^ ((fiEnable && (4717 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_22_io_in_control_0_shift_b <=( _mesh_30_22_io_out_control_0_shift) ^ ((fiEnable && (4718 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_22_io_in_control_0_dataflow_b <=( _mesh_30_22_io_out_control_0_dataflow) ^ ((fiEnable && (4719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_22_io_in_control_0_propagate_b <=( _mesh_30_22_io_out_control_0_propagate) ^ ((fiEnable && (4720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_23_0) begin
			b_736_0 <=( io_in_b_23_0) ^ ((fiEnable && (4721 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1760_0 <=( io_in_d_23_0) ^ ((fiEnable && (4722 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_23_io_in_control_0_shift_b <=( io_in_control_23_0_shift) ^ ((fiEnable && (4723 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_23_io_in_control_0_dataflow_b <=( io_in_control_23_0_dataflow) ^ ((fiEnable && (4724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_23_io_in_control_0_propagate_b <=( io_in_control_23_0_propagate) ^ ((fiEnable && (4725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_23_io_out_valid_0) begin
			b_737_0 <=( _mesh_0_23_io_out_b_0) ^ ((fiEnable && (4726 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1761_0 <=( _mesh_0_23_io_out_c_0) ^ ((fiEnable && (4727 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_23_io_in_control_0_shift_b <=( _mesh_0_23_io_out_control_0_shift) ^ ((fiEnable && (4728 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_23_io_in_control_0_dataflow_b <=( _mesh_0_23_io_out_control_0_dataflow) ^ ((fiEnable && (4729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_23_io_in_control_0_propagate_b <=( _mesh_0_23_io_out_control_0_propagate) ^ ((fiEnable && (4730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_23_io_out_valid_0) begin
			b_738_0 <=( _mesh_1_23_io_out_b_0) ^ ((fiEnable && (4731 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1762_0 <=( _mesh_1_23_io_out_c_0) ^ ((fiEnable && (4732 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_23_io_in_control_0_shift_b <=( _mesh_1_23_io_out_control_0_shift) ^ ((fiEnable && (4733 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_23_io_in_control_0_dataflow_b <=( _mesh_1_23_io_out_control_0_dataflow) ^ ((fiEnable && (4734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_23_io_in_control_0_propagate_b <=( _mesh_1_23_io_out_control_0_propagate) ^ ((fiEnable && (4735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_23_io_out_valid_0) begin
			b_739_0 <=( _mesh_2_23_io_out_b_0) ^ ((fiEnable && (4736 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1763_0 <=( _mesh_2_23_io_out_c_0) ^ ((fiEnable && (4737 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_23_io_in_control_0_shift_b <=( _mesh_2_23_io_out_control_0_shift) ^ ((fiEnable && (4738 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_23_io_in_control_0_dataflow_b <=( _mesh_2_23_io_out_control_0_dataflow) ^ ((fiEnable && (4739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_23_io_in_control_0_propagate_b <=( _mesh_2_23_io_out_control_0_propagate) ^ ((fiEnable && (4740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_23_io_out_valid_0) begin
			b_740_0 <=( _mesh_3_23_io_out_b_0) ^ ((fiEnable && (4741 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1764_0 <=( _mesh_3_23_io_out_c_0) ^ ((fiEnable && (4742 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_23_io_in_control_0_shift_b <=( _mesh_3_23_io_out_control_0_shift) ^ ((fiEnable && (4743 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_23_io_in_control_0_dataflow_b <=( _mesh_3_23_io_out_control_0_dataflow) ^ ((fiEnable && (4744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_23_io_in_control_0_propagate_b <=( _mesh_3_23_io_out_control_0_propagate) ^ ((fiEnable && (4745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_23_io_out_valid_0) begin
			b_741_0 <=( _mesh_4_23_io_out_b_0) ^ ((fiEnable && (4746 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1765_0 <=( _mesh_4_23_io_out_c_0) ^ ((fiEnable && (4747 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_23_io_in_control_0_shift_b <=( _mesh_4_23_io_out_control_0_shift) ^ ((fiEnable && (4748 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_23_io_in_control_0_dataflow_b <=( _mesh_4_23_io_out_control_0_dataflow) ^ ((fiEnable && (4749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_23_io_in_control_0_propagate_b <=( _mesh_4_23_io_out_control_0_propagate) ^ ((fiEnable && (4750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_23_io_out_valid_0) begin
			b_742_0 <=( _mesh_5_23_io_out_b_0) ^ ((fiEnable && (4751 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1766_0 <=( _mesh_5_23_io_out_c_0) ^ ((fiEnable && (4752 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_23_io_in_control_0_shift_b <=( _mesh_5_23_io_out_control_0_shift) ^ ((fiEnable && (4753 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_23_io_in_control_0_dataflow_b <=( _mesh_5_23_io_out_control_0_dataflow) ^ ((fiEnable && (4754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_23_io_in_control_0_propagate_b <=( _mesh_5_23_io_out_control_0_propagate) ^ ((fiEnable && (4755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_23_io_out_valid_0) begin
			b_743_0 <=( _mesh_6_23_io_out_b_0) ^ ((fiEnable && (4756 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1767_0 <=( _mesh_6_23_io_out_c_0) ^ ((fiEnable && (4757 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_23_io_in_control_0_shift_b <=( _mesh_6_23_io_out_control_0_shift) ^ ((fiEnable && (4758 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_23_io_in_control_0_dataflow_b <=( _mesh_6_23_io_out_control_0_dataflow) ^ ((fiEnable && (4759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_23_io_in_control_0_propagate_b <=( _mesh_6_23_io_out_control_0_propagate) ^ ((fiEnable && (4760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_23_io_out_valid_0) begin
			b_744_0 <=( _mesh_7_23_io_out_b_0) ^ ((fiEnable && (4761 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1768_0 <=( _mesh_7_23_io_out_c_0) ^ ((fiEnable && (4762 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_23_io_in_control_0_shift_b <=( _mesh_7_23_io_out_control_0_shift) ^ ((fiEnable && (4763 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_23_io_in_control_0_dataflow_b <=( _mesh_7_23_io_out_control_0_dataflow) ^ ((fiEnable && (4764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_23_io_in_control_0_propagate_b <=( _mesh_7_23_io_out_control_0_propagate) ^ ((fiEnable && (4765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_23_io_out_valid_0) begin
			b_745_0 <=( _mesh_8_23_io_out_b_0) ^ ((fiEnable && (4766 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1769_0 <=( _mesh_8_23_io_out_c_0) ^ ((fiEnable && (4767 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_23_io_in_control_0_shift_b <=( _mesh_8_23_io_out_control_0_shift) ^ ((fiEnable && (4768 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_23_io_in_control_0_dataflow_b <=( _mesh_8_23_io_out_control_0_dataflow) ^ ((fiEnable && (4769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_23_io_in_control_0_propagate_b <=( _mesh_8_23_io_out_control_0_propagate) ^ ((fiEnable && (4770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_23_io_out_valid_0) begin
			b_746_0 <=( _mesh_9_23_io_out_b_0) ^ ((fiEnable && (4771 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1770_0 <=( _mesh_9_23_io_out_c_0) ^ ((fiEnable && (4772 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_23_io_in_control_0_shift_b <=( _mesh_9_23_io_out_control_0_shift) ^ ((fiEnable && (4773 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_23_io_in_control_0_dataflow_b <=( _mesh_9_23_io_out_control_0_dataflow) ^ ((fiEnable && (4774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_23_io_in_control_0_propagate_b <=( _mesh_9_23_io_out_control_0_propagate) ^ ((fiEnable && (4775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_23_io_out_valid_0) begin
			b_747_0 <=( _mesh_10_23_io_out_b_0) ^ ((fiEnable && (4776 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1771_0 <=( _mesh_10_23_io_out_c_0) ^ ((fiEnable && (4777 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_23_io_in_control_0_shift_b <=( _mesh_10_23_io_out_control_0_shift) ^ ((fiEnable && (4778 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_23_io_in_control_0_dataflow_b <=( _mesh_10_23_io_out_control_0_dataflow) ^ ((fiEnable && (4779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_23_io_in_control_0_propagate_b <=( _mesh_10_23_io_out_control_0_propagate) ^ ((fiEnable && (4780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_23_io_out_valid_0) begin
			b_748_0 <=( _mesh_11_23_io_out_b_0) ^ ((fiEnable && (4781 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1772_0 <=( _mesh_11_23_io_out_c_0) ^ ((fiEnable && (4782 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_23_io_in_control_0_shift_b <=( _mesh_11_23_io_out_control_0_shift) ^ ((fiEnable && (4783 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_23_io_in_control_0_dataflow_b <=( _mesh_11_23_io_out_control_0_dataflow) ^ ((fiEnable && (4784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_23_io_in_control_0_propagate_b <=( _mesh_11_23_io_out_control_0_propagate) ^ ((fiEnable && (4785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_23_io_out_valid_0) begin
			b_749_0 <=( _mesh_12_23_io_out_b_0) ^ ((fiEnable && (4786 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1773_0 <=( _mesh_12_23_io_out_c_0) ^ ((fiEnable && (4787 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_23_io_in_control_0_shift_b <=( _mesh_12_23_io_out_control_0_shift) ^ ((fiEnable && (4788 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_23_io_in_control_0_dataflow_b <=( _mesh_12_23_io_out_control_0_dataflow) ^ ((fiEnable && (4789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_23_io_in_control_0_propagate_b <=( _mesh_12_23_io_out_control_0_propagate) ^ ((fiEnable && (4790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_23_io_out_valid_0) begin
			b_750_0 <=( _mesh_13_23_io_out_b_0) ^ ((fiEnable && (4791 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1774_0 <=( _mesh_13_23_io_out_c_0) ^ ((fiEnable && (4792 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_23_io_in_control_0_shift_b <=( _mesh_13_23_io_out_control_0_shift) ^ ((fiEnable && (4793 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_23_io_in_control_0_dataflow_b <=( _mesh_13_23_io_out_control_0_dataflow) ^ ((fiEnable && (4794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_23_io_in_control_0_propagate_b <=( _mesh_13_23_io_out_control_0_propagate) ^ ((fiEnable && (4795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_23_io_out_valid_0) begin
			b_751_0 <=( _mesh_14_23_io_out_b_0) ^ ((fiEnable && (4796 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1775_0 <=( _mesh_14_23_io_out_c_0) ^ ((fiEnable && (4797 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_23_io_in_control_0_shift_b <=( _mesh_14_23_io_out_control_0_shift) ^ ((fiEnable && (4798 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_23_io_in_control_0_dataflow_b <=( _mesh_14_23_io_out_control_0_dataflow) ^ ((fiEnable && (4799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_23_io_in_control_0_propagate_b <=( _mesh_14_23_io_out_control_0_propagate) ^ ((fiEnable && (4800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_23_io_out_valid_0) begin
			b_752_0 <=( _mesh_15_23_io_out_b_0) ^ ((fiEnable && (4801 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1776_0 <=( _mesh_15_23_io_out_c_0) ^ ((fiEnable && (4802 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_23_io_in_control_0_shift_b <=( _mesh_15_23_io_out_control_0_shift) ^ ((fiEnable && (4803 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_23_io_in_control_0_dataflow_b <=( _mesh_15_23_io_out_control_0_dataflow) ^ ((fiEnable && (4804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_23_io_in_control_0_propagate_b <=( _mesh_15_23_io_out_control_0_propagate) ^ ((fiEnable && (4805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_23_io_out_valid_0) begin
			b_753_0 <=( _mesh_16_23_io_out_b_0) ^ ((fiEnable && (4806 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1777_0 <=( _mesh_16_23_io_out_c_0) ^ ((fiEnable && (4807 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_23_io_in_control_0_shift_b <=( _mesh_16_23_io_out_control_0_shift) ^ ((fiEnable && (4808 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_23_io_in_control_0_dataflow_b <=( _mesh_16_23_io_out_control_0_dataflow) ^ ((fiEnable && (4809 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_23_io_in_control_0_propagate_b <=( _mesh_16_23_io_out_control_0_propagate) ^ ((fiEnable && (4810 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_23_io_out_valid_0) begin
			b_754_0 <=( _mesh_17_23_io_out_b_0) ^ ((fiEnable && (4811 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1778_0 <=( _mesh_17_23_io_out_c_0) ^ ((fiEnable && (4812 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_23_io_in_control_0_shift_b <=( _mesh_17_23_io_out_control_0_shift) ^ ((fiEnable && (4813 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_23_io_in_control_0_dataflow_b <=( _mesh_17_23_io_out_control_0_dataflow) ^ ((fiEnable && (4814 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_23_io_in_control_0_propagate_b <=( _mesh_17_23_io_out_control_0_propagate) ^ ((fiEnable && (4815 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_23_io_out_valid_0) begin
			b_755_0 <=( _mesh_18_23_io_out_b_0) ^ ((fiEnable && (4816 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1779_0 <=( _mesh_18_23_io_out_c_0) ^ ((fiEnable && (4817 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_23_io_in_control_0_shift_b <=( _mesh_18_23_io_out_control_0_shift) ^ ((fiEnable && (4818 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_23_io_in_control_0_dataflow_b <=( _mesh_18_23_io_out_control_0_dataflow) ^ ((fiEnable && (4819 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_23_io_in_control_0_propagate_b <=( _mesh_18_23_io_out_control_0_propagate) ^ ((fiEnable && (4820 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_23_io_out_valid_0) begin
			b_756_0 <=( _mesh_19_23_io_out_b_0) ^ ((fiEnable && (4821 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1780_0 <=( _mesh_19_23_io_out_c_0) ^ ((fiEnable && (4822 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_23_io_in_control_0_shift_b <=( _mesh_19_23_io_out_control_0_shift) ^ ((fiEnable && (4823 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_23_io_in_control_0_dataflow_b <=( _mesh_19_23_io_out_control_0_dataflow) ^ ((fiEnable && (4824 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_23_io_in_control_0_propagate_b <=( _mesh_19_23_io_out_control_0_propagate) ^ ((fiEnable && (4825 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_23_io_out_valid_0) begin
			b_757_0 <=( _mesh_20_23_io_out_b_0) ^ ((fiEnable && (4826 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1781_0 <=( _mesh_20_23_io_out_c_0) ^ ((fiEnable && (4827 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_23_io_in_control_0_shift_b <=( _mesh_20_23_io_out_control_0_shift) ^ ((fiEnable && (4828 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_23_io_in_control_0_dataflow_b <=( _mesh_20_23_io_out_control_0_dataflow) ^ ((fiEnable && (4829 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_23_io_in_control_0_propagate_b <=( _mesh_20_23_io_out_control_0_propagate) ^ ((fiEnable && (4830 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_23_io_out_valid_0) begin
			b_758_0 <=( _mesh_21_23_io_out_b_0) ^ ((fiEnable && (4831 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1782_0 <=( _mesh_21_23_io_out_c_0) ^ ((fiEnable && (4832 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_23_io_in_control_0_shift_b <=( _mesh_21_23_io_out_control_0_shift) ^ ((fiEnable && (4833 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_23_io_in_control_0_dataflow_b <=( _mesh_21_23_io_out_control_0_dataflow) ^ ((fiEnable && (4834 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_23_io_in_control_0_propagate_b <=( _mesh_21_23_io_out_control_0_propagate) ^ ((fiEnable && (4835 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_23_io_out_valid_0) begin
			b_759_0 <=( _mesh_22_23_io_out_b_0) ^ ((fiEnable && (4836 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1783_0 <=( _mesh_22_23_io_out_c_0) ^ ((fiEnable && (4837 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_23_io_in_control_0_shift_b <=( _mesh_22_23_io_out_control_0_shift) ^ ((fiEnable && (4838 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_23_io_in_control_0_dataflow_b <=( _mesh_22_23_io_out_control_0_dataflow) ^ ((fiEnable && (4839 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_23_io_in_control_0_propagate_b <=( _mesh_22_23_io_out_control_0_propagate) ^ ((fiEnable && (4840 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_23_io_out_valid_0) begin
			b_760_0 <=( _mesh_23_23_io_out_b_0) ^ ((fiEnable && (4841 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1784_0 <=( _mesh_23_23_io_out_c_0) ^ ((fiEnable && (4842 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_23_io_in_control_0_shift_b <=( _mesh_23_23_io_out_control_0_shift) ^ ((fiEnable && (4843 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_23_io_in_control_0_dataflow_b <=( _mesh_23_23_io_out_control_0_dataflow) ^ ((fiEnable && (4844 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_23_io_in_control_0_propagate_b <=( _mesh_23_23_io_out_control_0_propagate) ^ ((fiEnable && (4845 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_23_io_out_valid_0) begin
			b_761_0 <=( _mesh_24_23_io_out_b_0) ^ ((fiEnable && (4846 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1785_0 <=( _mesh_24_23_io_out_c_0) ^ ((fiEnable && (4847 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_23_io_in_control_0_shift_b <=( _mesh_24_23_io_out_control_0_shift) ^ ((fiEnable && (4848 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_23_io_in_control_0_dataflow_b <=( _mesh_24_23_io_out_control_0_dataflow) ^ ((fiEnable && (4849 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_23_io_in_control_0_propagate_b <=( _mesh_24_23_io_out_control_0_propagate) ^ ((fiEnable && (4850 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_23_io_out_valid_0) begin
			b_762_0 <=( _mesh_25_23_io_out_b_0) ^ ((fiEnable && (4851 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1786_0 <=( _mesh_25_23_io_out_c_0) ^ ((fiEnable && (4852 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_23_io_in_control_0_shift_b <=( _mesh_25_23_io_out_control_0_shift) ^ ((fiEnable && (4853 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_23_io_in_control_0_dataflow_b <=( _mesh_25_23_io_out_control_0_dataflow) ^ ((fiEnable && (4854 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_23_io_in_control_0_propagate_b <=( _mesh_25_23_io_out_control_0_propagate) ^ ((fiEnable && (4855 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_23_io_out_valid_0) begin
			b_763_0 <=( _mesh_26_23_io_out_b_0) ^ ((fiEnable && (4856 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1787_0 <=( _mesh_26_23_io_out_c_0) ^ ((fiEnable && (4857 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_23_io_in_control_0_shift_b <=( _mesh_26_23_io_out_control_0_shift) ^ ((fiEnable && (4858 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_23_io_in_control_0_dataflow_b <=( _mesh_26_23_io_out_control_0_dataflow) ^ ((fiEnable && (4859 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_23_io_in_control_0_propagate_b <=( _mesh_26_23_io_out_control_0_propagate) ^ ((fiEnable && (4860 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_23_io_out_valid_0) begin
			b_764_0 <=( _mesh_27_23_io_out_b_0) ^ ((fiEnable && (4861 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1788_0 <=( _mesh_27_23_io_out_c_0) ^ ((fiEnable && (4862 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_23_io_in_control_0_shift_b <=( _mesh_27_23_io_out_control_0_shift) ^ ((fiEnable && (4863 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_23_io_in_control_0_dataflow_b <=( _mesh_27_23_io_out_control_0_dataflow) ^ ((fiEnable && (4864 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_23_io_in_control_0_propagate_b <=( _mesh_27_23_io_out_control_0_propagate) ^ ((fiEnable && (4865 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_23_io_out_valid_0) begin
			b_765_0 <=( _mesh_28_23_io_out_b_0) ^ ((fiEnable && (4866 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1789_0 <=( _mesh_28_23_io_out_c_0) ^ ((fiEnable && (4867 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_23_io_in_control_0_shift_b <=( _mesh_28_23_io_out_control_0_shift) ^ ((fiEnable && (4868 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_23_io_in_control_0_dataflow_b <=( _mesh_28_23_io_out_control_0_dataflow) ^ ((fiEnable && (4869 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_23_io_in_control_0_propagate_b <=( _mesh_28_23_io_out_control_0_propagate) ^ ((fiEnable && (4870 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_23_io_out_valid_0) begin
			b_766_0 <=( _mesh_29_23_io_out_b_0) ^ ((fiEnable && (4871 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1790_0 <=( _mesh_29_23_io_out_c_0) ^ ((fiEnable && (4872 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_23_io_in_control_0_shift_b <=( _mesh_29_23_io_out_control_0_shift) ^ ((fiEnable && (4873 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_23_io_in_control_0_dataflow_b <=( _mesh_29_23_io_out_control_0_dataflow) ^ ((fiEnable && (4874 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_23_io_in_control_0_propagate_b <=( _mesh_29_23_io_out_control_0_propagate) ^ ((fiEnable && (4875 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_23_io_out_valid_0) begin
			b_767_0 <=( _mesh_30_23_io_out_b_0) ^ ((fiEnable && (4876 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1791_0 <=( _mesh_30_23_io_out_c_0) ^ ((fiEnable && (4877 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_23_io_in_control_0_shift_b <=( _mesh_30_23_io_out_control_0_shift) ^ ((fiEnable && (4878 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_23_io_in_control_0_dataflow_b <=( _mesh_30_23_io_out_control_0_dataflow) ^ ((fiEnable && (4879 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_23_io_in_control_0_propagate_b <=( _mesh_30_23_io_out_control_0_propagate) ^ ((fiEnable && (4880 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_24_0) begin
			b_768_0 <=( io_in_b_24_0) ^ ((fiEnable && (4881 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1792_0 <=( io_in_d_24_0) ^ ((fiEnable && (4882 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_24_io_in_control_0_shift_b <=( io_in_control_24_0_shift) ^ ((fiEnable && (4883 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_24_io_in_control_0_dataflow_b <=( io_in_control_24_0_dataflow) ^ ((fiEnable && (4884 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_24_io_in_control_0_propagate_b <=( io_in_control_24_0_propagate) ^ ((fiEnable && (4885 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_24_io_out_valid_0) begin
			b_769_0 <=( _mesh_0_24_io_out_b_0) ^ ((fiEnable && (4886 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1793_0 <=( _mesh_0_24_io_out_c_0) ^ ((fiEnable && (4887 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_24_io_in_control_0_shift_b <=( _mesh_0_24_io_out_control_0_shift) ^ ((fiEnable && (4888 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_24_io_in_control_0_dataflow_b <=( _mesh_0_24_io_out_control_0_dataflow) ^ ((fiEnable && (4889 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_24_io_in_control_0_propagate_b <=( _mesh_0_24_io_out_control_0_propagate) ^ ((fiEnable && (4890 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_24_io_out_valid_0) begin
			b_770_0 <=( _mesh_1_24_io_out_b_0) ^ ((fiEnable && (4891 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1794_0 <=( _mesh_1_24_io_out_c_0) ^ ((fiEnable && (4892 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_24_io_in_control_0_shift_b <=( _mesh_1_24_io_out_control_0_shift) ^ ((fiEnable && (4893 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_24_io_in_control_0_dataflow_b <=( _mesh_1_24_io_out_control_0_dataflow) ^ ((fiEnable && (4894 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_24_io_in_control_0_propagate_b <=( _mesh_1_24_io_out_control_0_propagate) ^ ((fiEnable && (4895 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_24_io_out_valid_0) begin
			b_771_0 <=( _mesh_2_24_io_out_b_0) ^ ((fiEnable && (4896 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1795_0 <=( _mesh_2_24_io_out_c_0) ^ ((fiEnable && (4897 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_24_io_in_control_0_shift_b <=( _mesh_2_24_io_out_control_0_shift) ^ ((fiEnable && (4898 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_24_io_in_control_0_dataflow_b <=( _mesh_2_24_io_out_control_0_dataflow) ^ ((fiEnable && (4899 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_24_io_in_control_0_propagate_b <=( _mesh_2_24_io_out_control_0_propagate) ^ ((fiEnable && (4900 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_24_io_out_valid_0) begin
			b_772_0 <=( _mesh_3_24_io_out_b_0) ^ ((fiEnable && (4901 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1796_0 <=( _mesh_3_24_io_out_c_0) ^ ((fiEnable && (4902 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_24_io_in_control_0_shift_b <=( _mesh_3_24_io_out_control_0_shift) ^ ((fiEnable && (4903 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_24_io_in_control_0_dataflow_b <=( _mesh_3_24_io_out_control_0_dataflow) ^ ((fiEnable && (4904 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_24_io_in_control_0_propagate_b <=( _mesh_3_24_io_out_control_0_propagate) ^ ((fiEnable && (4905 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_24_io_out_valid_0) begin
			b_773_0 <=( _mesh_4_24_io_out_b_0) ^ ((fiEnable && (4906 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1797_0 <=( _mesh_4_24_io_out_c_0) ^ ((fiEnable && (4907 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_24_io_in_control_0_shift_b <=( _mesh_4_24_io_out_control_0_shift) ^ ((fiEnable && (4908 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_24_io_in_control_0_dataflow_b <=( _mesh_4_24_io_out_control_0_dataflow) ^ ((fiEnable && (4909 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_24_io_in_control_0_propagate_b <=( _mesh_4_24_io_out_control_0_propagate) ^ ((fiEnable && (4910 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_24_io_out_valid_0) begin
			b_774_0 <=( _mesh_5_24_io_out_b_0) ^ ((fiEnable && (4911 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1798_0 <=( _mesh_5_24_io_out_c_0) ^ ((fiEnable && (4912 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_24_io_in_control_0_shift_b <=( _mesh_5_24_io_out_control_0_shift) ^ ((fiEnable && (4913 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_24_io_in_control_0_dataflow_b <=( _mesh_5_24_io_out_control_0_dataflow) ^ ((fiEnable && (4914 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_24_io_in_control_0_propagate_b <=( _mesh_5_24_io_out_control_0_propagate) ^ ((fiEnable && (4915 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_24_io_out_valid_0) begin
			b_775_0 <=( _mesh_6_24_io_out_b_0) ^ ((fiEnable && (4916 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1799_0 <=( _mesh_6_24_io_out_c_0) ^ ((fiEnable && (4917 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_24_io_in_control_0_shift_b <=( _mesh_6_24_io_out_control_0_shift) ^ ((fiEnable && (4918 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_24_io_in_control_0_dataflow_b <=( _mesh_6_24_io_out_control_0_dataflow) ^ ((fiEnable && (4919 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_24_io_in_control_0_propagate_b <=( _mesh_6_24_io_out_control_0_propagate) ^ ((fiEnable && (4920 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_24_io_out_valid_0) begin
			b_776_0 <=( _mesh_7_24_io_out_b_0) ^ ((fiEnable && (4921 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1800_0 <=( _mesh_7_24_io_out_c_0) ^ ((fiEnable && (4922 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_24_io_in_control_0_shift_b <=( _mesh_7_24_io_out_control_0_shift) ^ ((fiEnable && (4923 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_24_io_in_control_0_dataflow_b <=( _mesh_7_24_io_out_control_0_dataflow) ^ ((fiEnable && (4924 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_24_io_in_control_0_propagate_b <=( _mesh_7_24_io_out_control_0_propagate) ^ ((fiEnable && (4925 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_24_io_out_valid_0) begin
			b_777_0 <=( _mesh_8_24_io_out_b_0) ^ ((fiEnable && (4926 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1801_0 <=( _mesh_8_24_io_out_c_0) ^ ((fiEnable && (4927 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_24_io_in_control_0_shift_b <=( _mesh_8_24_io_out_control_0_shift) ^ ((fiEnable && (4928 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_24_io_in_control_0_dataflow_b <=( _mesh_8_24_io_out_control_0_dataflow) ^ ((fiEnable && (4929 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_24_io_in_control_0_propagate_b <=( _mesh_8_24_io_out_control_0_propagate) ^ ((fiEnable && (4930 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_24_io_out_valid_0) begin
			b_778_0 <=( _mesh_9_24_io_out_b_0) ^ ((fiEnable && (4931 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1802_0 <=( _mesh_9_24_io_out_c_0) ^ ((fiEnable && (4932 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_24_io_in_control_0_shift_b <=( _mesh_9_24_io_out_control_0_shift) ^ ((fiEnable && (4933 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_24_io_in_control_0_dataflow_b <=( _mesh_9_24_io_out_control_0_dataflow) ^ ((fiEnable && (4934 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_24_io_in_control_0_propagate_b <=( _mesh_9_24_io_out_control_0_propagate) ^ ((fiEnable && (4935 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_24_io_out_valid_0) begin
			b_779_0 <=( _mesh_10_24_io_out_b_0) ^ ((fiEnable && (4936 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1803_0 <=( _mesh_10_24_io_out_c_0) ^ ((fiEnable && (4937 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_24_io_in_control_0_shift_b <=( _mesh_10_24_io_out_control_0_shift) ^ ((fiEnable && (4938 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_24_io_in_control_0_dataflow_b <=( _mesh_10_24_io_out_control_0_dataflow) ^ ((fiEnable && (4939 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_24_io_in_control_0_propagate_b <=( _mesh_10_24_io_out_control_0_propagate) ^ ((fiEnable && (4940 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_24_io_out_valid_0) begin
			b_780_0 <=( _mesh_11_24_io_out_b_0) ^ ((fiEnable && (4941 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1804_0 <=( _mesh_11_24_io_out_c_0) ^ ((fiEnable && (4942 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_24_io_in_control_0_shift_b <=( _mesh_11_24_io_out_control_0_shift) ^ ((fiEnable && (4943 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_24_io_in_control_0_dataflow_b <=( _mesh_11_24_io_out_control_0_dataflow) ^ ((fiEnable && (4944 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_24_io_in_control_0_propagate_b <=( _mesh_11_24_io_out_control_0_propagate) ^ ((fiEnable && (4945 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_24_io_out_valid_0) begin
			b_781_0 <=( _mesh_12_24_io_out_b_0) ^ ((fiEnable && (4946 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1805_0 <=( _mesh_12_24_io_out_c_0) ^ ((fiEnable && (4947 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_24_io_in_control_0_shift_b <=( _mesh_12_24_io_out_control_0_shift) ^ ((fiEnable && (4948 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_24_io_in_control_0_dataflow_b <=( _mesh_12_24_io_out_control_0_dataflow) ^ ((fiEnable && (4949 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_24_io_in_control_0_propagate_b <=( _mesh_12_24_io_out_control_0_propagate) ^ ((fiEnable && (4950 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_24_io_out_valid_0) begin
			b_782_0 <=( _mesh_13_24_io_out_b_0) ^ ((fiEnable && (4951 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1806_0 <=( _mesh_13_24_io_out_c_0) ^ ((fiEnable && (4952 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_24_io_in_control_0_shift_b <=( _mesh_13_24_io_out_control_0_shift) ^ ((fiEnable && (4953 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_24_io_in_control_0_dataflow_b <=( _mesh_13_24_io_out_control_0_dataflow) ^ ((fiEnable && (4954 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_24_io_in_control_0_propagate_b <=( _mesh_13_24_io_out_control_0_propagate) ^ ((fiEnable && (4955 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_24_io_out_valid_0) begin
			b_783_0 <=( _mesh_14_24_io_out_b_0) ^ ((fiEnable && (4956 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1807_0 <=( _mesh_14_24_io_out_c_0) ^ ((fiEnable && (4957 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_24_io_in_control_0_shift_b <=( _mesh_14_24_io_out_control_0_shift) ^ ((fiEnable && (4958 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_24_io_in_control_0_dataflow_b <=( _mesh_14_24_io_out_control_0_dataflow) ^ ((fiEnable && (4959 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_24_io_in_control_0_propagate_b <=( _mesh_14_24_io_out_control_0_propagate) ^ ((fiEnable && (4960 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_24_io_out_valid_0) begin
			b_784_0 <=( _mesh_15_24_io_out_b_0) ^ ((fiEnable && (4961 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1808_0 <=( _mesh_15_24_io_out_c_0) ^ ((fiEnable && (4962 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_24_io_in_control_0_shift_b <=( _mesh_15_24_io_out_control_0_shift) ^ ((fiEnable && (4963 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_24_io_in_control_0_dataflow_b <=( _mesh_15_24_io_out_control_0_dataflow) ^ ((fiEnable && (4964 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_24_io_in_control_0_propagate_b <=( _mesh_15_24_io_out_control_0_propagate) ^ ((fiEnable && (4965 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_24_io_out_valid_0) begin
			b_785_0 <=( _mesh_16_24_io_out_b_0) ^ ((fiEnable && (4966 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1809_0 <=( _mesh_16_24_io_out_c_0) ^ ((fiEnable && (4967 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_24_io_in_control_0_shift_b <=( _mesh_16_24_io_out_control_0_shift) ^ ((fiEnable && (4968 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_24_io_in_control_0_dataflow_b <=( _mesh_16_24_io_out_control_0_dataflow) ^ ((fiEnable && (4969 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_24_io_in_control_0_propagate_b <=( _mesh_16_24_io_out_control_0_propagate) ^ ((fiEnable && (4970 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_24_io_out_valid_0) begin
			b_786_0 <=( _mesh_17_24_io_out_b_0) ^ ((fiEnable && (4971 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1810_0 <=( _mesh_17_24_io_out_c_0) ^ ((fiEnable && (4972 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_24_io_in_control_0_shift_b <=( _mesh_17_24_io_out_control_0_shift) ^ ((fiEnable && (4973 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_24_io_in_control_0_dataflow_b <=( _mesh_17_24_io_out_control_0_dataflow) ^ ((fiEnable && (4974 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_24_io_in_control_0_propagate_b <=( _mesh_17_24_io_out_control_0_propagate) ^ ((fiEnable && (4975 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_24_io_out_valid_0) begin
			b_787_0 <=( _mesh_18_24_io_out_b_0) ^ ((fiEnable && (4976 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1811_0 <=( _mesh_18_24_io_out_c_0) ^ ((fiEnable && (4977 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_24_io_in_control_0_shift_b <=( _mesh_18_24_io_out_control_0_shift) ^ ((fiEnable && (4978 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_24_io_in_control_0_dataflow_b <=( _mesh_18_24_io_out_control_0_dataflow) ^ ((fiEnable && (4979 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_24_io_in_control_0_propagate_b <=( _mesh_18_24_io_out_control_0_propagate) ^ ((fiEnable && (4980 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_24_io_out_valid_0) begin
			b_788_0 <=( _mesh_19_24_io_out_b_0) ^ ((fiEnable && (4981 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1812_0 <=( _mesh_19_24_io_out_c_0) ^ ((fiEnable && (4982 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_24_io_in_control_0_shift_b <=( _mesh_19_24_io_out_control_0_shift) ^ ((fiEnable && (4983 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_24_io_in_control_0_dataflow_b <=( _mesh_19_24_io_out_control_0_dataflow) ^ ((fiEnable && (4984 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_24_io_in_control_0_propagate_b <=( _mesh_19_24_io_out_control_0_propagate) ^ ((fiEnable && (4985 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_24_io_out_valid_0) begin
			b_789_0 <=( _mesh_20_24_io_out_b_0) ^ ((fiEnable && (4986 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1813_0 <=( _mesh_20_24_io_out_c_0) ^ ((fiEnable && (4987 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_24_io_in_control_0_shift_b <=( _mesh_20_24_io_out_control_0_shift) ^ ((fiEnable && (4988 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_24_io_in_control_0_dataflow_b <=( _mesh_20_24_io_out_control_0_dataflow) ^ ((fiEnable && (4989 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_24_io_in_control_0_propagate_b <=( _mesh_20_24_io_out_control_0_propagate) ^ ((fiEnable && (4990 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_24_io_out_valid_0) begin
			b_790_0 <=( _mesh_21_24_io_out_b_0) ^ ((fiEnable && (4991 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1814_0 <=( _mesh_21_24_io_out_c_0) ^ ((fiEnable && (4992 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_24_io_in_control_0_shift_b <=( _mesh_21_24_io_out_control_0_shift) ^ ((fiEnable && (4993 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_24_io_in_control_0_dataflow_b <=( _mesh_21_24_io_out_control_0_dataflow) ^ ((fiEnable && (4994 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_24_io_in_control_0_propagate_b <=( _mesh_21_24_io_out_control_0_propagate) ^ ((fiEnable && (4995 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_24_io_out_valid_0) begin
			b_791_0 <=( _mesh_22_24_io_out_b_0) ^ ((fiEnable && (4996 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1815_0 <=( _mesh_22_24_io_out_c_0) ^ ((fiEnable && (4997 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_24_io_in_control_0_shift_b <=( _mesh_22_24_io_out_control_0_shift) ^ ((fiEnable && (4998 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_24_io_in_control_0_dataflow_b <=( _mesh_22_24_io_out_control_0_dataflow) ^ ((fiEnable && (4999 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_24_io_in_control_0_propagate_b <=( _mesh_22_24_io_out_control_0_propagate) ^ ((fiEnable && (5000 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_24_io_out_valid_0) begin
			b_792_0 <=( _mesh_23_24_io_out_b_0) ^ ((fiEnable && (5001 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1816_0 <=( _mesh_23_24_io_out_c_0) ^ ((fiEnable && (5002 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_24_io_in_control_0_shift_b <=( _mesh_23_24_io_out_control_0_shift) ^ ((fiEnable && (5003 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_24_io_in_control_0_dataflow_b <=( _mesh_23_24_io_out_control_0_dataflow) ^ ((fiEnable && (5004 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_24_io_in_control_0_propagate_b <=( _mesh_23_24_io_out_control_0_propagate) ^ ((fiEnable && (5005 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_24_io_out_valid_0) begin
			b_793_0 <=( _mesh_24_24_io_out_b_0) ^ ((fiEnable && (5006 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1817_0 <=( _mesh_24_24_io_out_c_0) ^ ((fiEnable && (5007 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_24_io_in_control_0_shift_b <=( _mesh_24_24_io_out_control_0_shift) ^ ((fiEnable && (5008 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_24_io_in_control_0_dataflow_b <=( _mesh_24_24_io_out_control_0_dataflow) ^ ((fiEnable && (5009 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_24_io_in_control_0_propagate_b <=( _mesh_24_24_io_out_control_0_propagate) ^ ((fiEnable && (5010 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_24_io_out_valid_0) begin
			b_794_0 <=( _mesh_25_24_io_out_b_0) ^ ((fiEnable && (5011 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1818_0 <=( _mesh_25_24_io_out_c_0) ^ ((fiEnable && (5012 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_24_io_in_control_0_shift_b <=( _mesh_25_24_io_out_control_0_shift) ^ ((fiEnable && (5013 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_24_io_in_control_0_dataflow_b <=( _mesh_25_24_io_out_control_0_dataflow) ^ ((fiEnable && (5014 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_24_io_in_control_0_propagate_b <=( _mesh_25_24_io_out_control_0_propagate) ^ ((fiEnable && (5015 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_24_io_out_valid_0) begin
			b_795_0 <=( _mesh_26_24_io_out_b_0) ^ ((fiEnable && (5016 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1819_0 <=( _mesh_26_24_io_out_c_0) ^ ((fiEnable && (5017 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_24_io_in_control_0_shift_b <=( _mesh_26_24_io_out_control_0_shift) ^ ((fiEnable && (5018 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_24_io_in_control_0_dataflow_b <=( _mesh_26_24_io_out_control_0_dataflow) ^ ((fiEnable && (5019 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_24_io_in_control_0_propagate_b <=( _mesh_26_24_io_out_control_0_propagate) ^ ((fiEnable && (5020 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_24_io_out_valid_0) begin
			b_796_0 <=( _mesh_27_24_io_out_b_0) ^ ((fiEnable && (5021 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1820_0 <=( _mesh_27_24_io_out_c_0) ^ ((fiEnable && (5022 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_24_io_in_control_0_shift_b <=( _mesh_27_24_io_out_control_0_shift) ^ ((fiEnable && (5023 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_24_io_in_control_0_dataflow_b <=( _mesh_27_24_io_out_control_0_dataflow) ^ ((fiEnable && (5024 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_24_io_in_control_0_propagate_b <=( _mesh_27_24_io_out_control_0_propagate) ^ ((fiEnable && (5025 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_24_io_out_valid_0) begin
			b_797_0 <=( _mesh_28_24_io_out_b_0) ^ ((fiEnable && (5026 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1821_0 <=( _mesh_28_24_io_out_c_0) ^ ((fiEnable && (5027 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_24_io_in_control_0_shift_b <=( _mesh_28_24_io_out_control_0_shift) ^ ((fiEnable && (5028 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_24_io_in_control_0_dataflow_b <=( _mesh_28_24_io_out_control_0_dataflow) ^ ((fiEnable && (5029 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_24_io_in_control_0_propagate_b <=( _mesh_28_24_io_out_control_0_propagate) ^ ((fiEnable && (5030 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_24_io_out_valid_0) begin
			b_798_0 <=( _mesh_29_24_io_out_b_0) ^ ((fiEnable && (5031 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1822_0 <=( _mesh_29_24_io_out_c_0) ^ ((fiEnable && (5032 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_24_io_in_control_0_shift_b <=( _mesh_29_24_io_out_control_0_shift) ^ ((fiEnable && (5033 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_24_io_in_control_0_dataflow_b <=( _mesh_29_24_io_out_control_0_dataflow) ^ ((fiEnable && (5034 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_24_io_in_control_0_propagate_b <=( _mesh_29_24_io_out_control_0_propagate) ^ ((fiEnable && (5035 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_24_io_out_valid_0) begin
			b_799_0 <=( _mesh_30_24_io_out_b_0) ^ ((fiEnable && (5036 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1823_0 <=( _mesh_30_24_io_out_c_0) ^ ((fiEnable && (5037 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_24_io_in_control_0_shift_b <=( _mesh_30_24_io_out_control_0_shift) ^ ((fiEnable && (5038 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_24_io_in_control_0_dataflow_b <=( _mesh_30_24_io_out_control_0_dataflow) ^ ((fiEnable && (5039 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_24_io_in_control_0_propagate_b <=( _mesh_30_24_io_out_control_0_propagate) ^ ((fiEnable && (5040 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_25_0) begin
			b_800_0 <=( io_in_b_25_0) ^ ((fiEnable && (5041 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1824_0 <=( io_in_d_25_0) ^ ((fiEnable && (5042 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_25_io_in_control_0_shift_b <=( io_in_control_25_0_shift) ^ ((fiEnable && (5043 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_25_io_in_control_0_dataflow_b <=( io_in_control_25_0_dataflow) ^ ((fiEnable && (5044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_25_io_in_control_0_propagate_b <=( io_in_control_25_0_propagate) ^ ((fiEnable && (5045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_25_io_out_valid_0) begin
			b_801_0 <=( _mesh_0_25_io_out_b_0) ^ ((fiEnable && (5046 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1825_0 <=( _mesh_0_25_io_out_c_0) ^ ((fiEnable && (5047 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_25_io_in_control_0_shift_b <=( _mesh_0_25_io_out_control_0_shift) ^ ((fiEnable && (5048 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_25_io_in_control_0_dataflow_b <=( _mesh_0_25_io_out_control_0_dataflow) ^ ((fiEnable && (5049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_25_io_in_control_0_propagate_b <=( _mesh_0_25_io_out_control_0_propagate) ^ ((fiEnable && (5050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_25_io_out_valid_0) begin
			b_802_0 <=( _mesh_1_25_io_out_b_0) ^ ((fiEnable && (5051 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1826_0 <=( _mesh_1_25_io_out_c_0) ^ ((fiEnable && (5052 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_25_io_in_control_0_shift_b <=( _mesh_1_25_io_out_control_0_shift) ^ ((fiEnable && (5053 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_25_io_in_control_0_dataflow_b <=( _mesh_1_25_io_out_control_0_dataflow) ^ ((fiEnable && (5054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_25_io_in_control_0_propagate_b <=( _mesh_1_25_io_out_control_0_propagate) ^ ((fiEnable && (5055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_25_io_out_valid_0) begin
			b_803_0 <=( _mesh_2_25_io_out_b_0) ^ ((fiEnable && (5056 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1827_0 <=( _mesh_2_25_io_out_c_0) ^ ((fiEnable && (5057 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_25_io_in_control_0_shift_b <=( _mesh_2_25_io_out_control_0_shift) ^ ((fiEnable && (5058 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_25_io_in_control_0_dataflow_b <=( _mesh_2_25_io_out_control_0_dataflow) ^ ((fiEnable && (5059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_25_io_in_control_0_propagate_b <=( _mesh_2_25_io_out_control_0_propagate) ^ ((fiEnable && (5060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_25_io_out_valid_0) begin
			b_804_0 <=( _mesh_3_25_io_out_b_0) ^ ((fiEnable && (5061 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1828_0 <=( _mesh_3_25_io_out_c_0) ^ ((fiEnable && (5062 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_25_io_in_control_0_shift_b <=( _mesh_3_25_io_out_control_0_shift) ^ ((fiEnable && (5063 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_25_io_in_control_0_dataflow_b <=( _mesh_3_25_io_out_control_0_dataflow) ^ ((fiEnable && (5064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_25_io_in_control_0_propagate_b <=( _mesh_3_25_io_out_control_0_propagate) ^ ((fiEnable && (5065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_25_io_out_valid_0) begin
			b_805_0 <=( _mesh_4_25_io_out_b_0) ^ ((fiEnable && (5066 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1829_0 <=( _mesh_4_25_io_out_c_0) ^ ((fiEnable && (5067 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_25_io_in_control_0_shift_b <=( _mesh_4_25_io_out_control_0_shift) ^ ((fiEnable && (5068 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_25_io_in_control_0_dataflow_b <=( _mesh_4_25_io_out_control_0_dataflow) ^ ((fiEnable && (5069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_25_io_in_control_0_propagate_b <=( _mesh_4_25_io_out_control_0_propagate) ^ ((fiEnable && (5070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_25_io_out_valid_0) begin
			b_806_0 <=( _mesh_5_25_io_out_b_0) ^ ((fiEnable && (5071 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1830_0 <=( _mesh_5_25_io_out_c_0) ^ ((fiEnable && (5072 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_25_io_in_control_0_shift_b <=( _mesh_5_25_io_out_control_0_shift) ^ ((fiEnable && (5073 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_25_io_in_control_0_dataflow_b <=( _mesh_5_25_io_out_control_0_dataflow) ^ ((fiEnable && (5074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_25_io_in_control_0_propagate_b <=( _mesh_5_25_io_out_control_0_propagate) ^ ((fiEnable && (5075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_25_io_out_valid_0) begin
			b_807_0 <=( _mesh_6_25_io_out_b_0) ^ ((fiEnable && (5076 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1831_0 <=( _mesh_6_25_io_out_c_0) ^ ((fiEnable && (5077 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_25_io_in_control_0_shift_b <=( _mesh_6_25_io_out_control_0_shift) ^ ((fiEnable && (5078 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_25_io_in_control_0_dataflow_b <=( _mesh_6_25_io_out_control_0_dataflow) ^ ((fiEnable && (5079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_25_io_in_control_0_propagate_b <=( _mesh_6_25_io_out_control_0_propagate) ^ ((fiEnable && (5080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_25_io_out_valid_0) begin
			b_808_0 <=( _mesh_7_25_io_out_b_0) ^ ((fiEnable && (5081 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1832_0 <=( _mesh_7_25_io_out_c_0) ^ ((fiEnable && (5082 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_25_io_in_control_0_shift_b <=( _mesh_7_25_io_out_control_0_shift) ^ ((fiEnable && (5083 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_25_io_in_control_0_dataflow_b <=( _mesh_7_25_io_out_control_0_dataflow) ^ ((fiEnable && (5084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_25_io_in_control_0_propagate_b <=( _mesh_7_25_io_out_control_0_propagate) ^ ((fiEnable && (5085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_25_io_out_valid_0) begin
			b_809_0 <=( _mesh_8_25_io_out_b_0) ^ ((fiEnable && (5086 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1833_0 <=( _mesh_8_25_io_out_c_0) ^ ((fiEnable && (5087 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_25_io_in_control_0_shift_b <=( _mesh_8_25_io_out_control_0_shift) ^ ((fiEnable && (5088 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_25_io_in_control_0_dataflow_b <=( _mesh_8_25_io_out_control_0_dataflow) ^ ((fiEnable && (5089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_25_io_in_control_0_propagate_b <=( _mesh_8_25_io_out_control_0_propagate) ^ ((fiEnable && (5090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_25_io_out_valid_0) begin
			b_810_0 <=( _mesh_9_25_io_out_b_0) ^ ((fiEnable && (5091 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1834_0 <=( _mesh_9_25_io_out_c_0) ^ ((fiEnable && (5092 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_25_io_in_control_0_shift_b <=( _mesh_9_25_io_out_control_0_shift) ^ ((fiEnable && (5093 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_25_io_in_control_0_dataflow_b <=( _mesh_9_25_io_out_control_0_dataflow) ^ ((fiEnable && (5094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_25_io_in_control_0_propagate_b <=( _mesh_9_25_io_out_control_0_propagate) ^ ((fiEnable && (5095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_25_io_out_valid_0) begin
			b_811_0 <=( _mesh_10_25_io_out_b_0) ^ ((fiEnable && (5096 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1835_0 <=( _mesh_10_25_io_out_c_0) ^ ((fiEnable && (5097 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_25_io_in_control_0_shift_b <=( _mesh_10_25_io_out_control_0_shift) ^ ((fiEnable && (5098 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_25_io_in_control_0_dataflow_b <=( _mesh_10_25_io_out_control_0_dataflow) ^ ((fiEnable && (5099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_25_io_in_control_0_propagate_b <=( _mesh_10_25_io_out_control_0_propagate) ^ ((fiEnable && (5100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_25_io_out_valid_0) begin
			b_812_0 <=( _mesh_11_25_io_out_b_0) ^ ((fiEnable && (5101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1836_0 <=( _mesh_11_25_io_out_c_0) ^ ((fiEnable && (5102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_25_io_in_control_0_shift_b <=( _mesh_11_25_io_out_control_0_shift) ^ ((fiEnable && (5103 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_25_io_in_control_0_dataflow_b <=( _mesh_11_25_io_out_control_0_dataflow) ^ ((fiEnable && (5104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_25_io_in_control_0_propagate_b <=( _mesh_11_25_io_out_control_0_propagate) ^ ((fiEnable && (5105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_25_io_out_valid_0) begin
			b_813_0 <=( _mesh_12_25_io_out_b_0) ^ ((fiEnable && (5106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1837_0 <=( _mesh_12_25_io_out_c_0) ^ ((fiEnable && (5107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_25_io_in_control_0_shift_b <=( _mesh_12_25_io_out_control_0_shift) ^ ((fiEnable && (5108 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_25_io_in_control_0_dataflow_b <=( _mesh_12_25_io_out_control_0_dataflow) ^ ((fiEnable && (5109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_25_io_in_control_0_propagate_b <=( _mesh_12_25_io_out_control_0_propagate) ^ ((fiEnable && (5110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_25_io_out_valid_0) begin
			b_814_0 <=( _mesh_13_25_io_out_b_0) ^ ((fiEnable && (5111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1838_0 <=( _mesh_13_25_io_out_c_0) ^ ((fiEnable && (5112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_25_io_in_control_0_shift_b <=( _mesh_13_25_io_out_control_0_shift) ^ ((fiEnable && (5113 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_25_io_in_control_0_dataflow_b <=( _mesh_13_25_io_out_control_0_dataflow) ^ ((fiEnable && (5114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_25_io_in_control_0_propagate_b <=( _mesh_13_25_io_out_control_0_propagate) ^ ((fiEnable && (5115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_25_io_out_valid_0) begin
			b_815_0 <=( _mesh_14_25_io_out_b_0) ^ ((fiEnable && (5116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1839_0 <=( _mesh_14_25_io_out_c_0) ^ ((fiEnable && (5117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_25_io_in_control_0_shift_b <=( _mesh_14_25_io_out_control_0_shift) ^ ((fiEnable && (5118 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_25_io_in_control_0_dataflow_b <=( _mesh_14_25_io_out_control_0_dataflow) ^ ((fiEnable && (5119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_25_io_in_control_0_propagate_b <=( _mesh_14_25_io_out_control_0_propagate) ^ ((fiEnable && (5120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_25_io_out_valid_0) begin
			b_816_0 <=( _mesh_15_25_io_out_b_0) ^ ((fiEnable && (5121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1840_0 <=( _mesh_15_25_io_out_c_0) ^ ((fiEnable && (5122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_25_io_in_control_0_shift_b <=( _mesh_15_25_io_out_control_0_shift) ^ ((fiEnable && (5123 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_25_io_in_control_0_dataflow_b <=( _mesh_15_25_io_out_control_0_dataflow) ^ ((fiEnable && (5124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_25_io_in_control_0_propagate_b <=( _mesh_15_25_io_out_control_0_propagate) ^ ((fiEnable && (5125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_25_io_out_valid_0) begin
			b_817_0 <=( _mesh_16_25_io_out_b_0) ^ ((fiEnable && (5126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1841_0 <=( _mesh_16_25_io_out_c_0) ^ ((fiEnable && (5127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_25_io_in_control_0_shift_b <=( _mesh_16_25_io_out_control_0_shift) ^ ((fiEnable && (5128 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_25_io_in_control_0_dataflow_b <=( _mesh_16_25_io_out_control_0_dataflow) ^ ((fiEnable && (5129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_25_io_in_control_0_propagate_b <=( _mesh_16_25_io_out_control_0_propagate) ^ ((fiEnable && (5130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_25_io_out_valid_0) begin
			b_818_0 <=( _mesh_17_25_io_out_b_0) ^ ((fiEnable && (5131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1842_0 <=( _mesh_17_25_io_out_c_0) ^ ((fiEnable && (5132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_25_io_in_control_0_shift_b <=( _mesh_17_25_io_out_control_0_shift) ^ ((fiEnable && (5133 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_25_io_in_control_0_dataflow_b <=( _mesh_17_25_io_out_control_0_dataflow) ^ ((fiEnable && (5134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_25_io_in_control_0_propagate_b <=( _mesh_17_25_io_out_control_0_propagate) ^ ((fiEnable && (5135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_25_io_out_valid_0) begin
			b_819_0 <=( _mesh_18_25_io_out_b_0) ^ ((fiEnable && (5136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1843_0 <=( _mesh_18_25_io_out_c_0) ^ ((fiEnable && (5137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_25_io_in_control_0_shift_b <=( _mesh_18_25_io_out_control_0_shift) ^ ((fiEnable && (5138 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_25_io_in_control_0_dataflow_b <=( _mesh_18_25_io_out_control_0_dataflow) ^ ((fiEnable && (5139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_25_io_in_control_0_propagate_b <=( _mesh_18_25_io_out_control_0_propagate) ^ ((fiEnable && (5140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_25_io_out_valid_0) begin
			b_820_0 <=( _mesh_19_25_io_out_b_0) ^ ((fiEnable && (5141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1844_0 <=( _mesh_19_25_io_out_c_0) ^ ((fiEnable && (5142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_25_io_in_control_0_shift_b <=( _mesh_19_25_io_out_control_0_shift) ^ ((fiEnable && (5143 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_25_io_in_control_0_dataflow_b <=( _mesh_19_25_io_out_control_0_dataflow) ^ ((fiEnable && (5144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_25_io_in_control_0_propagate_b <=( _mesh_19_25_io_out_control_0_propagate) ^ ((fiEnable && (5145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_25_io_out_valid_0) begin
			b_821_0 <=( _mesh_20_25_io_out_b_0) ^ ((fiEnable && (5146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1845_0 <=( _mesh_20_25_io_out_c_0) ^ ((fiEnable && (5147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_25_io_in_control_0_shift_b <=( _mesh_20_25_io_out_control_0_shift) ^ ((fiEnable && (5148 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_25_io_in_control_0_dataflow_b <=( _mesh_20_25_io_out_control_0_dataflow) ^ ((fiEnable && (5149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_25_io_in_control_0_propagate_b <=( _mesh_20_25_io_out_control_0_propagate) ^ ((fiEnable && (5150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_25_io_out_valid_0) begin
			b_822_0 <=( _mesh_21_25_io_out_b_0) ^ ((fiEnable && (5151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1846_0 <=( _mesh_21_25_io_out_c_0) ^ ((fiEnable && (5152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_25_io_in_control_0_shift_b <=( _mesh_21_25_io_out_control_0_shift) ^ ((fiEnable && (5153 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_25_io_in_control_0_dataflow_b <=( _mesh_21_25_io_out_control_0_dataflow) ^ ((fiEnable && (5154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_25_io_in_control_0_propagate_b <=( _mesh_21_25_io_out_control_0_propagate) ^ ((fiEnable && (5155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_25_io_out_valid_0) begin
			b_823_0 <=( _mesh_22_25_io_out_b_0) ^ ((fiEnable && (5156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1847_0 <=( _mesh_22_25_io_out_c_0) ^ ((fiEnable && (5157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_25_io_in_control_0_shift_b <=( _mesh_22_25_io_out_control_0_shift) ^ ((fiEnable && (5158 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_25_io_in_control_0_dataflow_b <=( _mesh_22_25_io_out_control_0_dataflow) ^ ((fiEnable && (5159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_25_io_in_control_0_propagate_b <=( _mesh_22_25_io_out_control_0_propagate) ^ ((fiEnable && (5160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_25_io_out_valid_0) begin
			b_824_0 <=( _mesh_23_25_io_out_b_0) ^ ((fiEnable && (5161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1848_0 <=( _mesh_23_25_io_out_c_0) ^ ((fiEnable && (5162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_25_io_in_control_0_shift_b <=( _mesh_23_25_io_out_control_0_shift) ^ ((fiEnable && (5163 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_25_io_in_control_0_dataflow_b <=( _mesh_23_25_io_out_control_0_dataflow) ^ ((fiEnable && (5164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_25_io_in_control_0_propagate_b <=( _mesh_23_25_io_out_control_0_propagate) ^ ((fiEnable && (5165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_25_io_out_valid_0) begin
			b_825_0 <=( _mesh_24_25_io_out_b_0) ^ ((fiEnable && (5166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1849_0 <=( _mesh_24_25_io_out_c_0) ^ ((fiEnable && (5167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_25_io_in_control_0_shift_b <=( _mesh_24_25_io_out_control_0_shift) ^ ((fiEnable && (5168 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_25_io_in_control_0_dataflow_b <=( _mesh_24_25_io_out_control_0_dataflow) ^ ((fiEnable && (5169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_25_io_in_control_0_propagate_b <=( _mesh_24_25_io_out_control_0_propagate) ^ ((fiEnable && (5170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_25_io_out_valid_0) begin
			b_826_0 <=( _mesh_25_25_io_out_b_0) ^ ((fiEnable && (5171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1850_0 <=( _mesh_25_25_io_out_c_0) ^ ((fiEnable && (5172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_25_io_in_control_0_shift_b <=( _mesh_25_25_io_out_control_0_shift) ^ ((fiEnable && (5173 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_25_io_in_control_0_dataflow_b <=( _mesh_25_25_io_out_control_0_dataflow) ^ ((fiEnable && (5174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_25_io_in_control_0_propagate_b <=( _mesh_25_25_io_out_control_0_propagate) ^ ((fiEnable && (5175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_25_io_out_valid_0) begin
			b_827_0 <=( _mesh_26_25_io_out_b_0) ^ ((fiEnable && (5176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1851_0 <=( _mesh_26_25_io_out_c_0) ^ ((fiEnable && (5177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_25_io_in_control_0_shift_b <=( _mesh_26_25_io_out_control_0_shift) ^ ((fiEnable && (5178 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_25_io_in_control_0_dataflow_b <=( _mesh_26_25_io_out_control_0_dataflow) ^ ((fiEnable && (5179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_25_io_in_control_0_propagate_b <=( _mesh_26_25_io_out_control_0_propagate) ^ ((fiEnable && (5180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_25_io_out_valid_0) begin
			b_828_0 <=( _mesh_27_25_io_out_b_0) ^ ((fiEnable && (5181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1852_0 <=( _mesh_27_25_io_out_c_0) ^ ((fiEnable && (5182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_25_io_in_control_0_shift_b <=( _mesh_27_25_io_out_control_0_shift) ^ ((fiEnable && (5183 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_25_io_in_control_0_dataflow_b <=( _mesh_27_25_io_out_control_0_dataflow) ^ ((fiEnable && (5184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_25_io_in_control_0_propagate_b <=( _mesh_27_25_io_out_control_0_propagate) ^ ((fiEnable && (5185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_25_io_out_valid_0) begin
			b_829_0 <=( _mesh_28_25_io_out_b_0) ^ ((fiEnable && (5186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1853_0 <=( _mesh_28_25_io_out_c_0) ^ ((fiEnable && (5187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_25_io_in_control_0_shift_b <=( _mesh_28_25_io_out_control_0_shift) ^ ((fiEnable && (5188 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_25_io_in_control_0_dataflow_b <=( _mesh_28_25_io_out_control_0_dataflow) ^ ((fiEnable && (5189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_25_io_in_control_0_propagate_b <=( _mesh_28_25_io_out_control_0_propagate) ^ ((fiEnable && (5190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_25_io_out_valid_0) begin
			b_830_0 <=( _mesh_29_25_io_out_b_0) ^ ((fiEnable && (5191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1854_0 <=( _mesh_29_25_io_out_c_0) ^ ((fiEnable && (5192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_25_io_in_control_0_shift_b <=( _mesh_29_25_io_out_control_0_shift) ^ ((fiEnable && (5193 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_25_io_in_control_0_dataflow_b <=( _mesh_29_25_io_out_control_0_dataflow) ^ ((fiEnable && (5194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_25_io_in_control_0_propagate_b <=( _mesh_29_25_io_out_control_0_propagate) ^ ((fiEnable && (5195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_25_io_out_valid_0) begin
			b_831_0 <=( _mesh_30_25_io_out_b_0) ^ ((fiEnable && (5196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1855_0 <=( _mesh_30_25_io_out_c_0) ^ ((fiEnable && (5197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_25_io_in_control_0_shift_b <=( _mesh_30_25_io_out_control_0_shift) ^ ((fiEnable && (5198 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_25_io_in_control_0_dataflow_b <=( _mesh_30_25_io_out_control_0_dataflow) ^ ((fiEnable && (5199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_25_io_in_control_0_propagate_b <=( _mesh_30_25_io_out_control_0_propagate) ^ ((fiEnable && (5200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_26_0) begin
			b_832_0 <=( io_in_b_26_0) ^ ((fiEnable && (5201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1856_0 <=( io_in_d_26_0) ^ ((fiEnable && (5202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_26_io_in_control_0_shift_b <=( io_in_control_26_0_shift) ^ ((fiEnable && (5203 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_26_io_in_control_0_dataflow_b <=( io_in_control_26_0_dataflow) ^ ((fiEnable && (5204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_26_io_in_control_0_propagate_b <=( io_in_control_26_0_propagate) ^ ((fiEnable && (5205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_26_io_out_valid_0) begin
			b_833_0 <=( _mesh_0_26_io_out_b_0) ^ ((fiEnable && (5206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1857_0 <=( _mesh_0_26_io_out_c_0) ^ ((fiEnable && (5207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_26_io_in_control_0_shift_b <=( _mesh_0_26_io_out_control_0_shift) ^ ((fiEnable && (5208 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_26_io_in_control_0_dataflow_b <=( _mesh_0_26_io_out_control_0_dataflow) ^ ((fiEnable && (5209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_26_io_in_control_0_propagate_b <=( _mesh_0_26_io_out_control_0_propagate) ^ ((fiEnable && (5210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_26_io_out_valid_0) begin
			b_834_0 <=( _mesh_1_26_io_out_b_0) ^ ((fiEnable && (5211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1858_0 <=( _mesh_1_26_io_out_c_0) ^ ((fiEnable && (5212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_26_io_in_control_0_shift_b <=( _mesh_1_26_io_out_control_0_shift) ^ ((fiEnable && (5213 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_26_io_in_control_0_dataflow_b <=( _mesh_1_26_io_out_control_0_dataflow) ^ ((fiEnable && (5214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_26_io_in_control_0_propagate_b <=( _mesh_1_26_io_out_control_0_propagate) ^ ((fiEnable && (5215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_26_io_out_valid_0) begin
			b_835_0 <=( _mesh_2_26_io_out_b_0) ^ ((fiEnable && (5216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1859_0 <=( _mesh_2_26_io_out_c_0) ^ ((fiEnable && (5217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_26_io_in_control_0_shift_b <=( _mesh_2_26_io_out_control_0_shift) ^ ((fiEnable && (5218 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_26_io_in_control_0_dataflow_b <=( _mesh_2_26_io_out_control_0_dataflow) ^ ((fiEnable && (5219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_26_io_in_control_0_propagate_b <=( _mesh_2_26_io_out_control_0_propagate) ^ ((fiEnable && (5220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_26_io_out_valid_0) begin
			b_836_0 <=( _mesh_3_26_io_out_b_0) ^ ((fiEnable && (5221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1860_0 <=( _mesh_3_26_io_out_c_0) ^ ((fiEnable && (5222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_26_io_in_control_0_shift_b <=( _mesh_3_26_io_out_control_0_shift) ^ ((fiEnable && (5223 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_26_io_in_control_0_dataflow_b <=( _mesh_3_26_io_out_control_0_dataflow) ^ ((fiEnable && (5224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_26_io_in_control_0_propagate_b <=( _mesh_3_26_io_out_control_0_propagate) ^ ((fiEnable && (5225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_26_io_out_valid_0) begin
			b_837_0 <=( _mesh_4_26_io_out_b_0) ^ ((fiEnable && (5226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1861_0 <=( _mesh_4_26_io_out_c_0) ^ ((fiEnable && (5227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_26_io_in_control_0_shift_b <=( _mesh_4_26_io_out_control_0_shift) ^ ((fiEnable && (5228 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_26_io_in_control_0_dataflow_b <=( _mesh_4_26_io_out_control_0_dataflow) ^ ((fiEnable && (5229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_26_io_in_control_0_propagate_b <=( _mesh_4_26_io_out_control_0_propagate) ^ ((fiEnable && (5230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_26_io_out_valid_0) begin
			b_838_0 <=( _mesh_5_26_io_out_b_0) ^ ((fiEnable && (5231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1862_0 <=( _mesh_5_26_io_out_c_0) ^ ((fiEnable && (5232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_26_io_in_control_0_shift_b <=( _mesh_5_26_io_out_control_0_shift) ^ ((fiEnable && (5233 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_26_io_in_control_0_dataflow_b <=( _mesh_5_26_io_out_control_0_dataflow) ^ ((fiEnable && (5234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_26_io_in_control_0_propagate_b <=( _mesh_5_26_io_out_control_0_propagate) ^ ((fiEnable && (5235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_26_io_out_valid_0) begin
			b_839_0 <=( _mesh_6_26_io_out_b_0) ^ ((fiEnable && (5236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1863_0 <=( _mesh_6_26_io_out_c_0) ^ ((fiEnable && (5237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_26_io_in_control_0_shift_b <=( _mesh_6_26_io_out_control_0_shift) ^ ((fiEnable && (5238 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_26_io_in_control_0_dataflow_b <=( _mesh_6_26_io_out_control_0_dataflow) ^ ((fiEnable && (5239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_26_io_in_control_0_propagate_b <=( _mesh_6_26_io_out_control_0_propagate) ^ ((fiEnable && (5240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_26_io_out_valid_0) begin
			b_840_0 <=( _mesh_7_26_io_out_b_0) ^ ((fiEnable && (5241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1864_0 <=( _mesh_7_26_io_out_c_0) ^ ((fiEnable && (5242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_26_io_in_control_0_shift_b <=( _mesh_7_26_io_out_control_0_shift) ^ ((fiEnable && (5243 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_26_io_in_control_0_dataflow_b <=( _mesh_7_26_io_out_control_0_dataflow) ^ ((fiEnable && (5244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_26_io_in_control_0_propagate_b <=( _mesh_7_26_io_out_control_0_propagate) ^ ((fiEnable && (5245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_26_io_out_valid_0) begin
			b_841_0 <=( _mesh_8_26_io_out_b_0) ^ ((fiEnable && (5246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1865_0 <=( _mesh_8_26_io_out_c_0) ^ ((fiEnable && (5247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_26_io_in_control_0_shift_b <=( _mesh_8_26_io_out_control_0_shift) ^ ((fiEnable && (5248 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_26_io_in_control_0_dataflow_b <=( _mesh_8_26_io_out_control_0_dataflow) ^ ((fiEnable && (5249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_26_io_in_control_0_propagate_b <=( _mesh_8_26_io_out_control_0_propagate) ^ ((fiEnable && (5250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_26_io_out_valid_0) begin
			b_842_0 <=( _mesh_9_26_io_out_b_0) ^ ((fiEnable && (5251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1866_0 <=( _mesh_9_26_io_out_c_0) ^ ((fiEnable && (5252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_26_io_in_control_0_shift_b <=( _mesh_9_26_io_out_control_0_shift) ^ ((fiEnable && (5253 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_26_io_in_control_0_dataflow_b <=( _mesh_9_26_io_out_control_0_dataflow) ^ ((fiEnable && (5254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_26_io_in_control_0_propagate_b <=( _mesh_9_26_io_out_control_0_propagate) ^ ((fiEnable && (5255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_26_io_out_valid_0) begin
			b_843_0 <=( _mesh_10_26_io_out_b_0) ^ ((fiEnable && (5256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1867_0 <=( _mesh_10_26_io_out_c_0) ^ ((fiEnable && (5257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_26_io_in_control_0_shift_b <=( _mesh_10_26_io_out_control_0_shift) ^ ((fiEnable && (5258 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_26_io_in_control_0_dataflow_b <=( _mesh_10_26_io_out_control_0_dataflow) ^ ((fiEnable && (5259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_26_io_in_control_0_propagate_b <=( _mesh_10_26_io_out_control_0_propagate) ^ ((fiEnable && (5260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_26_io_out_valid_0) begin
			b_844_0 <=( _mesh_11_26_io_out_b_0) ^ ((fiEnable && (5261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1868_0 <=( _mesh_11_26_io_out_c_0) ^ ((fiEnable && (5262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_26_io_in_control_0_shift_b <=( _mesh_11_26_io_out_control_0_shift) ^ ((fiEnable && (5263 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_26_io_in_control_0_dataflow_b <=( _mesh_11_26_io_out_control_0_dataflow) ^ ((fiEnable && (5264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_26_io_in_control_0_propagate_b <=( _mesh_11_26_io_out_control_0_propagate) ^ ((fiEnable && (5265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_26_io_out_valid_0) begin
			b_845_0 <=( _mesh_12_26_io_out_b_0) ^ ((fiEnable && (5266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1869_0 <=( _mesh_12_26_io_out_c_0) ^ ((fiEnable && (5267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_26_io_in_control_0_shift_b <=( _mesh_12_26_io_out_control_0_shift) ^ ((fiEnable && (5268 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_26_io_in_control_0_dataflow_b <=( _mesh_12_26_io_out_control_0_dataflow) ^ ((fiEnable && (5269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_26_io_in_control_0_propagate_b <=( _mesh_12_26_io_out_control_0_propagate) ^ ((fiEnable && (5270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_26_io_out_valid_0) begin
			b_846_0 <=( _mesh_13_26_io_out_b_0) ^ ((fiEnable && (5271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1870_0 <=( _mesh_13_26_io_out_c_0) ^ ((fiEnable && (5272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_26_io_in_control_0_shift_b <=( _mesh_13_26_io_out_control_0_shift) ^ ((fiEnable && (5273 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_26_io_in_control_0_dataflow_b <=( _mesh_13_26_io_out_control_0_dataflow) ^ ((fiEnable && (5274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_26_io_in_control_0_propagate_b <=( _mesh_13_26_io_out_control_0_propagate) ^ ((fiEnable && (5275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_26_io_out_valid_0) begin
			b_847_0 <=( _mesh_14_26_io_out_b_0) ^ ((fiEnable && (5276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1871_0 <=( _mesh_14_26_io_out_c_0) ^ ((fiEnable && (5277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_26_io_in_control_0_shift_b <=( _mesh_14_26_io_out_control_0_shift) ^ ((fiEnable && (5278 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_26_io_in_control_0_dataflow_b <=( _mesh_14_26_io_out_control_0_dataflow) ^ ((fiEnable && (5279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_26_io_in_control_0_propagate_b <=( _mesh_14_26_io_out_control_0_propagate) ^ ((fiEnable && (5280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_26_io_out_valid_0) begin
			b_848_0 <=( _mesh_15_26_io_out_b_0) ^ ((fiEnable && (5281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1872_0 <=( _mesh_15_26_io_out_c_0) ^ ((fiEnable && (5282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_26_io_in_control_0_shift_b <=( _mesh_15_26_io_out_control_0_shift) ^ ((fiEnable && (5283 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_26_io_in_control_0_dataflow_b <=( _mesh_15_26_io_out_control_0_dataflow) ^ ((fiEnable && (5284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_26_io_in_control_0_propagate_b <=( _mesh_15_26_io_out_control_0_propagate) ^ ((fiEnable && (5285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_26_io_out_valid_0) begin
			b_849_0 <=( _mesh_16_26_io_out_b_0) ^ ((fiEnable && (5286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1873_0 <=( _mesh_16_26_io_out_c_0) ^ ((fiEnable && (5287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_26_io_in_control_0_shift_b <=( _mesh_16_26_io_out_control_0_shift) ^ ((fiEnable && (5288 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_26_io_in_control_0_dataflow_b <=( _mesh_16_26_io_out_control_0_dataflow) ^ ((fiEnable && (5289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_26_io_in_control_0_propagate_b <=( _mesh_16_26_io_out_control_0_propagate) ^ ((fiEnable && (5290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_26_io_out_valid_0) begin
			b_850_0 <=( _mesh_17_26_io_out_b_0) ^ ((fiEnable && (5291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1874_0 <=( _mesh_17_26_io_out_c_0) ^ ((fiEnable && (5292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_26_io_in_control_0_shift_b <=( _mesh_17_26_io_out_control_0_shift) ^ ((fiEnable && (5293 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_26_io_in_control_0_dataflow_b <=( _mesh_17_26_io_out_control_0_dataflow) ^ ((fiEnable && (5294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_26_io_in_control_0_propagate_b <=( _mesh_17_26_io_out_control_0_propagate) ^ ((fiEnable && (5295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_26_io_out_valid_0) begin
			b_851_0 <=( _mesh_18_26_io_out_b_0) ^ ((fiEnable && (5296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1875_0 <=( _mesh_18_26_io_out_c_0) ^ ((fiEnable && (5297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_26_io_in_control_0_shift_b <=( _mesh_18_26_io_out_control_0_shift) ^ ((fiEnable && (5298 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_26_io_in_control_0_dataflow_b <=( _mesh_18_26_io_out_control_0_dataflow) ^ ((fiEnable && (5299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_26_io_in_control_0_propagate_b <=( _mesh_18_26_io_out_control_0_propagate) ^ ((fiEnable && (5300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_26_io_out_valid_0) begin
			b_852_0 <=( _mesh_19_26_io_out_b_0) ^ ((fiEnable && (5301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1876_0 <=( _mesh_19_26_io_out_c_0) ^ ((fiEnable && (5302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_26_io_in_control_0_shift_b <=( _mesh_19_26_io_out_control_0_shift) ^ ((fiEnable && (5303 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_26_io_in_control_0_dataflow_b <=( _mesh_19_26_io_out_control_0_dataflow) ^ ((fiEnable && (5304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_26_io_in_control_0_propagate_b <=( _mesh_19_26_io_out_control_0_propagate) ^ ((fiEnable && (5305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_26_io_out_valid_0) begin
			b_853_0 <=( _mesh_20_26_io_out_b_0) ^ ((fiEnable && (5306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1877_0 <=( _mesh_20_26_io_out_c_0) ^ ((fiEnable && (5307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_26_io_in_control_0_shift_b <=( _mesh_20_26_io_out_control_0_shift) ^ ((fiEnable && (5308 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_26_io_in_control_0_dataflow_b <=( _mesh_20_26_io_out_control_0_dataflow) ^ ((fiEnable && (5309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_26_io_in_control_0_propagate_b <=( _mesh_20_26_io_out_control_0_propagate) ^ ((fiEnable && (5310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_26_io_out_valid_0) begin
			b_854_0 <=( _mesh_21_26_io_out_b_0) ^ ((fiEnable && (5311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1878_0 <=( _mesh_21_26_io_out_c_0) ^ ((fiEnable && (5312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_26_io_in_control_0_shift_b <=( _mesh_21_26_io_out_control_0_shift) ^ ((fiEnable && (5313 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_26_io_in_control_0_dataflow_b <=( _mesh_21_26_io_out_control_0_dataflow) ^ ((fiEnable && (5314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_26_io_in_control_0_propagate_b <=( _mesh_21_26_io_out_control_0_propagate) ^ ((fiEnable && (5315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_26_io_out_valid_0) begin
			b_855_0 <=( _mesh_22_26_io_out_b_0) ^ ((fiEnable && (5316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1879_0 <=( _mesh_22_26_io_out_c_0) ^ ((fiEnable && (5317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_26_io_in_control_0_shift_b <=( _mesh_22_26_io_out_control_0_shift) ^ ((fiEnable && (5318 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_26_io_in_control_0_dataflow_b <=( _mesh_22_26_io_out_control_0_dataflow) ^ ((fiEnable && (5319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_26_io_in_control_0_propagate_b <=( _mesh_22_26_io_out_control_0_propagate) ^ ((fiEnable && (5320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_26_io_out_valid_0) begin
			b_856_0 <=( _mesh_23_26_io_out_b_0) ^ ((fiEnable && (5321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1880_0 <=( _mesh_23_26_io_out_c_0) ^ ((fiEnable && (5322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_26_io_in_control_0_shift_b <=( _mesh_23_26_io_out_control_0_shift) ^ ((fiEnable && (5323 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_26_io_in_control_0_dataflow_b <=( _mesh_23_26_io_out_control_0_dataflow) ^ ((fiEnable && (5324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_26_io_in_control_0_propagate_b <=( _mesh_23_26_io_out_control_0_propagate) ^ ((fiEnable && (5325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_26_io_out_valid_0) begin
			b_857_0 <=( _mesh_24_26_io_out_b_0) ^ ((fiEnable && (5326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1881_0 <=( _mesh_24_26_io_out_c_0) ^ ((fiEnable && (5327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_26_io_in_control_0_shift_b <=( _mesh_24_26_io_out_control_0_shift) ^ ((fiEnable && (5328 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_26_io_in_control_0_dataflow_b <=( _mesh_24_26_io_out_control_0_dataflow) ^ ((fiEnable && (5329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_26_io_in_control_0_propagate_b <=( _mesh_24_26_io_out_control_0_propagate) ^ ((fiEnable && (5330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_26_io_out_valid_0) begin
			b_858_0 <=( _mesh_25_26_io_out_b_0) ^ ((fiEnable && (5331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1882_0 <=( _mesh_25_26_io_out_c_0) ^ ((fiEnable && (5332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_26_io_in_control_0_shift_b <=( _mesh_25_26_io_out_control_0_shift) ^ ((fiEnable && (5333 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_26_io_in_control_0_dataflow_b <=( _mesh_25_26_io_out_control_0_dataflow) ^ ((fiEnable && (5334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_26_io_in_control_0_propagate_b <=( _mesh_25_26_io_out_control_0_propagate) ^ ((fiEnable && (5335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_26_io_out_valid_0) begin
			b_859_0 <=( _mesh_26_26_io_out_b_0) ^ ((fiEnable && (5336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1883_0 <=( _mesh_26_26_io_out_c_0) ^ ((fiEnable && (5337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_26_io_in_control_0_shift_b <=( _mesh_26_26_io_out_control_0_shift) ^ ((fiEnable && (5338 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_26_io_in_control_0_dataflow_b <=( _mesh_26_26_io_out_control_0_dataflow) ^ ((fiEnable && (5339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_26_io_in_control_0_propagate_b <=( _mesh_26_26_io_out_control_0_propagate) ^ ((fiEnable && (5340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_26_io_out_valid_0) begin
			b_860_0 <=( _mesh_27_26_io_out_b_0) ^ ((fiEnable && (5341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1884_0 <=( _mesh_27_26_io_out_c_0) ^ ((fiEnable && (5342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_26_io_in_control_0_shift_b <=( _mesh_27_26_io_out_control_0_shift) ^ ((fiEnable && (5343 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_26_io_in_control_0_dataflow_b <=( _mesh_27_26_io_out_control_0_dataflow) ^ ((fiEnable && (5344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_26_io_in_control_0_propagate_b <=( _mesh_27_26_io_out_control_0_propagate) ^ ((fiEnable && (5345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_26_io_out_valid_0) begin
			b_861_0 <=( _mesh_28_26_io_out_b_0) ^ ((fiEnable && (5346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1885_0 <=( _mesh_28_26_io_out_c_0) ^ ((fiEnable && (5347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_26_io_in_control_0_shift_b <=( _mesh_28_26_io_out_control_0_shift) ^ ((fiEnable && (5348 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_26_io_in_control_0_dataflow_b <=( _mesh_28_26_io_out_control_0_dataflow) ^ ((fiEnable && (5349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_26_io_in_control_0_propagate_b <=( _mesh_28_26_io_out_control_0_propagate) ^ ((fiEnable && (5350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_26_io_out_valid_0) begin
			b_862_0 <=( _mesh_29_26_io_out_b_0) ^ ((fiEnable && (5351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1886_0 <=( _mesh_29_26_io_out_c_0) ^ ((fiEnable && (5352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_26_io_in_control_0_shift_b <=( _mesh_29_26_io_out_control_0_shift) ^ ((fiEnable && (5353 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_26_io_in_control_0_dataflow_b <=( _mesh_29_26_io_out_control_0_dataflow) ^ ((fiEnable && (5354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_26_io_in_control_0_propagate_b <=( _mesh_29_26_io_out_control_0_propagate) ^ ((fiEnable && (5355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_26_io_out_valid_0) begin
			b_863_0 <=( _mesh_30_26_io_out_b_0) ^ ((fiEnable && (5356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1887_0 <=( _mesh_30_26_io_out_c_0) ^ ((fiEnable && (5357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_26_io_in_control_0_shift_b <=( _mesh_30_26_io_out_control_0_shift) ^ ((fiEnable && (5358 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_26_io_in_control_0_dataflow_b <=( _mesh_30_26_io_out_control_0_dataflow) ^ ((fiEnable && (5359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_26_io_in_control_0_propagate_b <=( _mesh_30_26_io_out_control_0_propagate) ^ ((fiEnable && (5360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_27_0) begin
			b_864_0 <=( io_in_b_27_0) ^ ((fiEnable && (5361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1888_0 <=( io_in_d_27_0) ^ ((fiEnable && (5362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_27_io_in_control_0_shift_b <=( io_in_control_27_0_shift) ^ ((fiEnable && (5363 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_27_io_in_control_0_dataflow_b <=( io_in_control_27_0_dataflow) ^ ((fiEnable && (5364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_27_io_in_control_0_propagate_b <=( io_in_control_27_0_propagate) ^ ((fiEnable && (5365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_27_io_out_valid_0) begin
			b_865_0 <=( _mesh_0_27_io_out_b_0) ^ ((fiEnable && (5366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1889_0 <=( _mesh_0_27_io_out_c_0) ^ ((fiEnable && (5367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_27_io_in_control_0_shift_b <=( _mesh_0_27_io_out_control_0_shift) ^ ((fiEnable && (5368 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_27_io_in_control_0_dataflow_b <=( _mesh_0_27_io_out_control_0_dataflow) ^ ((fiEnable && (5369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_27_io_in_control_0_propagate_b <=( _mesh_0_27_io_out_control_0_propagate) ^ ((fiEnable && (5370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_27_io_out_valid_0) begin
			b_866_0 <=( _mesh_1_27_io_out_b_0) ^ ((fiEnable && (5371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1890_0 <=( _mesh_1_27_io_out_c_0) ^ ((fiEnable && (5372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_27_io_in_control_0_shift_b <=( _mesh_1_27_io_out_control_0_shift) ^ ((fiEnable && (5373 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_27_io_in_control_0_dataflow_b <=( _mesh_1_27_io_out_control_0_dataflow) ^ ((fiEnable && (5374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_27_io_in_control_0_propagate_b <=( _mesh_1_27_io_out_control_0_propagate) ^ ((fiEnable && (5375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_27_io_out_valid_0) begin
			b_867_0 <=( _mesh_2_27_io_out_b_0) ^ ((fiEnable && (5376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1891_0 <=( _mesh_2_27_io_out_c_0) ^ ((fiEnable && (5377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_27_io_in_control_0_shift_b <=( _mesh_2_27_io_out_control_0_shift) ^ ((fiEnable && (5378 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_27_io_in_control_0_dataflow_b <=( _mesh_2_27_io_out_control_0_dataflow) ^ ((fiEnable && (5379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_27_io_in_control_0_propagate_b <=( _mesh_2_27_io_out_control_0_propagate) ^ ((fiEnable && (5380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_27_io_out_valid_0) begin
			b_868_0 <=( _mesh_3_27_io_out_b_0) ^ ((fiEnable && (5381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1892_0 <=( _mesh_3_27_io_out_c_0) ^ ((fiEnable && (5382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_27_io_in_control_0_shift_b <=( _mesh_3_27_io_out_control_0_shift) ^ ((fiEnable && (5383 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_27_io_in_control_0_dataflow_b <=( _mesh_3_27_io_out_control_0_dataflow) ^ ((fiEnable && (5384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_27_io_in_control_0_propagate_b <=( _mesh_3_27_io_out_control_0_propagate) ^ ((fiEnable && (5385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_27_io_out_valid_0) begin
			b_869_0 <=( _mesh_4_27_io_out_b_0) ^ ((fiEnable && (5386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1893_0 <=( _mesh_4_27_io_out_c_0) ^ ((fiEnable && (5387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_27_io_in_control_0_shift_b <=( _mesh_4_27_io_out_control_0_shift) ^ ((fiEnable && (5388 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_27_io_in_control_0_dataflow_b <=( _mesh_4_27_io_out_control_0_dataflow) ^ ((fiEnable && (5389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_27_io_in_control_0_propagate_b <=( _mesh_4_27_io_out_control_0_propagate) ^ ((fiEnable && (5390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_27_io_out_valid_0) begin
			b_870_0 <=( _mesh_5_27_io_out_b_0) ^ ((fiEnable && (5391 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1894_0 <=( _mesh_5_27_io_out_c_0) ^ ((fiEnable && (5392 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_27_io_in_control_0_shift_b <=( _mesh_5_27_io_out_control_0_shift) ^ ((fiEnable && (5393 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_27_io_in_control_0_dataflow_b <=( _mesh_5_27_io_out_control_0_dataflow) ^ ((fiEnable && (5394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_27_io_in_control_0_propagate_b <=( _mesh_5_27_io_out_control_0_propagate) ^ ((fiEnable && (5395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_27_io_out_valid_0) begin
			b_871_0 <=( _mesh_6_27_io_out_b_0) ^ ((fiEnable && (5396 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1895_0 <=( _mesh_6_27_io_out_c_0) ^ ((fiEnable && (5397 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_27_io_in_control_0_shift_b <=( _mesh_6_27_io_out_control_0_shift) ^ ((fiEnable && (5398 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_27_io_in_control_0_dataflow_b <=( _mesh_6_27_io_out_control_0_dataflow) ^ ((fiEnable && (5399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_27_io_in_control_0_propagate_b <=( _mesh_6_27_io_out_control_0_propagate) ^ ((fiEnable && (5400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_27_io_out_valid_0) begin
			b_872_0 <=( _mesh_7_27_io_out_b_0) ^ ((fiEnable && (5401 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1896_0 <=( _mesh_7_27_io_out_c_0) ^ ((fiEnable && (5402 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_27_io_in_control_0_shift_b <=( _mesh_7_27_io_out_control_0_shift) ^ ((fiEnable && (5403 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_27_io_in_control_0_dataflow_b <=( _mesh_7_27_io_out_control_0_dataflow) ^ ((fiEnable && (5404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_27_io_in_control_0_propagate_b <=( _mesh_7_27_io_out_control_0_propagate) ^ ((fiEnable && (5405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_27_io_out_valid_0) begin
			b_873_0 <=( _mesh_8_27_io_out_b_0) ^ ((fiEnable && (5406 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1897_0 <=( _mesh_8_27_io_out_c_0) ^ ((fiEnable && (5407 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_27_io_in_control_0_shift_b <=( _mesh_8_27_io_out_control_0_shift) ^ ((fiEnable && (5408 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_27_io_in_control_0_dataflow_b <=( _mesh_8_27_io_out_control_0_dataflow) ^ ((fiEnable && (5409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_27_io_in_control_0_propagate_b <=( _mesh_8_27_io_out_control_0_propagate) ^ ((fiEnable && (5410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_27_io_out_valid_0) begin
			b_874_0 <=( _mesh_9_27_io_out_b_0) ^ ((fiEnable && (5411 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1898_0 <=( _mesh_9_27_io_out_c_0) ^ ((fiEnable && (5412 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_27_io_in_control_0_shift_b <=( _mesh_9_27_io_out_control_0_shift) ^ ((fiEnable && (5413 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_27_io_in_control_0_dataflow_b <=( _mesh_9_27_io_out_control_0_dataflow) ^ ((fiEnable && (5414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_27_io_in_control_0_propagate_b <=( _mesh_9_27_io_out_control_0_propagate) ^ ((fiEnable && (5415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_27_io_out_valid_0) begin
			b_875_0 <=( _mesh_10_27_io_out_b_0) ^ ((fiEnable && (5416 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1899_0 <=( _mesh_10_27_io_out_c_0) ^ ((fiEnable && (5417 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_27_io_in_control_0_shift_b <=( _mesh_10_27_io_out_control_0_shift) ^ ((fiEnable && (5418 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_27_io_in_control_0_dataflow_b <=( _mesh_10_27_io_out_control_0_dataflow) ^ ((fiEnable && (5419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_27_io_in_control_0_propagate_b <=( _mesh_10_27_io_out_control_0_propagate) ^ ((fiEnable && (5420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_27_io_out_valid_0) begin
			b_876_0 <=( _mesh_11_27_io_out_b_0) ^ ((fiEnable && (5421 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1900_0 <=( _mesh_11_27_io_out_c_0) ^ ((fiEnable && (5422 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_27_io_in_control_0_shift_b <=( _mesh_11_27_io_out_control_0_shift) ^ ((fiEnable && (5423 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_27_io_in_control_0_dataflow_b <=( _mesh_11_27_io_out_control_0_dataflow) ^ ((fiEnable && (5424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_27_io_in_control_0_propagate_b <=( _mesh_11_27_io_out_control_0_propagate) ^ ((fiEnable && (5425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_27_io_out_valid_0) begin
			b_877_0 <=( _mesh_12_27_io_out_b_0) ^ ((fiEnable && (5426 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1901_0 <=( _mesh_12_27_io_out_c_0) ^ ((fiEnable && (5427 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_27_io_in_control_0_shift_b <=( _mesh_12_27_io_out_control_0_shift) ^ ((fiEnable && (5428 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_27_io_in_control_0_dataflow_b <=( _mesh_12_27_io_out_control_0_dataflow) ^ ((fiEnable && (5429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_27_io_in_control_0_propagate_b <=( _mesh_12_27_io_out_control_0_propagate) ^ ((fiEnable && (5430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_27_io_out_valid_0) begin
			b_878_0 <=( _mesh_13_27_io_out_b_0) ^ ((fiEnable && (5431 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1902_0 <=( _mesh_13_27_io_out_c_0) ^ ((fiEnable && (5432 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_27_io_in_control_0_shift_b <=( _mesh_13_27_io_out_control_0_shift) ^ ((fiEnable && (5433 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_27_io_in_control_0_dataflow_b <=( _mesh_13_27_io_out_control_0_dataflow) ^ ((fiEnable && (5434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_27_io_in_control_0_propagate_b <=( _mesh_13_27_io_out_control_0_propagate) ^ ((fiEnable && (5435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_27_io_out_valid_0) begin
			b_879_0 <=( _mesh_14_27_io_out_b_0) ^ ((fiEnable && (5436 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1903_0 <=( _mesh_14_27_io_out_c_0) ^ ((fiEnable && (5437 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_27_io_in_control_0_shift_b <=( _mesh_14_27_io_out_control_0_shift) ^ ((fiEnable && (5438 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_27_io_in_control_0_dataflow_b <=( _mesh_14_27_io_out_control_0_dataflow) ^ ((fiEnable && (5439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_27_io_in_control_0_propagate_b <=( _mesh_14_27_io_out_control_0_propagate) ^ ((fiEnable && (5440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_27_io_out_valid_0) begin
			b_880_0 <=( _mesh_15_27_io_out_b_0) ^ ((fiEnable && (5441 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1904_0 <=( _mesh_15_27_io_out_c_0) ^ ((fiEnable && (5442 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_27_io_in_control_0_shift_b <=( _mesh_15_27_io_out_control_0_shift) ^ ((fiEnable && (5443 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_27_io_in_control_0_dataflow_b <=( _mesh_15_27_io_out_control_0_dataflow) ^ ((fiEnable && (5444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_27_io_in_control_0_propagate_b <=( _mesh_15_27_io_out_control_0_propagate) ^ ((fiEnable && (5445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_27_io_out_valid_0) begin
			b_881_0 <=( _mesh_16_27_io_out_b_0) ^ ((fiEnable && (5446 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1905_0 <=( _mesh_16_27_io_out_c_0) ^ ((fiEnable && (5447 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_27_io_in_control_0_shift_b <=( _mesh_16_27_io_out_control_0_shift) ^ ((fiEnable && (5448 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_27_io_in_control_0_dataflow_b <=( _mesh_16_27_io_out_control_0_dataflow) ^ ((fiEnable && (5449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_27_io_in_control_0_propagate_b <=( _mesh_16_27_io_out_control_0_propagate) ^ ((fiEnable && (5450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_27_io_out_valid_0) begin
			b_882_0 <=( _mesh_17_27_io_out_b_0) ^ ((fiEnable && (5451 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1906_0 <=( _mesh_17_27_io_out_c_0) ^ ((fiEnable && (5452 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_27_io_in_control_0_shift_b <=( _mesh_17_27_io_out_control_0_shift) ^ ((fiEnable && (5453 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_27_io_in_control_0_dataflow_b <=( _mesh_17_27_io_out_control_0_dataflow) ^ ((fiEnable && (5454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_27_io_in_control_0_propagate_b <=( _mesh_17_27_io_out_control_0_propagate) ^ ((fiEnable && (5455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_27_io_out_valid_0) begin
			b_883_0 <=( _mesh_18_27_io_out_b_0) ^ ((fiEnable && (5456 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1907_0 <=( _mesh_18_27_io_out_c_0) ^ ((fiEnable && (5457 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_27_io_in_control_0_shift_b <=( _mesh_18_27_io_out_control_0_shift) ^ ((fiEnable && (5458 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_27_io_in_control_0_dataflow_b <=( _mesh_18_27_io_out_control_0_dataflow) ^ ((fiEnable && (5459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_27_io_in_control_0_propagate_b <=( _mesh_18_27_io_out_control_0_propagate) ^ ((fiEnable && (5460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_27_io_out_valid_0) begin
			b_884_0 <=( _mesh_19_27_io_out_b_0) ^ ((fiEnable && (5461 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1908_0 <=( _mesh_19_27_io_out_c_0) ^ ((fiEnable && (5462 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_27_io_in_control_0_shift_b <=( _mesh_19_27_io_out_control_0_shift) ^ ((fiEnable && (5463 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_27_io_in_control_0_dataflow_b <=( _mesh_19_27_io_out_control_0_dataflow) ^ ((fiEnable && (5464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_27_io_in_control_0_propagate_b <=( _mesh_19_27_io_out_control_0_propagate) ^ ((fiEnable && (5465 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_27_io_out_valid_0) begin
			b_885_0 <=( _mesh_20_27_io_out_b_0) ^ ((fiEnable && (5466 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1909_0 <=( _mesh_20_27_io_out_c_0) ^ ((fiEnable && (5467 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_27_io_in_control_0_shift_b <=( _mesh_20_27_io_out_control_0_shift) ^ ((fiEnable && (5468 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_27_io_in_control_0_dataflow_b <=( _mesh_20_27_io_out_control_0_dataflow) ^ ((fiEnable && (5469 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_27_io_in_control_0_propagate_b <=( _mesh_20_27_io_out_control_0_propagate) ^ ((fiEnable && (5470 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_27_io_out_valid_0) begin
			b_886_0 <=( _mesh_21_27_io_out_b_0) ^ ((fiEnable && (5471 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1910_0 <=( _mesh_21_27_io_out_c_0) ^ ((fiEnable && (5472 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_27_io_in_control_0_shift_b <=( _mesh_21_27_io_out_control_0_shift) ^ ((fiEnable && (5473 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_27_io_in_control_0_dataflow_b <=( _mesh_21_27_io_out_control_0_dataflow) ^ ((fiEnable && (5474 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_27_io_in_control_0_propagate_b <=( _mesh_21_27_io_out_control_0_propagate) ^ ((fiEnable && (5475 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_27_io_out_valid_0) begin
			b_887_0 <=( _mesh_22_27_io_out_b_0) ^ ((fiEnable && (5476 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1911_0 <=( _mesh_22_27_io_out_c_0) ^ ((fiEnable && (5477 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_27_io_in_control_0_shift_b <=( _mesh_22_27_io_out_control_0_shift) ^ ((fiEnable && (5478 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_27_io_in_control_0_dataflow_b <=( _mesh_22_27_io_out_control_0_dataflow) ^ ((fiEnable && (5479 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_27_io_in_control_0_propagate_b <=( _mesh_22_27_io_out_control_0_propagate) ^ ((fiEnable && (5480 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_27_io_out_valid_0) begin
			b_888_0 <=( _mesh_23_27_io_out_b_0) ^ ((fiEnable && (5481 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1912_0 <=( _mesh_23_27_io_out_c_0) ^ ((fiEnable && (5482 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_27_io_in_control_0_shift_b <=( _mesh_23_27_io_out_control_0_shift) ^ ((fiEnable && (5483 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_27_io_in_control_0_dataflow_b <=( _mesh_23_27_io_out_control_0_dataflow) ^ ((fiEnable && (5484 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_27_io_in_control_0_propagate_b <=( _mesh_23_27_io_out_control_0_propagate) ^ ((fiEnable && (5485 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_27_io_out_valid_0) begin
			b_889_0 <=( _mesh_24_27_io_out_b_0) ^ ((fiEnable && (5486 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1913_0 <=( _mesh_24_27_io_out_c_0) ^ ((fiEnable && (5487 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_27_io_in_control_0_shift_b <=( _mesh_24_27_io_out_control_0_shift) ^ ((fiEnable && (5488 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_27_io_in_control_0_dataflow_b <=( _mesh_24_27_io_out_control_0_dataflow) ^ ((fiEnable && (5489 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_27_io_in_control_0_propagate_b <=( _mesh_24_27_io_out_control_0_propagate) ^ ((fiEnable && (5490 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_27_io_out_valid_0) begin
			b_890_0 <=( _mesh_25_27_io_out_b_0) ^ ((fiEnable && (5491 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1914_0 <=( _mesh_25_27_io_out_c_0) ^ ((fiEnable && (5492 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_27_io_in_control_0_shift_b <=( _mesh_25_27_io_out_control_0_shift) ^ ((fiEnable && (5493 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_27_io_in_control_0_dataflow_b <=( _mesh_25_27_io_out_control_0_dataflow) ^ ((fiEnable && (5494 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_27_io_in_control_0_propagate_b <=( _mesh_25_27_io_out_control_0_propagate) ^ ((fiEnable && (5495 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_27_io_out_valid_0) begin
			b_891_0 <=( _mesh_26_27_io_out_b_0) ^ ((fiEnable && (5496 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1915_0 <=( _mesh_26_27_io_out_c_0) ^ ((fiEnable && (5497 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_27_io_in_control_0_shift_b <=( _mesh_26_27_io_out_control_0_shift) ^ ((fiEnable && (5498 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_27_io_in_control_0_dataflow_b <=( _mesh_26_27_io_out_control_0_dataflow) ^ ((fiEnable && (5499 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_27_io_in_control_0_propagate_b <=( _mesh_26_27_io_out_control_0_propagate) ^ ((fiEnable && (5500 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_27_io_out_valid_0) begin
			b_892_0 <=( _mesh_27_27_io_out_b_0) ^ ((fiEnable && (5501 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1916_0 <=( _mesh_27_27_io_out_c_0) ^ ((fiEnable && (5502 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_27_io_in_control_0_shift_b <=( _mesh_27_27_io_out_control_0_shift) ^ ((fiEnable && (5503 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_27_io_in_control_0_dataflow_b <=( _mesh_27_27_io_out_control_0_dataflow) ^ ((fiEnable && (5504 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_27_io_in_control_0_propagate_b <=( _mesh_27_27_io_out_control_0_propagate) ^ ((fiEnable && (5505 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_27_io_out_valid_0) begin
			b_893_0 <=( _mesh_28_27_io_out_b_0) ^ ((fiEnable && (5506 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1917_0 <=( _mesh_28_27_io_out_c_0) ^ ((fiEnable && (5507 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_27_io_in_control_0_shift_b <=( _mesh_28_27_io_out_control_0_shift) ^ ((fiEnable && (5508 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_27_io_in_control_0_dataflow_b <=( _mesh_28_27_io_out_control_0_dataflow) ^ ((fiEnable && (5509 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_27_io_in_control_0_propagate_b <=( _mesh_28_27_io_out_control_0_propagate) ^ ((fiEnable && (5510 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_27_io_out_valid_0) begin
			b_894_0 <=( _mesh_29_27_io_out_b_0) ^ ((fiEnable && (5511 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1918_0 <=( _mesh_29_27_io_out_c_0) ^ ((fiEnable && (5512 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_27_io_in_control_0_shift_b <=( _mesh_29_27_io_out_control_0_shift) ^ ((fiEnable && (5513 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_27_io_in_control_0_dataflow_b <=( _mesh_29_27_io_out_control_0_dataflow) ^ ((fiEnable && (5514 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_27_io_in_control_0_propagate_b <=( _mesh_29_27_io_out_control_0_propagate) ^ ((fiEnable && (5515 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_27_io_out_valid_0) begin
			b_895_0 <=( _mesh_30_27_io_out_b_0) ^ ((fiEnable && (5516 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1919_0 <=( _mesh_30_27_io_out_c_0) ^ ((fiEnable && (5517 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_27_io_in_control_0_shift_b <=( _mesh_30_27_io_out_control_0_shift) ^ ((fiEnable && (5518 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_27_io_in_control_0_dataflow_b <=( _mesh_30_27_io_out_control_0_dataflow) ^ ((fiEnable && (5519 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_27_io_in_control_0_propagate_b <=( _mesh_30_27_io_out_control_0_propagate) ^ ((fiEnable && (5520 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_28_0) begin
			b_896_0 <=( io_in_b_28_0) ^ ((fiEnable && (5521 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1920_0 <=( io_in_d_28_0) ^ ((fiEnable && (5522 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_28_io_in_control_0_shift_b <=( io_in_control_28_0_shift) ^ ((fiEnable && (5523 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_28_io_in_control_0_dataflow_b <=( io_in_control_28_0_dataflow) ^ ((fiEnable && (5524 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_28_io_in_control_0_propagate_b <=( io_in_control_28_0_propagate) ^ ((fiEnable && (5525 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_28_io_out_valid_0) begin
			b_897_0 <=( _mesh_0_28_io_out_b_0) ^ ((fiEnable && (5526 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1921_0 <=( _mesh_0_28_io_out_c_0) ^ ((fiEnable && (5527 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_28_io_in_control_0_shift_b <=( _mesh_0_28_io_out_control_0_shift) ^ ((fiEnable && (5528 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_28_io_in_control_0_dataflow_b <=( _mesh_0_28_io_out_control_0_dataflow) ^ ((fiEnable && (5529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_28_io_in_control_0_propagate_b <=( _mesh_0_28_io_out_control_0_propagate) ^ ((fiEnable && (5530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_28_io_out_valid_0) begin
			b_898_0 <=( _mesh_1_28_io_out_b_0) ^ ((fiEnable && (5531 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1922_0 <=( _mesh_1_28_io_out_c_0) ^ ((fiEnable && (5532 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_28_io_in_control_0_shift_b <=( _mesh_1_28_io_out_control_0_shift) ^ ((fiEnable && (5533 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_28_io_in_control_0_dataflow_b <=( _mesh_1_28_io_out_control_0_dataflow) ^ ((fiEnable && (5534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_28_io_in_control_0_propagate_b <=( _mesh_1_28_io_out_control_0_propagate) ^ ((fiEnable && (5535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_28_io_out_valid_0) begin
			b_899_0 <=( _mesh_2_28_io_out_b_0) ^ ((fiEnable && (5536 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1923_0 <=( _mesh_2_28_io_out_c_0) ^ ((fiEnable && (5537 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_28_io_in_control_0_shift_b <=( _mesh_2_28_io_out_control_0_shift) ^ ((fiEnable && (5538 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_28_io_in_control_0_dataflow_b <=( _mesh_2_28_io_out_control_0_dataflow) ^ ((fiEnable && (5539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_28_io_in_control_0_propagate_b <=( _mesh_2_28_io_out_control_0_propagate) ^ ((fiEnable && (5540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_28_io_out_valid_0) begin
			b_900_0 <=( _mesh_3_28_io_out_b_0) ^ ((fiEnable && (5541 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1924_0 <=( _mesh_3_28_io_out_c_0) ^ ((fiEnable && (5542 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_28_io_in_control_0_shift_b <=( _mesh_3_28_io_out_control_0_shift) ^ ((fiEnable && (5543 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_28_io_in_control_0_dataflow_b <=( _mesh_3_28_io_out_control_0_dataflow) ^ ((fiEnable && (5544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_28_io_in_control_0_propagate_b <=( _mesh_3_28_io_out_control_0_propagate) ^ ((fiEnable && (5545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_28_io_out_valid_0) begin
			b_901_0 <=( _mesh_4_28_io_out_b_0) ^ ((fiEnable && (5546 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1925_0 <=( _mesh_4_28_io_out_c_0) ^ ((fiEnable && (5547 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_28_io_in_control_0_shift_b <=( _mesh_4_28_io_out_control_0_shift) ^ ((fiEnable && (5548 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_28_io_in_control_0_dataflow_b <=( _mesh_4_28_io_out_control_0_dataflow) ^ ((fiEnable && (5549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_28_io_in_control_0_propagate_b <=( _mesh_4_28_io_out_control_0_propagate) ^ ((fiEnable && (5550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_28_io_out_valid_0) begin
			b_902_0 <=( _mesh_5_28_io_out_b_0) ^ ((fiEnable && (5551 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1926_0 <=( _mesh_5_28_io_out_c_0) ^ ((fiEnable && (5552 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_28_io_in_control_0_shift_b <=( _mesh_5_28_io_out_control_0_shift) ^ ((fiEnable && (5553 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_28_io_in_control_0_dataflow_b <=( _mesh_5_28_io_out_control_0_dataflow) ^ ((fiEnable && (5554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_28_io_in_control_0_propagate_b <=( _mesh_5_28_io_out_control_0_propagate) ^ ((fiEnable && (5555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_28_io_out_valid_0) begin
			b_903_0 <=( _mesh_6_28_io_out_b_0) ^ ((fiEnable && (5556 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1927_0 <=( _mesh_6_28_io_out_c_0) ^ ((fiEnable && (5557 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_28_io_in_control_0_shift_b <=( _mesh_6_28_io_out_control_0_shift) ^ ((fiEnable && (5558 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_28_io_in_control_0_dataflow_b <=( _mesh_6_28_io_out_control_0_dataflow) ^ ((fiEnable && (5559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_28_io_in_control_0_propagate_b <=( _mesh_6_28_io_out_control_0_propagate) ^ ((fiEnable && (5560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_28_io_out_valid_0) begin
			b_904_0 <=( _mesh_7_28_io_out_b_0) ^ ((fiEnable && (5561 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1928_0 <=( _mesh_7_28_io_out_c_0) ^ ((fiEnable && (5562 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_28_io_in_control_0_shift_b <=( _mesh_7_28_io_out_control_0_shift) ^ ((fiEnable && (5563 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_28_io_in_control_0_dataflow_b <=( _mesh_7_28_io_out_control_0_dataflow) ^ ((fiEnable && (5564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_28_io_in_control_0_propagate_b <=( _mesh_7_28_io_out_control_0_propagate) ^ ((fiEnable && (5565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_28_io_out_valid_0) begin
			b_905_0 <=( _mesh_8_28_io_out_b_0) ^ ((fiEnable && (5566 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1929_0 <=( _mesh_8_28_io_out_c_0) ^ ((fiEnable && (5567 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_28_io_in_control_0_shift_b <=( _mesh_8_28_io_out_control_0_shift) ^ ((fiEnable && (5568 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_28_io_in_control_0_dataflow_b <=( _mesh_8_28_io_out_control_0_dataflow) ^ ((fiEnable && (5569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_28_io_in_control_0_propagate_b <=( _mesh_8_28_io_out_control_0_propagate) ^ ((fiEnable && (5570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_28_io_out_valid_0) begin
			b_906_0 <=( _mesh_9_28_io_out_b_0) ^ ((fiEnable && (5571 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1930_0 <=( _mesh_9_28_io_out_c_0) ^ ((fiEnable && (5572 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_28_io_in_control_0_shift_b <=( _mesh_9_28_io_out_control_0_shift) ^ ((fiEnable && (5573 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_28_io_in_control_0_dataflow_b <=( _mesh_9_28_io_out_control_0_dataflow) ^ ((fiEnable && (5574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_28_io_in_control_0_propagate_b <=( _mesh_9_28_io_out_control_0_propagate) ^ ((fiEnable && (5575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_28_io_out_valid_0) begin
			b_907_0 <=( _mesh_10_28_io_out_b_0) ^ ((fiEnable && (5576 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1931_0 <=( _mesh_10_28_io_out_c_0) ^ ((fiEnable && (5577 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_28_io_in_control_0_shift_b <=( _mesh_10_28_io_out_control_0_shift) ^ ((fiEnable && (5578 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_28_io_in_control_0_dataflow_b <=( _mesh_10_28_io_out_control_0_dataflow) ^ ((fiEnable && (5579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_28_io_in_control_0_propagate_b <=( _mesh_10_28_io_out_control_0_propagate) ^ ((fiEnable && (5580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_28_io_out_valid_0) begin
			b_908_0 <=( _mesh_11_28_io_out_b_0) ^ ((fiEnable && (5581 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1932_0 <=( _mesh_11_28_io_out_c_0) ^ ((fiEnable && (5582 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_28_io_in_control_0_shift_b <=( _mesh_11_28_io_out_control_0_shift) ^ ((fiEnable && (5583 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_28_io_in_control_0_dataflow_b <=( _mesh_11_28_io_out_control_0_dataflow) ^ ((fiEnable && (5584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_28_io_in_control_0_propagate_b <=( _mesh_11_28_io_out_control_0_propagate) ^ ((fiEnable && (5585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_28_io_out_valid_0) begin
			b_909_0 <=( _mesh_12_28_io_out_b_0) ^ ((fiEnable && (5586 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1933_0 <=( _mesh_12_28_io_out_c_0) ^ ((fiEnable && (5587 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_28_io_in_control_0_shift_b <=( _mesh_12_28_io_out_control_0_shift) ^ ((fiEnable && (5588 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_28_io_in_control_0_dataflow_b <=( _mesh_12_28_io_out_control_0_dataflow) ^ ((fiEnable && (5589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_28_io_in_control_0_propagate_b <=( _mesh_12_28_io_out_control_0_propagate) ^ ((fiEnable && (5590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_28_io_out_valid_0) begin
			b_910_0 <=( _mesh_13_28_io_out_b_0) ^ ((fiEnable && (5591 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1934_0 <=( _mesh_13_28_io_out_c_0) ^ ((fiEnable && (5592 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_28_io_in_control_0_shift_b <=( _mesh_13_28_io_out_control_0_shift) ^ ((fiEnable && (5593 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_28_io_in_control_0_dataflow_b <=( _mesh_13_28_io_out_control_0_dataflow) ^ ((fiEnable && (5594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_28_io_in_control_0_propagate_b <=( _mesh_13_28_io_out_control_0_propagate) ^ ((fiEnable && (5595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_28_io_out_valid_0) begin
			b_911_0 <=( _mesh_14_28_io_out_b_0) ^ ((fiEnable && (5596 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1935_0 <=( _mesh_14_28_io_out_c_0) ^ ((fiEnable && (5597 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_28_io_in_control_0_shift_b <=( _mesh_14_28_io_out_control_0_shift) ^ ((fiEnable && (5598 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_28_io_in_control_0_dataflow_b <=( _mesh_14_28_io_out_control_0_dataflow) ^ ((fiEnable && (5599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_28_io_in_control_0_propagate_b <=( _mesh_14_28_io_out_control_0_propagate) ^ ((fiEnable && (5600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_28_io_out_valid_0) begin
			b_912_0 <=( _mesh_15_28_io_out_b_0) ^ ((fiEnable && (5601 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1936_0 <=( _mesh_15_28_io_out_c_0) ^ ((fiEnable && (5602 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_28_io_in_control_0_shift_b <=( _mesh_15_28_io_out_control_0_shift) ^ ((fiEnable && (5603 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_28_io_in_control_0_dataflow_b <=( _mesh_15_28_io_out_control_0_dataflow) ^ ((fiEnable && (5604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_28_io_in_control_0_propagate_b <=( _mesh_15_28_io_out_control_0_propagate) ^ ((fiEnable && (5605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_28_io_out_valid_0) begin
			b_913_0 <=( _mesh_16_28_io_out_b_0) ^ ((fiEnable && (5606 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1937_0 <=( _mesh_16_28_io_out_c_0) ^ ((fiEnable && (5607 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_28_io_in_control_0_shift_b <=( _mesh_16_28_io_out_control_0_shift) ^ ((fiEnable && (5608 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_28_io_in_control_0_dataflow_b <=( _mesh_16_28_io_out_control_0_dataflow) ^ ((fiEnable && (5609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_28_io_in_control_0_propagate_b <=( _mesh_16_28_io_out_control_0_propagate) ^ ((fiEnable && (5610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_28_io_out_valid_0) begin
			b_914_0 <=( _mesh_17_28_io_out_b_0) ^ ((fiEnable && (5611 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1938_0 <=( _mesh_17_28_io_out_c_0) ^ ((fiEnable && (5612 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_28_io_in_control_0_shift_b <=( _mesh_17_28_io_out_control_0_shift) ^ ((fiEnable && (5613 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_28_io_in_control_0_dataflow_b <=( _mesh_17_28_io_out_control_0_dataflow) ^ ((fiEnable && (5614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_28_io_in_control_0_propagate_b <=( _mesh_17_28_io_out_control_0_propagate) ^ ((fiEnable && (5615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_28_io_out_valid_0) begin
			b_915_0 <=( _mesh_18_28_io_out_b_0) ^ ((fiEnable && (5616 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1939_0 <=( _mesh_18_28_io_out_c_0) ^ ((fiEnable && (5617 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_28_io_in_control_0_shift_b <=( _mesh_18_28_io_out_control_0_shift) ^ ((fiEnable && (5618 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_28_io_in_control_0_dataflow_b <=( _mesh_18_28_io_out_control_0_dataflow) ^ ((fiEnable && (5619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_28_io_in_control_0_propagate_b <=( _mesh_18_28_io_out_control_0_propagate) ^ ((fiEnable && (5620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_28_io_out_valid_0) begin
			b_916_0 <=( _mesh_19_28_io_out_b_0) ^ ((fiEnable && (5621 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1940_0 <=( _mesh_19_28_io_out_c_0) ^ ((fiEnable && (5622 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_28_io_in_control_0_shift_b <=( _mesh_19_28_io_out_control_0_shift) ^ ((fiEnable && (5623 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_28_io_in_control_0_dataflow_b <=( _mesh_19_28_io_out_control_0_dataflow) ^ ((fiEnable && (5624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_28_io_in_control_0_propagate_b <=( _mesh_19_28_io_out_control_0_propagate) ^ ((fiEnable && (5625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_28_io_out_valid_0) begin
			b_917_0 <=( _mesh_20_28_io_out_b_0) ^ ((fiEnable && (5626 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1941_0 <=( _mesh_20_28_io_out_c_0) ^ ((fiEnable && (5627 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_28_io_in_control_0_shift_b <=( _mesh_20_28_io_out_control_0_shift) ^ ((fiEnable && (5628 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_28_io_in_control_0_dataflow_b <=( _mesh_20_28_io_out_control_0_dataflow) ^ ((fiEnable && (5629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_28_io_in_control_0_propagate_b <=( _mesh_20_28_io_out_control_0_propagate) ^ ((fiEnable && (5630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_28_io_out_valid_0) begin
			b_918_0 <=( _mesh_21_28_io_out_b_0) ^ ((fiEnable && (5631 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1942_0 <=( _mesh_21_28_io_out_c_0) ^ ((fiEnable && (5632 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_28_io_in_control_0_shift_b <=( _mesh_21_28_io_out_control_0_shift) ^ ((fiEnable && (5633 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_28_io_in_control_0_dataflow_b <=( _mesh_21_28_io_out_control_0_dataflow) ^ ((fiEnable && (5634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_28_io_in_control_0_propagate_b <=( _mesh_21_28_io_out_control_0_propagate) ^ ((fiEnable && (5635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_28_io_out_valid_0) begin
			b_919_0 <=( _mesh_22_28_io_out_b_0) ^ ((fiEnable && (5636 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1943_0 <=( _mesh_22_28_io_out_c_0) ^ ((fiEnable && (5637 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_28_io_in_control_0_shift_b <=( _mesh_22_28_io_out_control_0_shift) ^ ((fiEnable && (5638 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_28_io_in_control_0_dataflow_b <=( _mesh_22_28_io_out_control_0_dataflow) ^ ((fiEnable && (5639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_28_io_in_control_0_propagate_b <=( _mesh_22_28_io_out_control_0_propagate) ^ ((fiEnable && (5640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_28_io_out_valid_0) begin
			b_920_0 <=( _mesh_23_28_io_out_b_0) ^ ((fiEnable && (5641 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1944_0 <=( _mesh_23_28_io_out_c_0) ^ ((fiEnable && (5642 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_28_io_in_control_0_shift_b <=( _mesh_23_28_io_out_control_0_shift) ^ ((fiEnable && (5643 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_28_io_in_control_0_dataflow_b <=( _mesh_23_28_io_out_control_0_dataflow) ^ ((fiEnable && (5644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_28_io_in_control_0_propagate_b <=( _mesh_23_28_io_out_control_0_propagate) ^ ((fiEnable && (5645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_28_io_out_valid_0) begin
			b_921_0 <=( _mesh_24_28_io_out_b_0) ^ ((fiEnable && (5646 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1945_0 <=( _mesh_24_28_io_out_c_0) ^ ((fiEnable && (5647 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_28_io_in_control_0_shift_b <=( _mesh_24_28_io_out_control_0_shift) ^ ((fiEnable && (5648 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_28_io_in_control_0_dataflow_b <=( _mesh_24_28_io_out_control_0_dataflow) ^ ((fiEnable && (5649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_28_io_in_control_0_propagate_b <=( _mesh_24_28_io_out_control_0_propagate) ^ ((fiEnable && (5650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_28_io_out_valid_0) begin
			b_922_0 <=( _mesh_25_28_io_out_b_0) ^ ((fiEnable && (5651 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1946_0 <=( _mesh_25_28_io_out_c_0) ^ ((fiEnable && (5652 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_28_io_in_control_0_shift_b <=( _mesh_25_28_io_out_control_0_shift) ^ ((fiEnable && (5653 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_28_io_in_control_0_dataflow_b <=( _mesh_25_28_io_out_control_0_dataflow) ^ ((fiEnable && (5654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_28_io_in_control_0_propagate_b <=( _mesh_25_28_io_out_control_0_propagate) ^ ((fiEnable && (5655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_28_io_out_valid_0) begin
			b_923_0 <=( _mesh_26_28_io_out_b_0) ^ ((fiEnable && (5656 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1947_0 <=( _mesh_26_28_io_out_c_0) ^ ((fiEnable && (5657 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_28_io_in_control_0_shift_b <=( _mesh_26_28_io_out_control_0_shift) ^ ((fiEnable && (5658 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_28_io_in_control_0_dataflow_b <=( _mesh_26_28_io_out_control_0_dataflow) ^ ((fiEnable && (5659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_28_io_in_control_0_propagate_b <=( _mesh_26_28_io_out_control_0_propagate) ^ ((fiEnable && (5660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_28_io_out_valid_0) begin
			b_924_0 <=( _mesh_27_28_io_out_b_0) ^ ((fiEnable && (5661 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1948_0 <=( _mesh_27_28_io_out_c_0) ^ ((fiEnable && (5662 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_28_io_in_control_0_shift_b <=( _mesh_27_28_io_out_control_0_shift) ^ ((fiEnable && (5663 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_28_io_in_control_0_dataflow_b <=( _mesh_27_28_io_out_control_0_dataflow) ^ ((fiEnable && (5664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_28_io_in_control_0_propagate_b <=( _mesh_27_28_io_out_control_0_propagate) ^ ((fiEnable && (5665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_28_io_out_valid_0) begin
			b_925_0 <=( _mesh_28_28_io_out_b_0) ^ ((fiEnable && (5666 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1949_0 <=( _mesh_28_28_io_out_c_0) ^ ((fiEnable && (5667 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_28_io_in_control_0_shift_b <=( _mesh_28_28_io_out_control_0_shift) ^ ((fiEnable && (5668 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_28_io_in_control_0_dataflow_b <=( _mesh_28_28_io_out_control_0_dataflow) ^ ((fiEnable && (5669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_28_io_in_control_0_propagate_b <=( _mesh_28_28_io_out_control_0_propagate) ^ ((fiEnable && (5670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_28_io_out_valid_0) begin
			b_926_0 <=( _mesh_29_28_io_out_b_0) ^ ((fiEnable && (5671 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1950_0 <=( _mesh_29_28_io_out_c_0) ^ ((fiEnable && (5672 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_28_io_in_control_0_shift_b <=( _mesh_29_28_io_out_control_0_shift) ^ ((fiEnable && (5673 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_28_io_in_control_0_dataflow_b <=( _mesh_29_28_io_out_control_0_dataflow) ^ ((fiEnable && (5674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_28_io_in_control_0_propagate_b <=( _mesh_29_28_io_out_control_0_propagate) ^ ((fiEnable && (5675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_28_io_out_valid_0) begin
			b_927_0 <=( _mesh_30_28_io_out_b_0) ^ ((fiEnable && (5676 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1951_0 <=( _mesh_30_28_io_out_c_0) ^ ((fiEnable && (5677 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_28_io_in_control_0_shift_b <=( _mesh_30_28_io_out_control_0_shift) ^ ((fiEnable && (5678 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_28_io_in_control_0_dataflow_b <=( _mesh_30_28_io_out_control_0_dataflow) ^ ((fiEnable && (5679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_28_io_in_control_0_propagate_b <=( _mesh_30_28_io_out_control_0_propagate) ^ ((fiEnable && (5680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_29_0) begin
			b_928_0 <=( io_in_b_29_0) ^ ((fiEnable && (5681 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1952_0 <=( io_in_d_29_0) ^ ((fiEnable && (5682 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_29_io_in_control_0_shift_b <=( io_in_control_29_0_shift) ^ ((fiEnable && (5683 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_29_io_in_control_0_dataflow_b <=( io_in_control_29_0_dataflow) ^ ((fiEnable && (5684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_29_io_in_control_0_propagate_b <=( io_in_control_29_0_propagate) ^ ((fiEnable && (5685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_29_io_out_valid_0) begin
			b_929_0 <=( _mesh_0_29_io_out_b_0) ^ ((fiEnable && (5686 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1953_0 <=( _mesh_0_29_io_out_c_0) ^ ((fiEnable && (5687 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_29_io_in_control_0_shift_b <=( _mesh_0_29_io_out_control_0_shift) ^ ((fiEnable && (5688 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_29_io_in_control_0_dataflow_b <=( _mesh_0_29_io_out_control_0_dataflow) ^ ((fiEnable && (5689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_29_io_in_control_0_propagate_b <=( _mesh_0_29_io_out_control_0_propagate) ^ ((fiEnable && (5690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_29_io_out_valid_0) begin
			b_930_0 <=( _mesh_1_29_io_out_b_0) ^ ((fiEnable && (5691 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1954_0 <=( _mesh_1_29_io_out_c_0) ^ ((fiEnable && (5692 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_29_io_in_control_0_shift_b <=( _mesh_1_29_io_out_control_0_shift) ^ ((fiEnable && (5693 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_29_io_in_control_0_dataflow_b <=( _mesh_1_29_io_out_control_0_dataflow) ^ ((fiEnable && (5694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_29_io_in_control_0_propagate_b <=( _mesh_1_29_io_out_control_0_propagate) ^ ((fiEnable && (5695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_29_io_out_valid_0) begin
			b_931_0 <=( _mesh_2_29_io_out_b_0) ^ ((fiEnable && (5696 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1955_0 <=( _mesh_2_29_io_out_c_0) ^ ((fiEnable && (5697 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_29_io_in_control_0_shift_b <=( _mesh_2_29_io_out_control_0_shift) ^ ((fiEnable && (5698 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_29_io_in_control_0_dataflow_b <=( _mesh_2_29_io_out_control_0_dataflow) ^ ((fiEnable && (5699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_29_io_in_control_0_propagate_b <=( _mesh_2_29_io_out_control_0_propagate) ^ ((fiEnable && (5700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_29_io_out_valid_0) begin
			b_932_0 <=( _mesh_3_29_io_out_b_0) ^ ((fiEnable && (5701 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1956_0 <=( _mesh_3_29_io_out_c_0) ^ ((fiEnable && (5702 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_29_io_in_control_0_shift_b <=( _mesh_3_29_io_out_control_0_shift) ^ ((fiEnable && (5703 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_29_io_in_control_0_dataflow_b <=( _mesh_3_29_io_out_control_0_dataflow) ^ ((fiEnable && (5704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_29_io_in_control_0_propagate_b <=( _mesh_3_29_io_out_control_0_propagate) ^ ((fiEnable && (5705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_29_io_out_valid_0) begin
			b_933_0 <=( _mesh_4_29_io_out_b_0) ^ ((fiEnable && (5706 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1957_0 <=( _mesh_4_29_io_out_c_0) ^ ((fiEnable && (5707 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_29_io_in_control_0_shift_b <=( _mesh_4_29_io_out_control_0_shift) ^ ((fiEnable && (5708 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_29_io_in_control_0_dataflow_b <=( _mesh_4_29_io_out_control_0_dataflow) ^ ((fiEnable && (5709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_29_io_in_control_0_propagate_b <=( _mesh_4_29_io_out_control_0_propagate) ^ ((fiEnable && (5710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_29_io_out_valid_0) begin
			b_934_0 <=( _mesh_5_29_io_out_b_0) ^ ((fiEnable && (5711 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1958_0 <=( _mesh_5_29_io_out_c_0) ^ ((fiEnable && (5712 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_29_io_in_control_0_shift_b <=( _mesh_5_29_io_out_control_0_shift) ^ ((fiEnable && (5713 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_29_io_in_control_0_dataflow_b <=( _mesh_5_29_io_out_control_0_dataflow) ^ ((fiEnable && (5714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_29_io_in_control_0_propagate_b <=( _mesh_5_29_io_out_control_0_propagate) ^ ((fiEnable && (5715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_29_io_out_valid_0) begin
			b_935_0 <=( _mesh_6_29_io_out_b_0) ^ ((fiEnable && (5716 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1959_0 <=( _mesh_6_29_io_out_c_0) ^ ((fiEnable && (5717 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_29_io_in_control_0_shift_b <=( _mesh_6_29_io_out_control_0_shift) ^ ((fiEnable && (5718 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_29_io_in_control_0_dataflow_b <=( _mesh_6_29_io_out_control_0_dataflow) ^ ((fiEnable && (5719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_29_io_in_control_0_propagate_b <=( _mesh_6_29_io_out_control_0_propagate) ^ ((fiEnable && (5720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_29_io_out_valid_0) begin
			b_936_0 <=( _mesh_7_29_io_out_b_0) ^ ((fiEnable && (5721 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1960_0 <=( _mesh_7_29_io_out_c_0) ^ ((fiEnable && (5722 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_29_io_in_control_0_shift_b <=( _mesh_7_29_io_out_control_0_shift) ^ ((fiEnable && (5723 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_29_io_in_control_0_dataflow_b <=( _mesh_7_29_io_out_control_0_dataflow) ^ ((fiEnable && (5724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_29_io_in_control_0_propagate_b <=( _mesh_7_29_io_out_control_0_propagate) ^ ((fiEnable && (5725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_29_io_out_valid_0) begin
			b_937_0 <=( _mesh_8_29_io_out_b_0) ^ ((fiEnable && (5726 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1961_0 <=( _mesh_8_29_io_out_c_0) ^ ((fiEnable && (5727 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_29_io_in_control_0_shift_b <=( _mesh_8_29_io_out_control_0_shift) ^ ((fiEnable && (5728 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_29_io_in_control_0_dataflow_b <=( _mesh_8_29_io_out_control_0_dataflow) ^ ((fiEnable && (5729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_29_io_in_control_0_propagate_b <=( _mesh_8_29_io_out_control_0_propagate) ^ ((fiEnable && (5730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_29_io_out_valid_0) begin
			b_938_0 <=( _mesh_9_29_io_out_b_0) ^ ((fiEnable && (5731 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1962_0 <=( _mesh_9_29_io_out_c_0) ^ ((fiEnable && (5732 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_29_io_in_control_0_shift_b <=( _mesh_9_29_io_out_control_0_shift) ^ ((fiEnable && (5733 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_29_io_in_control_0_dataflow_b <=( _mesh_9_29_io_out_control_0_dataflow) ^ ((fiEnable && (5734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_29_io_in_control_0_propagate_b <=( _mesh_9_29_io_out_control_0_propagate) ^ ((fiEnable && (5735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_29_io_out_valid_0) begin
			b_939_0 <=( _mesh_10_29_io_out_b_0) ^ ((fiEnable && (5736 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1963_0 <=( _mesh_10_29_io_out_c_0) ^ ((fiEnable && (5737 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_29_io_in_control_0_shift_b <=( _mesh_10_29_io_out_control_0_shift) ^ ((fiEnable && (5738 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_29_io_in_control_0_dataflow_b <=( _mesh_10_29_io_out_control_0_dataflow) ^ ((fiEnable && (5739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_29_io_in_control_0_propagate_b <=( _mesh_10_29_io_out_control_0_propagate) ^ ((fiEnable && (5740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_29_io_out_valid_0) begin
			b_940_0 <=( _mesh_11_29_io_out_b_0) ^ ((fiEnable && (5741 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1964_0 <=( _mesh_11_29_io_out_c_0) ^ ((fiEnable && (5742 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_29_io_in_control_0_shift_b <=( _mesh_11_29_io_out_control_0_shift) ^ ((fiEnable && (5743 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_29_io_in_control_0_dataflow_b <=( _mesh_11_29_io_out_control_0_dataflow) ^ ((fiEnable && (5744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_29_io_in_control_0_propagate_b <=( _mesh_11_29_io_out_control_0_propagate) ^ ((fiEnable && (5745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_29_io_out_valid_0) begin
			b_941_0 <=( _mesh_12_29_io_out_b_0) ^ ((fiEnable && (5746 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1965_0 <=( _mesh_12_29_io_out_c_0) ^ ((fiEnable && (5747 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_29_io_in_control_0_shift_b <=( _mesh_12_29_io_out_control_0_shift) ^ ((fiEnable && (5748 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_29_io_in_control_0_dataflow_b <=( _mesh_12_29_io_out_control_0_dataflow) ^ ((fiEnable && (5749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_29_io_in_control_0_propagate_b <=( _mesh_12_29_io_out_control_0_propagate) ^ ((fiEnable && (5750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_29_io_out_valid_0) begin
			b_942_0 <=( _mesh_13_29_io_out_b_0) ^ ((fiEnable && (5751 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1966_0 <=( _mesh_13_29_io_out_c_0) ^ ((fiEnable && (5752 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_29_io_in_control_0_shift_b <=( _mesh_13_29_io_out_control_0_shift) ^ ((fiEnable && (5753 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_29_io_in_control_0_dataflow_b <=( _mesh_13_29_io_out_control_0_dataflow) ^ ((fiEnable && (5754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_29_io_in_control_0_propagate_b <=( _mesh_13_29_io_out_control_0_propagate) ^ ((fiEnable && (5755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_29_io_out_valid_0) begin
			b_943_0 <=( _mesh_14_29_io_out_b_0) ^ ((fiEnable && (5756 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1967_0 <=( _mesh_14_29_io_out_c_0) ^ ((fiEnable && (5757 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_29_io_in_control_0_shift_b <=( _mesh_14_29_io_out_control_0_shift) ^ ((fiEnable && (5758 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_29_io_in_control_0_dataflow_b <=( _mesh_14_29_io_out_control_0_dataflow) ^ ((fiEnable && (5759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_29_io_in_control_0_propagate_b <=( _mesh_14_29_io_out_control_0_propagate) ^ ((fiEnable && (5760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_29_io_out_valid_0) begin
			b_944_0 <=( _mesh_15_29_io_out_b_0) ^ ((fiEnable && (5761 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1968_0 <=( _mesh_15_29_io_out_c_0) ^ ((fiEnable && (5762 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_29_io_in_control_0_shift_b <=( _mesh_15_29_io_out_control_0_shift) ^ ((fiEnable && (5763 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_29_io_in_control_0_dataflow_b <=( _mesh_15_29_io_out_control_0_dataflow) ^ ((fiEnable && (5764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_29_io_in_control_0_propagate_b <=( _mesh_15_29_io_out_control_0_propagate) ^ ((fiEnable && (5765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_29_io_out_valid_0) begin
			b_945_0 <=( _mesh_16_29_io_out_b_0) ^ ((fiEnable && (5766 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1969_0 <=( _mesh_16_29_io_out_c_0) ^ ((fiEnable && (5767 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_29_io_in_control_0_shift_b <=( _mesh_16_29_io_out_control_0_shift) ^ ((fiEnable && (5768 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_29_io_in_control_0_dataflow_b <=( _mesh_16_29_io_out_control_0_dataflow) ^ ((fiEnable && (5769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_29_io_in_control_0_propagate_b <=( _mesh_16_29_io_out_control_0_propagate) ^ ((fiEnable && (5770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_29_io_out_valid_0) begin
			b_946_0 <=( _mesh_17_29_io_out_b_0) ^ ((fiEnable && (5771 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1970_0 <=( _mesh_17_29_io_out_c_0) ^ ((fiEnable && (5772 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_29_io_in_control_0_shift_b <=( _mesh_17_29_io_out_control_0_shift) ^ ((fiEnable && (5773 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_29_io_in_control_0_dataflow_b <=( _mesh_17_29_io_out_control_0_dataflow) ^ ((fiEnable && (5774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_29_io_in_control_0_propagate_b <=( _mesh_17_29_io_out_control_0_propagate) ^ ((fiEnable && (5775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_29_io_out_valid_0) begin
			b_947_0 <=( _mesh_18_29_io_out_b_0) ^ ((fiEnable && (5776 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1971_0 <=( _mesh_18_29_io_out_c_0) ^ ((fiEnable && (5777 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_29_io_in_control_0_shift_b <=( _mesh_18_29_io_out_control_0_shift) ^ ((fiEnable && (5778 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_29_io_in_control_0_dataflow_b <=( _mesh_18_29_io_out_control_0_dataflow) ^ ((fiEnable && (5779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_29_io_in_control_0_propagate_b <=( _mesh_18_29_io_out_control_0_propagate) ^ ((fiEnable && (5780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_29_io_out_valid_0) begin
			b_948_0 <=( _mesh_19_29_io_out_b_0) ^ ((fiEnable && (5781 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1972_0 <=( _mesh_19_29_io_out_c_0) ^ ((fiEnable && (5782 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_29_io_in_control_0_shift_b <=( _mesh_19_29_io_out_control_0_shift) ^ ((fiEnable && (5783 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_29_io_in_control_0_dataflow_b <=( _mesh_19_29_io_out_control_0_dataflow) ^ ((fiEnable && (5784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_29_io_in_control_0_propagate_b <=( _mesh_19_29_io_out_control_0_propagate) ^ ((fiEnable && (5785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_29_io_out_valid_0) begin
			b_949_0 <=( _mesh_20_29_io_out_b_0) ^ ((fiEnable && (5786 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1973_0 <=( _mesh_20_29_io_out_c_0) ^ ((fiEnable && (5787 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_29_io_in_control_0_shift_b <=( _mesh_20_29_io_out_control_0_shift) ^ ((fiEnable && (5788 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_29_io_in_control_0_dataflow_b <=( _mesh_20_29_io_out_control_0_dataflow) ^ ((fiEnable && (5789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_29_io_in_control_0_propagate_b <=( _mesh_20_29_io_out_control_0_propagate) ^ ((fiEnable && (5790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_29_io_out_valid_0) begin
			b_950_0 <=( _mesh_21_29_io_out_b_0) ^ ((fiEnable && (5791 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1974_0 <=( _mesh_21_29_io_out_c_0) ^ ((fiEnable && (5792 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_29_io_in_control_0_shift_b <=( _mesh_21_29_io_out_control_0_shift) ^ ((fiEnable && (5793 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_29_io_in_control_0_dataflow_b <=( _mesh_21_29_io_out_control_0_dataflow) ^ ((fiEnable && (5794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_29_io_in_control_0_propagate_b <=( _mesh_21_29_io_out_control_0_propagate) ^ ((fiEnable && (5795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_29_io_out_valid_0) begin
			b_951_0 <=( _mesh_22_29_io_out_b_0) ^ ((fiEnable && (5796 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1975_0 <=( _mesh_22_29_io_out_c_0) ^ ((fiEnable && (5797 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_29_io_in_control_0_shift_b <=( _mesh_22_29_io_out_control_0_shift) ^ ((fiEnable && (5798 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_29_io_in_control_0_dataflow_b <=( _mesh_22_29_io_out_control_0_dataflow) ^ ((fiEnable && (5799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_29_io_in_control_0_propagate_b <=( _mesh_22_29_io_out_control_0_propagate) ^ ((fiEnable && (5800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_29_io_out_valid_0) begin
			b_952_0 <=( _mesh_23_29_io_out_b_0) ^ ((fiEnable && (5801 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1976_0 <=( _mesh_23_29_io_out_c_0) ^ ((fiEnable && (5802 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_29_io_in_control_0_shift_b <=( _mesh_23_29_io_out_control_0_shift) ^ ((fiEnable && (5803 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_29_io_in_control_0_dataflow_b <=( _mesh_23_29_io_out_control_0_dataflow) ^ ((fiEnable && (5804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_29_io_in_control_0_propagate_b <=( _mesh_23_29_io_out_control_0_propagate) ^ ((fiEnable && (5805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_29_io_out_valid_0) begin
			b_953_0 <=( _mesh_24_29_io_out_b_0) ^ ((fiEnable && (5806 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1977_0 <=( _mesh_24_29_io_out_c_0) ^ ((fiEnable && (5807 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_29_io_in_control_0_shift_b <=( _mesh_24_29_io_out_control_0_shift) ^ ((fiEnable && (5808 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_29_io_in_control_0_dataflow_b <=( _mesh_24_29_io_out_control_0_dataflow) ^ ((fiEnable && (5809 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_29_io_in_control_0_propagate_b <=( _mesh_24_29_io_out_control_0_propagate) ^ ((fiEnable && (5810 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_29_io_out_valid_0) begin
			b_954_0 <=( _mesh_25_29_io_out_b_0) ^ ((fiEnable && (5811 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1978_0 <=( _mesh_25_29_io_out_c_0) ^ ((fiEnable && (5812 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_29_io_in_control_0_shift_b <=( _mesh_25_29_io_out_control_0_shift) ^ ((fiEnable && (5813 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_29_io_in_control_0_dataflow_b <=( _mesh_25_29_io_out_control_0_dataflow) ^ ((fiEnable && (5814 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_29_io_in_control_0_propagate_b <=( _mesh_25_29_io_out_control_0_propagate) ^ ((fiEnable && (5815 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_29_io_out_valid_0) begin
			b_955_0 <=( _mesh_26_29_io_out_b_0) ^ ((fiEnable && (5816 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1979_0 <=( _mesh_26_29_io_out_c_0) ^ ((fiEnable && (5817 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_29_io_in_control_0_shift_b <=( _mesh_26_29_io_out_control_0_shift) ^ ((fiEnable && (5818 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_29_io_in_control_0_dataflow_b <=( _mesh_26_29_io_out_control_0_dataflow) ^ ((fiEnable && (5819 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_29_io_in_control_0_propagate_b <=( _mesh_26_29_io_out_control_0_propagate) ^ ((fiEnable && (5820 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_29_io_out_valid_0) begin
			b_956_0 <=( _mesh_27_29_io_out_b_0) ^ ((fiEnable && (5821 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1980_0 <=( _mesh_27_29_io_out_c_0) ^ ((fiEnable && (5822 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_29_io_in_control_0_shift_b <=( _mesh_27_29_io_out_control_0_shift) ^ ((fiEnable && (5823 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_29_io_in_control_0_dataflow_b <=( _mesh_27_29_io_out_control_0_dataflow) ^ ((fiEnable && (5824 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_29_io_in_control_0_propagate_b <=( _mesh_27_29_io_out_control_0_propagate) ^ ((fiEnable && (5825 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_29_io_out_valid_0) begin
			b_957_0 <=( _mesh_28_29_io_out_b_0) ^ ((fiEnable && (5826 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1981_0 <=( _mesh_28_29_io_out_c_0) ^ ((fiEnable && (5827 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_29_io_in_control_0_shift_b <=( _mesh_28_29_io_out_control_0_shift) ^ ((fiEnable && (5828 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_29_io_in_control_0_dataflow_b <=( _mesh_28_29_io_out_control_0_dataflow) ^ ((fiEnable && (5829 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_29_io_in_control_0_propagate_b <=( _mesh_28_29_io_out_control_0_propagate) ^ ((fiEnable && (5830 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_29_io_out_valid_0) begin
			b_958_0 <=( _mesh_29_29_io_out_b_0) ^ ((fiEnable && (5831 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1982_0 <=( _mesh_29_29_io_out_c_0) ^ ((fiEnable && (5832 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_29_io_in_control_0_shift_b <=( _mesh_29_29_io_out_control_0_shift) ^ ((fiEnable && (5833 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_29_io_in_control_0_dataflow_b <=( _mesh_29_29_io_out_control_0_dataflow) ^ ((fiEnable && (5834 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_29_io_in_control_0_propagate_b <=( _mesh_29_29_io_out_control_0_propagate) ^ ((fiEnable && (5835 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_29_io_out_valid_0) begin
			b_959_0 <=( _mesh_30_29_io_out_b_0) ^ ((fiEnable && (5836 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1983_0 <=( _mesh_30_29_io_out_c_0) ^ ((fiEnable && (5837 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_29_io_in_control_0_shift_b <=( _mesh_30_29_io_out_control_0_shift) ^ ((fiEnable && (5838 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_29_io_in_control_0_dataflow_b <=( _mesh_30_29_io_out_control_0_dataflow) ^ ((fiEnable && (5839 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_29_io_in_control_0_propagate_b <=( _mesh_30_29_io_out_control_0_propagate) ^ ((fiEnable && (5840 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_30_0) begin
			b_960_0 <=( io_in_b_30_0) ^ ((fiEnable && (5841 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1984_0 <=( io_in_d_30_0) ^ ((fiEnable && (5842 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_30_io_in_control_0_shift_b <=( io_in_control_30_0_shift) ^ ((fiEnable && (5843 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_30_io_in_control_0_dataflow_b <=( io_in_control_30_0_dataflow) ^ ((fiEnable && (5844 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_30_io_in_control_0_propagate_b <=( io_in_control_30_0_propagate) ^ ((fiEnable && (5845 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_30_io_out_valid_0) begin
			b_961_0 <=( _mesh_0_30_io_out_b_0) ^ ((fiEnable && (5846 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1985_0 <=( _mesh_0_30_io_out_c_0) ^ ((fiEnable && (5847 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_30_io_in_control_0_shift_b <=( _mesh_0_30_io_out_control_0_shift) ^ ((fiEnable && (5848 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_30_io_in_control_0_dataflow_b <=( _mesh_0_30_io_out_control_0_dataflow) ^ ((fiEnable && (5849 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_30_io_in_control_0_propagate_b <=( _mesh_0_30_io_out_control_0_propagate) ^ ((fiEnable && (5850 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_30_io_out_valid_0) begin
			b_962_0 <=( _mesh_1_30_io_out_b_0) ^ ((fiEnable && (5851 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1986_0 <=( _mesh_1_30_io_out_c_0) ^ ((fiEnable && (5852 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_30_io_in_control_0_shift_b <=( _mesh_1_30_io_out_control_0_shift) ^ ((fiEnable && (5853 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_30_io_in_control_0_dataflow_b <=( _mesh_1_30_io_out_control_0_dataflow) ^ ((fiEnable && (5854 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_30_io_in_control_0_propagate_b <=( _mesh_1_30_io_out_control_0_propagate) ^ ((fiEnable && (5855 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_30_io_out_valid_0) begin
			b_963_0 <=( _mesh_2_30_io_out_b_0) ^ ((fiEnable && (5856 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1987_0 <=( _mesh_2_30_io_out_c_0) ^ ((fiEnable && (5857 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_30_io_in_control_0_shift_b <=( _mesh_2_30_io_out_control_0_shift) ^ ((fiEnable && (5858 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_30_io_in_control_0_dataflow_b <=( _mesh_2_30_io_out_control_0_dataflow) ^ ((fiEnable && (5859 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_30_io_in_control_0_propagate_b <=( _mesh_2_30_io_out_control_0_propagate) ^ ((fiEnable && (5860 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_30_io_out_valid_0) begin
			b_964_0 <=( _mesh_3_30_io_out_b_0) ^ ((fiEnable && (5861 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1988_0 <=( _mesh_3_30_io_out_c_0) ^ ((fiEnable && (5862 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_30_io_in_control_0_shift_b <=( _mesh_3_30_io_out_control_0_shift) ^ ((fiEnable && (5863 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_30_io_in_control_0_dataflow_b <=( _mesh_3_30_io_out_control_0_dataflow) ^ ((fiEnable && (5864 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_30_io_in_control_0_propagate_b <=( _mesh_3_30_io_out_control_0_propagate) ^ ((fiEnable && (5865 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_30_io_out_valid_0) begin
			b_965_0 <=( _mesh_4_30_io_out_b_0) ^ ((fiEnable && (5866 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1989_0 <=( _mesh_4_30_io_out_c_0) ^ ((fiEnable && (5867 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_30_io_in_control_0_shift_b <=( _mesh_4_30_io_out_control_0_shift) ^ ((fiEnable && (5868 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_30_io_in_control_0_dataflow_b <=( _mesh_4_30_io_out_control_0_dataflow) ^ ((fiEnable && (5869 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_30_io_in_control_0_propagate_b <=( _mesh_4_30_io_out_control_0_propagate) ^ ((fiEnable && (5870 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_30_io_out_valid_0) begin
			b_966_0 <=( _mesh_5_30_io_out_b_0) ^ ((fiEnable && (5871 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1990_0 <=( _mesh_5_30_io_out_c_0) ^ ((fiEnable && (5872 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_30_io_in_control_0_shift_b <=( _mesh_5_30_io_out_control_0_shift) ^ ((fiEnable && (5873 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_30_io_in_control_0_dataflow_b <=( _mesh_5_30_io_out_control_0_dataflow) ^ ((fiEnable && (5874 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_30_io_in_control_0_propagate_b <=( _mesh_5_30_io_out_control_0_propagate) ^ ((fiEnable && (5875 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_30_io_out_valid_0) begin
			b_967_0 <=( _mesh_6_30_io_out_b_0) ^ ((fiEnable && (5876 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1991_0 <=( _mesh_6_30_io_out_c_0) ^ ((fiEnable && (5877 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_30_io_in_control_0_shift_b <=( _mesh_6_30_io_out_control_0_shift) ^ ((fiEnable && (5878 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_30_io_in_control_0_dataflow_b <=( _mesh_6_30_io_out_control_0_dataflow) ^ ((fiEnable && (5879 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_30_io_in_control_0_propagate_b <=( _mesh_6_30_io_out_control_0_propagate) ^ ((fiEnable && (5880 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_30_io_out_valid_0) begin
			b_968_0 <=( _mesh_7_30_io_out_b_0) ^ ((fiEnable && (5881 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1992_0 <=( _mesh_7_30_io_out_c_0) ^ ((fiEnable && (5882 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_30_io_in_control_0_shift_b <=( _mesh_7_30_io_out_control_0_shift) ^ ((fiEnable && (5883 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_30_io_in_control_0_dataflow_b <=( _mesh_7_30_io_out_control_0_dataflow) ^ ((fiEnable && (5884 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_30_io_in_control_0_propagate_b <=( _mesh_7_30_io_out_control_0_propagate) ^ ((fiEnable && (5885 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_30_io_out_valid_0) begin
			b_969_0 <=( _mesh_8_30_io_out_b_0) ^ ((fiEnable && (5886 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1993_0 <=( _mesh_8_30_io_out_c_0) ^ ((fiEnable && (5887 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_30_io_in_control_0_shift_b <=( _mesh_8_30_io_out_control_0_shift) ^ ((fiEnable && (5888 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_30_io_in_control_0_dataflow_b <=( _mesh_8_30_io_out_control_0_dataflow) ^ ((fiEnable && (5889 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_30_io_in_control_0_propagate_b <=( _mesh_8_30_io_out_control_0_propagate) ^ ((fiEnable && (5890 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_30_io_out_valid_0) begin
			b_970_0 <=( _mesh_9_30_io_out_b_0) ^ ((fiEnable && (5891 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1994_0 <=( _mesh_9_30_io_out_c_0) ^ ((fiEnable && (5892 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_30_io_in_control_0_shift_b <=( _mesh_9_30_io_out_control_0_shift) ^ ((fiEnable && (5893 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_30_io_in_control_0_dataflow_b <=( _mesh_9_30_io_out_control_0_dataflow) ^ ((fiEnable && (5894 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_30_io_in_control_0_propagate_b <=( _mesh_9_30_io_out_control_0_propagate) ^ ((fiEnable && (5895 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_30_io_out_valid_0) begin
			b_971_0 <=( _mesh_10_30_io_out_b_0) ^ ((fiEnable && (5896 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1995_0 <=( _mesh_10_30_io_out_c_0) ^ ((fiEnable && (5897 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_30_io_in_control_0_shift_b <=( _mesh_10_30_io_out_control_0_shift) ^ ((fiEnable && (5898 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_30_io_in_control_0_dataflow_b <=( _mesh_10_30_io_out_control_0_dataflow) ^ ((fiEnable && (5899 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_30_io_in_control_0_propagate_b <=( _mesh_10_30_io_out_control_0_propagate) ^ ((fiEnable && (5900 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_30_io_out_valid_0) begin
			b_972_0 <=( _mesh_11_30_io_out_b_0) ^ ((fiEnable && (5901 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1996_0 <=( _mesh_11_30_io_out_c_0) ^ ((fiEnable && (5902 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_30_io_in_control_0_shift_b <=( _mesh_11_30_io_out_control_0_shift) ^ ((fiEnable && (5903 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_30_io_in_control_0_dataflow_b <=( _mesh_11_30_io_out_control_0_dataflow) ^ ((fiEnable && (5904 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_30_io_in_control_0_propagate_b <=( _mesh_11_30_io_out_control_0_propagate) ^ ((fiEnable && (5905 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_30_io_out_valid_0) begin
			b_973_0 <=( _mesh_12_30_io_out_b_0) ^ ((fiEnable && (5906 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1997_0 <=( _mesh_12_30_io_out_c_0) ^ ((fiEnable && (5907 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_30_io_in_control_0_shift_b <=( _mesh_12_30_io_out_control_0_shift) ^ ((fiEnable && (5908 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_30_io_in_control_0_dataflow_b <=( _mesh_12_30_io_out_control_0_dataflow) ^ ((fiEnable && (5909 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_30_io_in_control_0_propagate_b <=( _mesh_12_30_io_out_control_0_propagate) ^ ((fiEnable && (5910 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_30_io_out_valid_0) begin
			b_974_0 <=( _mesh_13_30_io_out_b_0) ^ ((fiEnable && (5911 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1998_0 <=( _mesh_13_30_io_out_c_0) ^ ((fiEnable && (5912 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_30_io_in_control_0_shift_b <=( _mesh_13_30_io_out_control_0_shift) ^ ((fiEnable && (5913 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_30_io_in_control_0_dataflow_b <=( _mesh_13_30_io_out_control_0_dataflow) ^ ((fiEnable && (5914 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_30_io_in_control_0_propagate_b <=( _mesh_13_30_io_out_control_0_propagate) ^ ((fiEnable && (5915 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_30_io_out_valid_0) begin
			b_975_0 <=( _mesh_14_30_io_out_b_0) ^ ((fiEnable && (5916 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_1999_0 <=( _mesh_14_30_io_out_c_0) ^ ((fiEnable && (5917 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_30_io_in_control_0_shift_b <=( _mesh_14_30_io_out_control_0_shift) ^ ((fiEnable && (5918 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_30_io_in_control_0_dataflow_b <=( _mesh_14_30_io_out_control_0_dataflow) ^ ((fiEnable && (5919 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_30_io_in_control_0_propagate_b <=( _mesh_14_30_io_out_control_0_propagate) ^ ((fiEnable && (5920 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_30_io_out_valid_0) begin
			b_976_0 <=( _mesh_15_30_io_out_b_0) ^ ((fiEnable && (5921 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2000_0 <=( _mesh_15_30_io_out_c_0) ^ ((fiEnable && (5922 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_30_io_in_control_0_shift_b <=( _mesh_15_30_io_out_control_0_shift) ^ ((fiEnable && (5923 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_30_io_in_control_0_dataflow_b <=( _mesh_15_30_io_out_control_0_dataflow) ^ ((fiEnable && (5924 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_30_io_in_control_0_propagate_b <=( _mesh_15_30_io_out_control_0_propagate) ^ ((fiEnable && (5925 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_30_io_out_valid_0) begin
			b_977_0 <=( _mesh_16_30_io_out_b_0) ^ ((fiEnable && (5926 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2001_0 <=( _mesh_16_30_io_out_c_0) ^ ((fiEnable && (5927 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_30_io_in_control_0_shift_b <=( _mesh_16_30_io_out_control_0_shift) ^ ((fiEnable && (5928 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_30_io_in_control_0_dataflow_b <=( _mesh_16_30_io_out_control_0_dataflow) ^ ((fiEnable && (5929 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_30_io_in_control_0_propagate_b <=( _mesh_16_30_io_out_control_0_propagate) ^ ((fiEnable && (5930 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_30_io_out_valid_0) begin
			b_978_0 <=( _mesh_17_30_io_out_b_0) ^ ((fiEnable && (5931 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2002_0 <=( _mesh_17_30_io_out_c_0) ^ ((fiEnable && (5932 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_30_io_in_control_0_shift_b <=( _mesh_17_30_io_out_control_0_shift) ^ ((fiEnable && (5933 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_30_io_in_control_0_dataflow_b <=( _mesh_17_30_io_out_control_0_dataflow) ^ ((fiEnable && (5934 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_30_io_in_control_0_propagate_b <=( _mesh_17_30_io_out_control_0_propagate) ^ ((fiEnable && (5935 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_30_io_out_valid_0) begin
			b_979_0 <=( _mesh_18_30_io_out_b_0) ^ ((fiEnable && (5936 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2003_0 <=( _mesh_18_30_io_out_c_0) ^ ((fiEnable && (5937 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_30_io_in_control_0_shift_b <=( _mesh_18_30_io_out_control_0_shift) ^ ((fiEnable && (5938 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_30_io_in_control_0_dataflow_b <=( _mesh_18_30_io_out_control_0_dataflow) ^ ((fiEnable && (5939 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_30_io_in_control_0_propagate_b <=( _mesh_18_30_io_out_control_0_propagate) ^ ((fiEnable && (5940 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_30_io_out_valid_0) begin
			b_980_0 <=( _mesh_19_30_io_out_b_0) ^ ((fiEnable && (5941 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2004_0 <=( _mesh_19_30_io_out_c_0) ^ ((fiEnable && (5942 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_30_io_in_control_0_shift_b <=( _mesh_19_30_io_out_control_0_shift) ^ ((fiEnable && (5943 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_30_io_in_control_0_dataflow_b <=( _mesh_19_30_io_out_control_0_dataflow) ^ ((fiEnable && (5944 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_30_io_in_control_0_propagate_b <=( _mesh_19_30_io_out_control_0_propagate) ^ ((fiEnable && (5945 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_30_io_out_valid_0) begin
			b_981_0 <=( _mesh_20_30_io_out_b_0) ^ ((fiEnable && (5946 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2005_0 <=( _mesh_20_30_io_out_c_0) ^ ((fiEnable && (5947 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_30_io_in_control_0_shift_b <=( _mesh_20_30_io_out_control_0_shift) ^ ((fiEnable && (5948 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_30_io_in_control_0_dataflow_b <=( _mesh_20_30_io_out_control_0_dataflow) ^ ((fiEnable && (5949 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_30_io_in_control_0_propagate_b <=( _mesh_20_30_io_out_control_0_propagate) ^ ((fiEnable && (5950 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_30_io_out_valid_0) begin
			b_982_0 <=( _mesh_21_30_io_out_b_0) ^ ((fiEnable && (5951 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2006_0 <=( _mesh_21_30_io_out_c_0) ^ ((fiEnable && (5952 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_30_io_in_control_0_shift_b <=( _mesh_21_30_io_out_control_0_shift) ^ ((fiEnable && (5953 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_30_io_in_control_0_dataflow_b <=( _mesh_21_30_io_out_control_0_dataflow) ^ ((fiEnable && (5954 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_30_io_in_control_0_propagate_b <=( _mesh_21_30_io_out_control_0_propagate) ^ ((fiEnable && (5955 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_30_io_out_valid_0) begin
			b_983_0 <=( _mesh_22_30_io_out_b_0) ^ ((fiEnable && (5956 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2007_0 <=( _mesh_22_30_io_out_c_0) ^ ((fiEnable && (5957 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_30_io_in_control_0_shift_b <=( _mesh_22_30_io_out_control_0_shift) ^ ((fiEnable && (5958 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_30_io_in_control_0_dataflow_b <=( _mesh_22_30_io_out_control_0_dataflow) ^ ((fiEnable && (5959 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_30_io_in_control_0_propagate_b <=( _mesh_22_30_io_out_control_0_propagate) ^ ((fiEnable && (5960 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_30_io_out_valid_0) begin
			b_984_0 <=( _mesh_23_30_io_out_b_0) ^ ((fiEnable && (5961 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2008_0 <=( _mesh_23_30_io_out_c_0) ^ ((fiEnable && (5962 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_30_io_in_control_0_shift_b <=( _mesh_23_30_io_out_control_0_shift) ^ ((fiEnable && (5963 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_30_io_in_control_0_dataflow_b <=( _mesh_23_30_io_out_control_0_dataflow) ^ ((fiEnable && (5964 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_30_io_in_control_0_propagate_b <=( _mesh_23_30_io_out_control_0_propagate) ^ ((fiEnable && (5965 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_30_io_out_valid_0) begin
			b_985_0 <=( _mesh_24_30_io_out_b_0) ^ ((fiEnable && (5966 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2009_0 <=( _mesh_24_30_io_out_c_0) ^ ((fiEnable && (5967 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_30_io_in_control_0_shift_b <=( _mesh_24_30_io_out_control_0_shift) ^ ((fiEnable && (5968 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_30_io_in_control_0_dataflow_b <=( _mesh_24_30_io_out_control_0_dataflow) ^ ((fiEnable && (5969 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_30_io_in_control_0_propagate_b <=( _mesh_24_30_io_out_control_0_propagate) ^ ((fiEnable && (5970 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_30_io_out_valid_0) begin
			b_986_0 <=( _mesh_25_30_io_out_b_0) ^ ((fiEnable && (5971 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2010_0 <=( _mesh_25_30_io_out_c_0) ^ ((fiEnable && (5972 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_30_io_in_control_0_shift_b <=( _mesh_25_30_io_out_control_0_shift) ^ ((fiEnable && (5973 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_30_io_in_control_0_dataflow_b <=( _mesh_25_30_io_out_control_0_dataflow) ^ ((fiEnable && (5974 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_30_io_in_control_0_propagate_b <=( _mesh_25_30_io_out_control_0_propagate) ^ ((fiEnable && (5975 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_30_io_out_valid_0) begin
			b_987_0 <=( _mesh_26_30_io_out_b_0) ^ ((fiEnable && (5976 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2011_0 <=( _mesh_26_30_io_out_c_0) ^ ((fiEnable && (5977 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_30_io_in_control_0_shift_b <=( _mesh_26_30_io_out_control_0_shift) ^ ((fiEnable && (5978 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_30_io_in_control_0_dataflow_b <=( _mesh_26_30_io_out_control_0_dataflow) ^ ((fiEnable && (5979 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_30_io_in_control_0_propagate_b <=( _mesh_26_30_io_out_control_0_propagate) ^ ((fiEnable && (5980 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_30_io_out_valid_0) begin
			b_988_0 <=( _mesh_27_30_io_out_b_0) ^ ((fiEnable && (5981 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2012_0 <=( _mesh_27_30_io_out_c_0) ^ ((fiEnable && (5982 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_30_io_in_control_0_shift_b <=( _mesh_27_30_io_out_control_0_shift) ^ ((fiEnable && (5983 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_30_io_in_control_0_dataflow_b <=( _mesh_27_30_io_out_control_0_dataflow) ^ ((fiEnable && (5984 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_30_io_in_control_0_propagate_b <=( _mesh_27_30_io_out_control_0_propagate) ^ ((fiEnable && (5985 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_30_io_out_valid_0) begin
			b_989_0 <=( _mesh_28_30_io_out_b_0) ^ ((fiEnable && (5986 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2013_0 <=( _mesh_28_30_io_out_c_0) ^ ((fiEnable && (5987 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_30_io_in_control_0_shift_b <=( _mesh_28_30_io_out_control_0_shift) ^ ((fiEnable && (5988 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_30_io_in_control_0_dataflow_b <=( _mesh_28_30_io_out_control_0_dataflow) ^ ((fiEnable && (5989 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_30_io_in_control_0_propagate_b <=( _mesh_28_30_io_out_control_0_propagate) ^ ((fiEnable && (5990 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_30_io_out_valid_0) begin
			b_990_0 <=( _mesh_29_30_io_out_b_0) ^ ((fiEnable && (5991 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2014_0 <=( _mesh_29_30_io_out_c_0) ^ ((fiEnable && (5992 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_30_io_in_control_0_shift_b <=( _mesh_29_30_io_out_control_0_shift) ^ ((fiEnable && (5993 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_30_io_in_control_0_dataflow_b <=( _mesh_29_30_io_out_control_0_dataflow) ^ ((fiEnable && (5994 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_30_io_in_control_0_propagate_b <=( _mesh_29_30_io_out_control_0_propagate) ^ ((fiEnable && (5995 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_30_io_out_valid_0) begin
			b_991_0 <=( _mesh_30_30_io_out_b_0) ^ ((fiEnable && (5996 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2015_0 <=( _mesh_30_30_io_out_c_0) ^ ((fiEnable && (5997 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_30_io_in_control_0_shift_b <=( _mesh_30_30_io_out_control_0_shift) ^ ((fiEnable && (5998 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_30_io_in_control_0_dataflow_b <=( _mesh_30_30_io_out_control_0_dataflow) ^ ((fiEnable && (5999 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_30_io_in_control_0_propagate_b <=( _mesh_30_30_io_out_control_0_propagate) ^ ((fiEnable && (6000 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_31_0) begin
			b_992_0 <=( io_in_b_31_0) ^ ((fiEnable && (6001 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2016_0 <=( io_in_d_31_0) ^ ((fiEnable && (6002 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_31_io_in_control_0_shift_b <=( io_in_control_31_0_shift) ^ ((fiEnable && (6003 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_31_io_in_control_0_dataflow_b <=( io_in_control_31_0_dataflow) ^ ((fiEnable && (6004 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_31_io_in_control_0_propagate_b <=( io_in_control_31_0_propagate) ^ ((fiEnable && (6005 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_31_io_out_valid_0) begin
			b_993_0 <=( _mesh_0_31_io_out_b_0) ^ ((fiEnable && (6006 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2017_0 <=( _mesh_0_31_io_out_c_0) ^ ((fiEnable && (6007 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_31_io_in_control_0_shift_b <=( _mesh_0_31_io_out_control_0_shift) ^ ((fiEnable && (6008 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_31_io_in_control_0_dataflow_b <=( _mesh_0_31_io_out_control_0_dataflow) ^ ((fiEnable && (6009 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_31_io_in_control_0_propagate_b <=( _mesh_0_31_io_out_control_0_propagate) ^ ((fiEnable && (6010 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_31_io_out_valid_0) begin
			b_994_0 <=( _mesh_1_31_io_out_b_0) ^ ((fiEnable && (6011 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2018_0 <=( _mesh_1_31_io_out_c_0) ^ ((fiEnable && (6012 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_31_io_in_control_0_shift_b <=( _mesh_1_31_io_out_control_0_shift) ^ ((fiEnable && (6013 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_31_io_in_control_0_dataflow_b <=( _mesh_1_31_io_out_control_0_dataflow) ^ ((fiEnable && (6014 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_31_io_in_control_0_propagate_b <=( _mesh_1_31_io_out_control_0_propagate) ^ ((fiEnable && (6015 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_31_io_out_valid_0) begin
			b_995_0 <=( _mesh_2_31_io_out_b_0) ^ ((fiEnable && (6016 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2019_0 <=( _mesh_2_31_io_out_c_0) ^ ((fiEnable && (6017 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_31_io_in_control_0_shift_b <=( _mesh_2_31_io_out_control_0_shift) ^ ((fiEnable && (6018 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_31_io_in_control_0_dataflow_b <=( _mesh_2_31_io_out_control_0_dataflow) ^ ((fiEnable && (6019 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_31_io_in_control_0_propagate_b <=( _mesh_2_31_io_out_control_0_propagate) ^ ((fiEnable && (6020 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_31_io_out_valid_0) begin
			b_996_0 <=( _mesh_3_31_io_out_b_0) ^ ((fiEnable && (6021 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2020_0 <=( _mesh_3_31_io_out_c_0) ^ ((fiEnable && (6022 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_31_io_in_control_0_shift_b <=( _mesh_3_31_io_out_control_0_shift) ^ ((fiEnable && (6023 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_31_io_in_control_0_dataflow_b <=( _mesh_3_31_io_out_control_0_dataflow) ^ ((fiEnable && (6024 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_31_io_in_control_0_propagate_b <=( _mesh_3_31_io_out_control_0_propagate) ^ ((fiEnable && (6025 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_31_io_out_valid_0) begin
			b_997_0 <=( _mesh_4_31_io_out_b_0) ^ ((fiEnable && (6026 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2021_0 <=( _mesh_4_31_io_out_c_0) ^ ((fiEnable && (6027 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_31_io_in_control_0_shift_b <=( _mesh_4_31_io_out_control_0_shift) ^ ((fiEnable && (6028 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_31_io_in_control_0_dataflow_b <=( _mesh_4_31_io_out_control_0_dataflow) ^ ((fiEnable && (6029 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_31_io_in_control_0_propagate_b <=( _mesh_4_31_io_out_control_0_propagate) ^ ((fiEnable && (6030 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_31_io_out_valid_0) begin
			b_998_0 <=( _mesh_5_31_io_out_b_0) ^ ((fiEnable && (6031 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2022_0 <=( _mesh_5_31_io_out_c_0) ^ ((fiEnable && (6032 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_31_io_in_control_0_shift_b <=( _mesh_5_31_io_out_control_0_shift) ^ ((fiEnable && (6033 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_31_io_in_control_0_dataflow_b <=( _mesh_5_31_io_out_control_0_dataflow) ^ ((fiEnable && (6034 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_31_io_in_control_0_propagate_b <=( _mesh_5_31_io_out_control_0_propagate) ^ ((fiEnable && (6035 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_31_io_out_valid_0) begin
			b_999_0 <=( _mesh_6_31_io_out_b_0) ^ ((fiEnable && (6036 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2023_0 <=( _mesh_6_31_io_out_c_0) ^ ((fiEnable && (6037 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_31_io_in_control_0_shift_b <=( _mesh_6_31_io_out_control_0_shift) ^ ((fiEnable && (6038 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_31_io_in_control_0_dataflow_b <=( _mesh_6_31_io_out_control_0_dataflow) ^ ((fiEnable && (6039 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_31_io_in_control_0_propagate_b <=( _mesh_6_31_io_out_control_0_propagate) ^ ((fiEnable && (6040 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_7_31_io_out_valid_0) begin
			b_1000_0 <=( _mesh_7_31_io_out_b_0) ^ ((fiEnable && (6041 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2024_0 <=( _mesh_7_31_io_out_c_0) ^ ((fiEnable && (6042 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_8_31_io_in_control_0_shift_b <=( _mesh_7_31_io_out_control_0_shift) ^ ((fiEnable && (6043 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_8_31_io_in_control_0_dataflow_b <=( _mesh_7_31_io_out_control_0_dataflow) ^ ((fiEnable && (6044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_8_31_io_in_control_0_propagate_b <=( _mesh_7_31_io_out_control_0_propagate) ^ ((fiEnable && (6045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_8_31_io_out_valid_0) begin
			b_1001_0 <=( _mesh_8_31_io_out_b_0) ^ ((fiEnable && (6046 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2025_0 <=( _mesh_8_31_io_out_c_0) ^ ((fiEnable && (6047 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_9_31_io_in_control_0_shift_b <=( _mesh_8_31_io_out_control_0_shift) ^ ((fiEnable && (6048 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_9_31_io_in_control_0_dataflow_b <=( _mesh_8_31_io_out_control_0_dataflow) ^ ((fiEnable && (6049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_9_31_io_in_control_0_propagate_b <=( _mesh_8_31_io_out_control_0_propagate) ^ ((fiEnable && (6050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_9_31_io_out_valid_0) begin
			b_1002_0 <=( _mesh_9_31_io_out_b_0) ^ ((fiEnable && (6051 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2026_0 <=( _mesh_9_31_io_out_c_0) ^ ((fiEnable && (6052 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_10_31_io_in_control_0_shift_b <=( _mesh_9_31_io_out_control_0_shift) ^ ((fiEnable && (6053 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_10_31_io_in_control_0_dataflow_b <=( _mesh_9_31_io_out_control_0_dataflow) ^ ((fiEnable && (6054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_10_31_io_in_control_0_propagate_b <=( _mesh_9_31_io_out_control_0_propagate) ^ ((fiEnable && (6055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_10_31_io_out_valid_0) begin
			b_1003_0 <=( _mesh_10_31_io_out_b_0) ^ ((fiEnable && (6056 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2027_0 <=( _mesh_10_31_io_out_c_0) ^ ((fiEnable && (6057 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_11_31_io_in_control_0_shift_b <=( _mesh_10_31_io_out_control_0_shift) ^ ((fiEnable && (6058 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_11_31_io_in_control_0_dataflow_b <=( _mesh_10_31_io_out_control_0_dataflow) ^ ((fiEnable && (6059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_11_31_io_in_control_0_propagate_b <=( _mesh_10_31_io_out_control_0_propagate) ^ ((fiEnable && (6060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_11_31_io_out_valid_0) begin
			b_1004_0 <=( _mesh_11_31_io_out_b_0) ^ ((fiEnable && (6061 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2028_0 <=( _mesh_11_31_io_out_c_0) ^ ((fiEnable && (6062 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_12_31_io_in_control_0_shift_b <=( _mesh_11_31_io_out_control_0_shift) ^ ((fiEnable && (6063 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_12_31_io_in_control_0_dataflow_b <=( _mesh_11_31_io_out_control_0_dataflow) ^ ((fiEnable && (6064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_12_31_io_in_control_0_propagate_b <=( _mesh_11_31_io_out_control_0_propagate) ^ ((fiEnable && (6065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_12_31_io_out_valid_0) begin
			b_1005_0 <=( _mesh_12_31_io_out_b_0) ^ ((fiEnable && (6066 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2029_0 <=( _mesh_12_31_io_out_c_0) ^ ((fiEnable && (6067 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_13_31_io_in_control_0_shift_b <=( _mesh_12_31_io_out_control_0_shift) ^ ((fiEnable && (6068 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_13_31_io_in_control_0_dataflow_b <=( _mesh_12_31_io_out_control_0_dataflow) ^ ((fiEnable && (6069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_13_31_io_in_control_0_propagate_b <=( _mesh_12_31_io_out_control_0_propagate) ^ ((fiEnable && (6070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_13_31_io_out_valid_0) begin
			b_1006_0 <=( _mesh_13_31_io_out_b_0) ^ ((fiEnable && (6071 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2030_0 <=( _mesh_13_31_io_out_c_0) ^ ((fiEnable && (6072 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_14_31_io_in_control_0_shift_b <=( _mesh_13_31_io_out_control_0_shift) ^ ((fiEnable && (6073 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_14_31_io_in_control_0_dataflow_b <=( _mesh_13_31_io_out_control_0_dataflow) ^ ((fiEnable && (6074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_14_31_io_in_control_0_propagate_b <=( _mesh_13_31_io_out_control_0_propagate) ^ ((fiEnable && (6075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_14_31_io_out_valid_0) begin
			b_1007_0 <=( _mesh_14_31_io_out_b_0) ^ ((fiEnable && (6076 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2031_0 <=( _mesh_14_31_io_out_c_0) ^ ((fiEnable && (6077 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_15_31_io_in_control_0_shift_b <=( _mesh_14_31_io_out_control_0_shift) ^ ((fiEnable && (6078 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_15_31_io_in_control_0_dataflow_b <=( _mesh_14_31_io_out_control_0_dataflow) ^ ((fiEnable && (6079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_15_31_io_in_control_0_propagate_b <=( _mesh_14_31_io_out_control_0_propagate) ^ ((fiEnable && (6080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_15_31_io_out_valid_0) begin
			b_1008_0 <=( _mesh_15_31_io_out_b_0) ^ ((fiEnable && (6081 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2032_0 <=( _mesh_15_31_io_out_c_0) ^ ((fiEnable && (6082 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_16_31_io_in_control_0_shift_b <=( _mesh_15_31_io_out_control_0_shift) ^ ((fiEnable && (6083 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_16_31_io_in_control_0_dataflow_b <=( _mesh_15_31_io_out_control_0_dataflow) ^ ((fiEnable && (6084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_16_31_io_in_control_0_propagate_b <=( _mesh_15_31_io_out_control_0_propagate) ^ ((fiEnable && (6085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_16_31_io_out_valid_0) begin
			b_1009_0 <=( _mesh_16_31_io_out_b_0) ^ ((fiEnable && (6086 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2033_0 <=( _mesh_16_31_io_out_c_0) ^ ((fiEnable && (6087 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_17_31_io_in_control_0_shift_b <=( _mesh_16_31_io_out_control_0_shift) ^ ((fiEnable && (6088 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_17_31_io_in_control_0_dataflow_b <=( _mesh_16_31_io_out_control_0_dataflow) ^ ((fiEnable && (6089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_17_31_io_in_control_0_propagate_b <=( _mesh_16_31_io_out_control_0_propagate) ^ ((fiEnable && (6090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_17_31_io_out_valid_0) begin
			b_1010_0 <=( _mesh_17_31_io_out_b_0) ^ ((fiEnable && (6091 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2034_0 <=( _mesh_17_31_io_out_c_0) ^ ((fiEnable && (6092 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_18_31_io_in_control_0_shift_b <=( _mesh_17_31_io_out_control_0_shift) ^ ((fiEnable && (6093 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_18_31_io_in_control_0_dataflow_b <=( _mesh_17_31_io_out_control_0_dataflow) ^ ((fiEnable && (6094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_18_31_io_in_control_0_propagate_b <=( _mesh_17_31_io_out_control_0_propagate) ^ ((fiEnable && (6095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_18_31_io_out_valid_0) begin
			b_1011_0 <=( _mesh_18_31_io_out_b_0) ^ ((fiEnable && (6096 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2035_0 <=( _mesh_18_31_io_out_c_0) ^ ((fiEnable && (6097 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_19_31_io_in_control_0_shift_b <=( _mesh_18_31_io_out_control_0_shift) ^ ((fiEnable && (6098 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_19_31_io_in_control_0_dataflow_b <=( _mesh_18_31_io_out_control_0_dataflow) ^ ((fiEnable && (6099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_19_31_io_in_control_0_propagate_b <=( _mesh_18_31_io_out_control_0_propagate) ^ ((fiEnable && (6100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_19_31_io_out_valid_0) begin
			b_1012_0 <=( _mesh_19_31_io_out_b_0) ^ ((fiEnable && (6101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2036_0 <=( _mesh_19_31_io_out_c_0) ^ ((fiEnable && (6102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_20_31_io_in_control_0_shift_b <=( _mesh_19_31_io_out_control_0_shift) ^ ((fiEnable && (6103 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_20_31_io_in_control_0_dataflow_b <=( _mesh_19_31_io_out_control_0_dataflow) ^ ((fiEnable && (6104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_20_31_io_in_control_0_propagate_b <=( _mesh_19_31_io_out_control_0_propagate) ^ ((fiEnable && (6105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_20_31_io_out_valid_0) begin
			b_1013_0 <=( _mesh_20_31_io_out_b_0) ^ ((fiEnable && (6106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2037_0 <=( _mesh_20_31_io_out_c_0) ^ ((fiEnable && (6107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_21_31_io_in_control_0_shift_b <=( _mesh_20_31_io_out_control_0_shift) ^ ((fiEnable && (6108 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_21_31_io_in_control_0_dataflow_b <=( _mesh_20_31_io_out_control_0_dataflow) ^ ((fiEnable && (6109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_21_31_io_in_control_0_propagate_b <=( _mesh_20_31_io_out_control_0_propagate) ^ ((fiEnable && (6110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_21_31_io_out_valid_0) begin
			b_1014_0 <=( _mesh_21_31_io_out_b_0) ^ ((fiEnable && (6111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2038_0 <=( _mesh_21_31_io_out_c_0) ^ ((fiEnable && (6112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_22_31_io_in_control_0_shift_b <=( _mesh_21_31_io_out_control_0_shift) ^ ((fiEnable && (6113 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_22_31_io_in_control_0_dataflow_b <=( _mesh_21_31_io_out_control_0_dataflow) ^ ((fiEnable && (6114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_22_31_io_in_control_0_propagate_b <=( _mesh_21_31_io_out_control_0_propagate) ^ ((fiEnable && (6115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_22_31_io_out_valid_0) begin
			b_1015_0 <=( _mesh_22_31_io_out_b_0) ^ ((fiEnable && (6116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2039_0 <=( _mesh_22_31_io_out_c_0) ^ ((fiEnable && (6117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_23_31_io_in_control_0_shift_b <=( _mesh_22_31_io_out_control_0_shift) ^ ((fiEnable && (6118 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_23_31_io_in_control_0_dataflow_b <=( _mesh_22_31_io_out_control_0_dataflow) ^ ((fiEnable && (6119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_23_31_io_in_control_0_propagate_b <=( _mesh_22_31_io_out_control_0_propagate) ^ ((fiEnable && (6120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_23_31_io_out_valid_0) begin
			b_1016_0 <=( _mesh_23_31_io_out_b_0) ^ ((fiEnable && (6121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2040_0 <=( _mesh_23_31_io_out_c_0) ^ ((fiEnable && (6122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_24_31_io_in_control_0_shift_b <=( _mesh_23_31_io_out_control_0_shift) ^ ((fiEnable && (6123 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_24_31_io_in_control_0_dataflow_b <=( _mesh_23_31_io_out_control_0_dataflow) ^ ((fiEnable && (6124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_24_31_io_in_control_0_propagate_b <=( _mesh_23_31_io_out_control_0_propagate) ^ ((fiEnable && (6125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_24_31_io_out_valid_0) begin
			b_1017_0 <=( _mesh_24_31_io_out_b_0) ^ ((fiEnable && (6126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2041_0 <=( _mesh_24_31_io_out_c_0) ^ ((fiEnable && (6127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_25_31_io_in_control_0_shift_b <=( _mesh_24_31_io_out_control_0_shift) ^ ((fiEnable && (6128 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_25_31_io_in_control_0_dataflow_b <=( _mesh_24_31_io_out_control_0_dataflow) ^ ((fiEnable && (6129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_25_31_io_in_control_0_propagate_b <=( _mesh_24_31_io_out_control_0_propagate) ^ ((fiEnable && (6130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_25_31_io_out_valid_0) begin
			b_1018_0 <=( _mesh_25_31_io_out_b_0) ^ ((fiEnable && (6131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2042_0 <=( _mesh_25_31_io_out_c_0) ^ ((fiEnable && (6132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_26_31_io_in_control_0_shift_b <=( _mesh_25_31_io_out_control_0_shift) ^ ((fiEnable && (6133 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_26_31_io_in_control_0_dataflow_b <=( _mesh_25_31_io_out_control_0_dataflow) ^ ((fiEnable && (6134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_26_31_io_in_control_0_propagate_b <=( _mesh_25_31_io_out_control_0_propagate) ^ ((fiEnable && (6135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_26_31_io_out_valid_0) begin
			b_1019_0 <=( _mesh_26_31_io_out_b_0) ^ ((fiEnable && (6136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2043_0 <=( _mesh_26_31_io_out_c_0) ^ ((fiEnable && (6137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_27_31_io_in_control_0_shift_b <=( _mesh_26_31_io_out_control_0_shift) ^ ((fiEnable && (6138 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_27_31_io_in_control_0_dataflow_b <=( _mesh_26_31_io_out_control_0_dataflow) ^ ((fiEnable && (6139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_27_31_io_in_control_0_propagate_b <=( _mesh_26_31_io_out_control_0_propagate) ^ ((fiEnable && (6140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_27_31_io_out_valid_0) begin
			b_1020_0 <=( _mesh_27_31_io_out_b_0) ^ ((fiEnable && (6141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2044_0 <=( _mesh_27_31_io_out_c_0) ^ ((fiEnable && (6142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_28_31_io_in_control_0_shift_b <=( _mesh_27_31_io_out_control_0_shift) ^ ((fiEnable && (6143 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_28_31_io_in_control_0_dataflow_b <=( _mesh_27_31_io_out_control_0_dataflow) ^ ((fiEnable && (6144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_28_31_io_in_control_0_propagate_b <=( _mesh_27_31_io_out_control_0_propagate) ^ ((fiEnable && (6145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_28_31_io_out_valid_0) begin
			b_1021_0 <=( _mesh_28_31_io_out_b_0) ^ ((fiEnable && (6146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2045_0 <=( _mesh_28_31_io_out_c_0) ^ ((fiEnable && (6147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_29_31_io_in_control_0_shift_b <=( _mesh_28_31_io_out_control_0_shift) ^ ((fiEnable && (6148 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_29_31_io_in_control_0_dataflow_b <=( _mesh_28_31_io_out_control_0_dataflow) ^ ((fiEnable && (6149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_29_31_io_in_control_0_propagate_b <=( _mesh_28_31_io_out_control_0_propagate) ^ ((fiEnable && (6150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_29_31_io_out_valid_0) begin
			b_1022_0 <=( _mesh_29_31_io_out_b_0) ^ ((fiEnable && (6151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2046_0 <=( _mesh_29_31_io_out_c_0) ^ ((fiEnable && (6152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_30_31_io_in_control_0_shift_b <=( _mesh_29_31_io_out_control_0_shift) ^ ((fiEnable && (6153 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_30_31_io_in_control_0_dataflow_b <=( _mesh_29_31_io_out_control_0_dataflow) ^ ((fiEnable && (6154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_30_31_io_in_control_0_propagate_b <=( _mesh_29_31_io_out_control_0_propagate) ^ ((fiEnable && (6155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_30_31_io_out_valid_0) begin
			b_1023_0 <=( _mesh_30_31_io_out_b_0) ^ ((fiEnable && (6156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_2047_0 <=( _mesh_30_31_io_out_c_0) ^ ((fiEnable && (6157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_31_31_io_in_control_0_shift_b <=( _mesh_30_31_io_out_control_0_shift) ^ ((fiEnable && (6158 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_31_31_io_in_control_0_dataflow_b <=( _mesh_30_31_io_out_control_0_dataflow) ^ ((fiEnable && (6159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_31_31_io_in_control_0_propagate_b <=( _mesh_30_31_io_out_control_0_propagate) ^ ((fiEnable && (6160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		r_1024_0 <=( io_in_valid_0_0) ^ ((fiEnable && (6161 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1025_0 <=( _mesh_0_0_io_out_valid_0) ^ ((fiEnable && (6162 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1026_0 <=( _mesh_1_0_io_out_valid_0) ^ ((fiEnable && (6163 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1027_0 <=( _mesh_2_0_io_out_valid_0) ^ ((fiEnable && (6164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1028_0 <=( _mesh_3_0_io_out_valid_0) ^ ((fiEnable && (6165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1029_0 <=( _mesh_4_0_io_out_valid_0) ^ ((fiEnable && (6166 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1030_0 <=( _mesh_5_0_io_out_valid_0) ^ ((fiEnable && (6167 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1031_0 <=( _mesh_6_0_io_out_valid_0) ^ ((fiEnable && (6168 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1032_0 <=( _mesh_7_0_io_out_valid_0) ^ ((fiEnable && (6169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1033_0 <=( _mesh_8_0_io_out_valid_0) ^ ((fiEnable && (6170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1034_0 <=( _mesh_9_0_io_out_valid_0) ^ ((fiEnable && (6171 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1035_0 <=( _mesh_10_0_io_out_valid_0) ^ ((fiEnable && (6172 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1036_0 <=( _mesh_11_0_io_out_valid_0) ^ ((fiEnable && (6173 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1037_0 <=( _mesh_12_0_io_out_valid_0) ^ ((fiEnable && (6174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1038_0 <=( _mesh_13_0_io_out_valid_0) ^ ((fiEnable && (6175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1039_0 <=( _mesh_14_0_io_out_valid_0) ^ ((fiEnable && (6176 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1040_0 <=( _mesh_15_0_io_out_valid_0) ^ ((fiEnable && (6177 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1041_0 <=( _mesh_16_0_io_out_valid_0) ^ ((fiEnable && (6178 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1042_0 <=( _mesh_17_0_io_out_valid_0) ^ ((fiEnable && (6179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1043_0 <=( _mesh_18_0_io_out_valid_0) ^ ((fiEnable && (6180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1044_0 <=( _mesh_19_0_io_out_valid_0) ^ ((fiEnable && (6181 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1045_0 <=( _mesh_20_0_io_out_valid_0) ^ ((fiEnable && (6182 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1046_0 <=( _mesh_21_0_io_out_valid_0) ^ ((fiEnable && (6183 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1047_0 <=( _mesh_22_0_io_out_valid_0) ^ ((fiEnable && (6184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1048_0 <=( _mesh_23_0_io_out_valid_0) ^ ((fiEnable && (6185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1049_0 <=( _mesh_24_0_io_out_valid_0) ^ ((fiEnable && (6186 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1050_0 <=( _mesh_25_0_io_out_valid_0) ^ ((fiEnable && (6187 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1051_0 <=( _mesh_26_0_io_out_valid_0) ^ ((fiEnable && (6188 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1052_0 <=( _mesh_27_0_io_out_valid_0) ^ ((fiEnable && (6189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1053_0 <=( _mesh_28_0_io_out_valid_0) ^ ((fiEnable && (6190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1054_0 <=( _mesh_29_0_io_out_valid_0) ^ ((fiEnable && (6191 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1055_0 <=( _mesh_30_0_io_out_valid_0) ^ ((fiEnable && (6192 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1056_0 <=( io_in_valid_1_0) ^ ((fiEnable && (6193 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1057_0 <=( _mesh_0_1_io_out_valid_0) ^ ((fiEnable && (6194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1058_0 <=( _mesh_1_1_io_out_valid_0) ^ ((fiEnable && (6195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1059_0 <=( _mesh_2_1_io_out_valid_0) ^ ((fiEnable && (6196 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1060_0 <=( _mesh_3_1_io_out_valid_0) ^ ((fiEnable && (6197 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1061_0 <=( _mesh_4_1_io_out_valid_0) ^ ((fiEnable && (6198 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1062_0 <=( _mesh_5_1_io_out_valid_0) ^ ((fiEnable && (6199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1063_0 <=( _mesh_6_1_io_out_valid_0) ^ ((fiEnable && (6200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1064_0 <=( _mesh_7_1_io_out_valid_0) ^ ((fiEnable && (6201 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1065_0 <=( _mesh_8_1_io_out_valid_0) ^ ((fiEnable && (6202 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1066_0 <=( _mesh_9_1_io_out_valid_0) ^ ((fiEnable && (6203 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1067_0 <=( _mesh_10_1_io_out_valid_0) ^ ((fiEnable && (6204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1068_0 <=( _mesh_11_1_io_out_valid_0) ^ ((fiEnable && (6205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1069_0 <=( _mesh_12_1_io_out_valid_0) ^ ((fiEnable && (6206 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1070_0 <=( _mesh_13_1_io_out_valid_0) ^ ((fiEnable && (6207 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1071_0 <=( _mesh_14_1_io_out_valid_0) ^ ((fiEnable && (6208 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1072_0 <=( _mesh_15_1_io_out_valid_0) ^ ((fiEnable && (6209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1073_0 <=( _mesh_16_1_io_out_valid_0) ^ ((fiEnable && (6210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1074_0 <=( _mesh_17_1_io_out_valid_0) ^ ((fiEnable && (6211 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1075_0 <=( _mesh_18_1_io_out_valid_0) ^ ((fiEnable && (6212 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1076_0 <=( _mesh_19_1_io_out_valid_0) ^ ((fiEnable && (6213 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1077_0 <=( _mesh_20_1_io_out_valid_0) ^ ((fiEnable && (6214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1078_0 <=( _mesh_21_1_io_out_valid_0) ^ ((fiEnable && (6215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1079_0 <=( _mesh_22_1_io_out_valid_0) ^ ((fiEnable && (6216 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1080_0 <=( _mesh_23_1_io_out_valid_0) ^ ((fiEnable && (6217 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1081_0 <=( _mesh_24_1_io_out_valid_0) ^ ((fiEnable && (6218 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1082_0 <=( _mesh_25_1_io_out_valid_0) ^ ((fiEnable && (6219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1083_0 <=( _mesh_26_1_io_out_valid_0) ^ ((fiEnable && (6220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1084_0 <=( _mesh_27_1_io_out_valid_0) ^ ((fiEnable && (6221 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1085_0 <=( _mesh_28_1_io_out_valid_0) ^ ((fiEnable && (6222 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1086_0 <=( _mesh_29_1_io_out_valid_0) ^ ((fiEnable && (6223 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1087_0 <=( _mesh_30_1_io_out_valid_0) ^ ((fiEnable && (6224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1088_0 <=( io_in_valid_2_0) ^ ((fiEnable && (6225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1089_0 <=( _mesh_0_2_io_out_valid_0) ^ ((fiEnable && (6226 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1090_0 <=( _mesh_1_2_io_out_valid_0) ^ ((fiEnable && (6227 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1091_0 <=( _mesh_2_2_io_out_valid_0) ^ ((fiEnable && (6228 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1092_0 <=( _mesh_3_2_io_out_valid_0) ^ ((fiEnable && (6229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1093_0 <=( _mesh_4_2_io_out_valid_0) ^ ((fiEnable && (6230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1094_0 <=( _mesh_5_2_io_out_valid_0) ^ ((fiEnable && (6231 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1095_0 <=( _mesh_6_2_io_out_valid_0) ^ ((fiEnable && (6232 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1096_0 <=( _mesh_7_2_io_out_valid_0) ^ ((fiEnable && (6233 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1097_0 <=( _mesh_8_2_io_out_valid_0) ^ ((fiEnable && (6234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1098_0 <=( _mesh_9_2_io_out_valid_0) ^ ((fiEnable && (6235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1099_0 <=( _mesh_10_2_io_out_valid_0) ^ ((fiEnable && (6236 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1100_0 <=( _mesh_11_2_io_out_valid_0) ^ ((fiEnable && (6237 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1101_0 <=( _mesh_12_2_io_out_valid_0) ^ ((fiEnable && (6238 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1102_0 <=( _mesh_13_2_io_out_valid_0) ^ ((fiEnable && (6239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1103_0 <=( _mesh_14_2_io_out_valid_0) ^ ((fiEnable && (6240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1104_0 <=( _mesh_15_2_io_out_valid_0) ^ ((fiEnable && (6241 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1105_0 <=( _mesh_16_2_io_out_valid_0) ^ ((fiEnable && (6242 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1106_0 <=( _mesh_17_2_io_out_valid_0) ^ ((fiEnable && (6243 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1107_0 <=( _mesh_18_2_io_out_valid_0) ^ ((fiEnable && (6244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1108_0 <=( _mesh_19_2_io_out_valid_0) ^ ((fiEnable && (6245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1109_0 <=( _mesh_20_2_io_out_valid_0) ^ ((fiEnable && (6246 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1110_0 <=( _mesh_21_2_io_out_valid_0) ^ ((fiEnable && (6247 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1111_0 <=( _mesh_22_2_io_out_valid_0) ^ ((fiEnable && (6248 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1112_0 <=( _mesh_23_2_io_out_valid_0) ^ ((fiEnable && (6249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1113_0 <=( _mesh_24_2_io_out_valid_0) ^ ((fiEnable && (6250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1114_0 <=( _mesh_25_2_io_out_valid_0) ^ ((fiEnable && (6251 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1115_0 <=( _mesh_26_2_io_out_valid_0) ^ ((fiEnable && (6252 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1116_0 <=( _mesh_27_2_io_out_valid_0) ^ ((fiEnable && (6253 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1117_0 <=( _mesh_28_2_io_out_valid_0) ^ ((fiEnable && (6254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1118_0 <=( _mesh_29_2_io_out_valid_0) ^ ((fiEnable && (6255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1119_0 <=( _mesh_30_2_io_out_valid_0) ^ ((fiEnable && (6256 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1120_0 <=( io_in_valid_3_0) ^ ((fiEnable && (6257 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1121_0 <=( _mesh_0_3_io_out_valid_0) ^ ((fiEnable && (6258 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1122_0 <=( _mesh_1_3_io_out_valid_0) ^ ((fiEnable && (6259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1123_0 <=( _mesh_2_3_io_out_valid_0) ^ ((fiEnable && (6260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1124_0 <=( _mesh_3_3_io_out_valid_0) ^ ((fiEnable && (6261 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1125_0 <=( _mesh_4_3_io_out_valid_0) ^ ((fiEnable && (6262 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1126_0 <=( _mesh_5_3_io_out_valid_0) ^ ((fiEnable && (6263 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1127_0 <=( _mesh_6_3_io_out_valid_0) ^ ((fiEnable && (6264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1128_0 <=( _mesh_7_3_io_out_valid_0) ^ ((fiEnable && (6265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1129_0 <=( _mesh_8_3_io_out_valid_0) ^ ((fiEnable && (6266 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1130_0 <=( _mesh_9_3_io_out_valid_0) ^ ((fiEnable && (6267 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1131_0 <=( _mesh_10_3_io_out_valid_0) ^ ((fiEnable && (6268 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1132_0 <=( _mesh_11_3_io_out_valid_0) ^ ((fiEnable && (6269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1133_0 <=( _mesh_12_3_io_out_valid_0) ^ ((fiEnable && (6270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1134_0 <=( _mesh_13_3_io_out_valid_0) ^ ((fiEnable && (6271 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1135_0 <=( _mesh_14_3_io_out_valid_0) ^ ((fiEnable && (6272 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1136_0 <=( _mesh_15_3_io_out_valid_0) ^ ((fiEnable && (6273 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1137_0 <=( _mesh_16_3_io_out_valid_0) ^ ((fiEnable && (6274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1138_0 <=( _mesh_17_3_io_out_valid_0) ^ ((fiEnable && (6275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1139_0 <=( _mesh_18_3_io_out_valid_0) ^ ((fiEnable && (6276 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1140_0 <=( _mesh_19_3_io_out_valid_0) ^ ((fiEnable && (6277 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1141_0 <=( _mesh_20_3_io_out_valid_0) ^ ((fiEnable && (6278 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1142_0 <=( _mesh_21_3_io_out_valid_0) ^ ((fiEnable && (6279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1143_0 <=( _mesh_22_3_io_out_valid_0) ^ ((fiEnable && (6280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1144_0 <=( _mesh_23_3_io_out_valid_0) ^ ((fiEnable && (6281 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1145_0 <=( _mesh_24_3_io_out_valid_0) ^ ((fiEnable && (6282 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1146_0 <=( _mesh_25_3_io_out_valid_0) ^ ((fiEnable && (6283 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1147_0 <=( _mesh_26_3_io_out_valid_0) ^ ((fiEnable && (6284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1148_0 <=( _mesh_27_3_io_out_valid_0) ^ ((fiEnable && (6285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1149_0 <=( _mesh_28_3_io_out_valid_0) ^ ((fiEnable && (6286 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1150_0 <=( _mesh_29_3_io_out_valid_0) ^ ((fiEnable && (6287 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1151_0 <=( _mesh_30_3_io_out_valid_0) ^ ((fiEnable && (6288 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1152_0 <=( io_in_valid_4_0) ^ ((fiEnable && (6289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1153_0 <=( _mesh_0_4_io_out_valid_0) ^ ((fiEnable && (6290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1154_0 <=( _mesh_1_4_io_out_valid_0) ^ ((fiEnable && (6291 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1155_0 <=( _mesh_2_4_io_out_valid_0) ^ ((fiEnable && (6292 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1156_0 <=( _mesh_3_4_io_out_valid_0) ^ ((fiEnable && (6293 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1157_0 <=( _mesh_4_4_io_out_valid_0) ^ ((fiEnable && (6294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1158_0 <=( _mesh_5_4_io_out_valid_0) ^ ((fiEnable && (6295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1159_0 <=( _mesh_6_4_io_out_valid_0) ^ ((fiEnable && (6296 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1160_0 <=( _mesh_7_4_io_out_valid_0) ^ ((fiEnable && (6297 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1161_0 <=( _mesh_8_4_io_out_valid_0) ^ ((fiEnable && (6298 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1162_0 <=( _mesh_9_4_io_out_valid_0) ^ ((fiEnable && (6299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1163_0 <=( _mesh_10_4_io_out_valid_0) ^ ((fiEnable && (6300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1164_0 <=( _mesh_11_4_io_out_valid_0) ^ ((fiEnable && (6301 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1165_0 <=( _mesh_12_4_io_out_valid_0) ^ ((fiEnable && (6302 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1166_0 <=( _mesh_13_4_io_out_valid_0) ^ ((fiEnable && (6303 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1167_0 <=( _mesh_14_4_io_out_valid_0) ^ ((fiEnable && (6304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1168_0 <=( _mesh_15_4_io_out_valid_0) ^ ((fiEnable && (6305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1169_0 <=( _mesh_16_4_io_out_valid_0) ^ ((fiEnable && (6306 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1170_0 <=( _mesh_17_4_io_out_valid_0) ^ ((fiEnable && (6307 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1171_0 <=( _mesh_18_4_io_out_valid_0) ^ ((fiEnable && (6308 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1172_0 <=( _mesh_19_4_io_out_valid_0) ^ ((fiEnable && (6309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1173_0 <=( _mesh_20_4_io_out_valid_0) ^ ((fiEnable && (6310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1174_0 <=( _mesh_21_4_io_out_valid_0) ^ ((fiEnable && (6311 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1175_0 <=( _mesh_22_4_io_out_valid_0) ^ ((fiEnable && (6312 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1176_0 <=( _mesh_23_4_io_out_valid_0) ^ ((fiEnable && (6313 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1177_0 <=( _mesh_24_4_io_out_valid_0) ^ ((fiEnable && (6314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1178_0 <=( _mesh_25_4_io_out_valid_0) ^ ((fiEnable && (6315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1179_0 <=( _mesh_26_4_io_out_valid_0) ^ ((fiEnable && (6316 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1180_0 <=( _mesh_27_4_io_out_valid_0) ^ ((fiEnable && (6317 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1181_0 <=( _mesh_28_4_io_out_valid_0) ^ ((fiEnable && (6318 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1182_0 <=( _mesh_29_4_io_out_valid_0) ^ ((fiEnable && (6319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1183_0 <=( _mesh_30_4_io_out_valid_0) ^ ((fiEnable && (6320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1184_0 <=( io_in_valid_5_0) ^ ((fiEnable && (6321 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1185_0 <=( _mesh_0_5_io_out_valid_0) ^ ((fiEnable && (6322 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1186_0 <=( _mesh_1_5_io_out_valid_0) ^ ((fiEnable && (6323 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1187_0 <=( _mesh_2_5_io_out_valid_0) ^ ((fiEnable && (6324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1188_0 <=( _mesh_3_5_io_out_valid_0) ^ ((fiEnable && (6325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1189_0 <=( _mesh_4_5_io_out_valid_0) ^ ((fiEnable && (6326 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1190_0 <=( _mesh_5_5_io_out_valid_0) ^ ((fiEnable && (6327 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1191_0 <=( _mesh_6_5_io_out_valid_0) ^ ((fiEnable && (6328 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1192_0 <=( _mesh_7_5_io_out_valid_0) ^ ((fiEnable && (6329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1193_0 <=( _mesh_8_5_io_out_valid_0) ^ ((fiEnable && (6330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1194_0 <=( _mesh_9_5_io_out_valid_0) ^ ((fiEnable && (6331 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1195_0 <=( _mesh_10_5_io_out_valid_0) ^ ((fiEnable && (6332 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1196_0 <=( _mesh_11_5_io_out_valid_0) ^ ((fiEnable && (6333 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1197_0 <=( _mesh_12_5_io_out_valid_0) ^ ((fiEnable && (6334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1198_0 <=( _mesh_13_5_io_out_valid_0) ^ ((fiEnable && (6335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1199_0 <=( _mesh_14_5_io_out_valid_0) ^ ((fiEnable && (6336 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1200_0 <=( _mesh_15_5_io_out_valid_0) ^ ((fiEnable && (6337 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1201_0 <=( _mesh_16_5_io_out_valid_0) ^ ((fiEnable && (6338 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1202_0 <=( _mesh_17_5_io_out_valid_0) ^ ((fiEnable && (6339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1203_0 <=( _mesh_18_5_io_out_valid_0) ^ ((fiEnable && (6340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1204_0 <=( _mesh_19_5_io_out_valid_0) ^ ((fiEnable && (6341 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1205_0 <=( _mesh_20_5_io_out_valid_0) ^ ((fiEnable && (6342 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1206_0 <=( _mesh_21_5_io_out_valid_0) ^ ((fiEnable && (6343 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1207_0 <=( _mesh_22_5_io_out_valid_0) ^ ((fiEnable && (6344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1208_0 <=( _mesh_23_5_io_out_valid_0) ^ ((fiEnable && (6345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1209_0 <=( _mesh_24_5_io_out_valid_0) ^ ((fiEnable && (6346 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1210_0 <=( _mesh_25_5_io_out_valid_0) ^ ((fiEnable && (6347 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1211_0 <=( _mesh_26_5_io_out_valid_0) ^ ((fiEnable && (6348 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1212_0 <=( _mesh_27_5_io_out_valid_0) ^ ((fiEnable && (6349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1213_0 <=( _mesh_28_5_io_out_valid_0) ^ ((fiEnable && (6350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1214_0 <=( _mesh_29_5_io_out_valid_0) ^ ((fiEnable && (6351 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1215_0 <=( _mesh_30_5_io_out_valid_0) ^ ((fiEnable && (6352 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1216_0 <=( io_in_valid_6_0) ^ ((fiEnable && (6353 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1217_0 <=( _mesh_0_6_io_out_valid_0) ^ ((fiEnable && (6354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1218_0 <=( _mesh_1_6_io_out_valid_0) ^ ((fiEnable && (6355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1219_0 <=( _mesh_2_6_io_out_valid_0) ^ ((fiEnable && (6356 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1220_0 <=( _mesh_3_6_io_out_valid_0) ^ ((fiEnable && (6357 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1221_0 <=( _mesh_4_6_io_out_valid_0) ^ ((fiEnable && (6358 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1222_0 <=( _mesh_5_6_io_out_valid_0) ^ ((fiEnable && (6359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1223_0 <=( _mesh_6_6_io_out_valid_0) ^ ((fiEnable && (6360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1224_0 <=( _mesh_7_6_io_out_valid_0) ^ ((fiEnable && (6361 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1225_0 <=( _mesh_8_6_io_out_valid_0) ^ ((fiEnable && (6362 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1226_0 <=( _mesh_9_6_io_out_valid_0) ^ ((fiEnable && (6363 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1227_0 <=( _mesh_10_6_io_out_valid_0) ^ ((fiEnable && (6364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1228_0 <=( _mesh_11_6_io_out_valid_0) ^ ((fiEnable && (6365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1229_0 <=( _mesh_12_6_io_out_valid_0) ^ ((fiEnable && (6366 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1230_0 <=( _mesh_13_6_io_out_valid_0) ^ ((fiEnable && (6367 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1231_0 <=( _mesh_14_6_io_out_valid_0) ^ ((fiEnable && (6368 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1232_0 <=( _mesh_15_6_io_out_valid_0) ^ ((fiEnable && (6369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1233_0 <=( _mesh_16_6_io_out_valid_0) ^ ((fiEnable && (6370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1234_0 <=( _mesh_17_6_io_out_valid_0) ^ ((fiEnable && (6371 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1235_0 <=( _mesh_18_6_io_out_valid_0) ^ ((fiEnable && (6372 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1236_0 <=( _mesh_19_6_io_out_valid_0) ^ ((fiEnable && (6373 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1237_0 <=( _mesh_20_6_io_out_valid_0) ^ ((fiEnable && (6374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1238_0 <=( _mesh_21_6_io_out_valid_0) ^ ((fiEnable && (6375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1239_0 <=( _mesh_22_6_io_out_valid_0) ^ ((fiEnable && (6376 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1240_0 <=( _mesh_23_6_io_out_valid_0) ^ ((fiEnable && (6377 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1241_0 <=( _mesh_24_6_io_out_valid_0) ^ ((fiEnable && (6378 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1242_0 <=( _mesh_25_6_io_out_valid_0) ^ ((fiEnable && (6379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1243_0 <=( _mesh_26_6_io_out_valid_0) ^ ((fiEnable && (6380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1244_0 <=( _mesh_27_6_io_out_valid_0) ^ ((fiEnable && (6381 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1245_0 <=( _mesh_28_6_io_out_valid_0) ^ ((fiEnable && (6382 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1246_0 <=( _mesh_29_6_io_out_valid_0) ^ ((fiEnable && (6383 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1247_0 <=( _mesh_30_6_io_out_valid_0) ^ ((fiEnable && (6384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1248_0 <=( io_in_valid_7_0) ^ ((fiEnable && (6385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1249_0 <=( _mesh_0_7_io_out_valid_0) ^ ((fiEnable && (6386 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1250_0 <=( _mesh_1_7_io_out_valid_0) ^ ((fiEnable && (6387 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1251_0 <=( _mesh_2_7_io_out_valid_0) ^ ((fiEnable && (6388 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1252_0 <=( _mesh_3_7_io_out_valid_0) ^ ((fiEnable && (6389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1253_0 <=( _mesh_4_7_io_out_valid_0) ^ ((fiEnable && (6390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1254_0 <=( _mesh_5_7_io_out_valid_0) ^ ((fiEnable && (6391 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1255_0 <=( _mesh_6_7_io_out_valid_0) ^ ((fiEnable && (6392 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1256_0 <=( _mesh_7_7_io_out_valid_0) ^ ((fiEnable && (6393 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1257_0 <=( _mesh_8_7_io_out_valid_0) ^ ((fiEnable && (6394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1258_0 <=( _mesh_9_7_io_out_valid_0) ^ ((fiEnable && (6395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1259_0 <=( _mesh_10_7_io_out_valid_0) ^ ((fiEnable && (6396 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1260_0 <=( _mesh_11_7_io_out_valid_0) ^ ((fiEnable && (6397 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1261_0 <=( _mesh_12_7_io_out_valid_0) ^ ((fiEnable && (6398 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1262_0 <=( _mesh_13_7_io_out_valid_0) ^ ((fiEnable && (6399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1263_0 <=( _mesh_14_7_io_out_valid_0) ^ ((fiEnable && (6400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1264_0 <=( _mesh_15_7_io_out_valid_0) ^ ((fiEnable && (6401 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1265_0 <=( _mesh_16_7_io_out_valid_0) ^ ((fiEnable && (6402 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1266_0 <=( _mesh_17_7_io_out_valid_0) ^ ((fiEnable && (6403 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1267_0 <=( _mesh_18_7_io_out_valid_0) ^ ((fiEnable && (6404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1268_0 <=( _mesh_19_7_io_out_valid_0) ^ ((fiEnable && (6405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1269_0 <=( _mesh_20_7_io_out_valid_0) ^ ((fiEnable && (6406 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1270_0 <=( _mesh_21_7_io_out_valid_0) ^ ((fiEnable && (6407 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1271_0 <=( _mesh_22_7_io_out_valid_0) ^ ((fiEnable && (6408 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1272_0 <=( _mesh_23_7_io_out_valid_0) ^ ((fiEnable && (6409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1273_0 <=( _mesh_24_7_io_out_valid_0) ^ ((fiEnable && (6410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1274_0 <=( _mesh_25_7_io_out_valid_0) ^ ((fiEnable && (6411 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1275_0 <=( _mesh_26_7_io_out_valid_0) ^ ((fiEnable && (6412 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1276_0 <=( _mesh_27_7_io_out_valid_0) ^ ((fiEnable && (6413 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1277_0 <=( _mesh_28_7_io_out_valid_0) ^ ((fiEnable && (6414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1278_0 <=( _mesh_29_7_io_out_valid_0) ^ ((fiEnable && (6415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1279_0 <=( _mesh_30_7_io_out_valid_0) ^ ((fiEnable && (6416 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1280_0 <=( io_in_valid_8_0) ^ ((fiEnable && (6417 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1281_0 <=( _mesh_0_8_io_out_valid_0) ^ ((fiEnable && (6418 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1282_0 <=( _mesh_1_8_io_out_valid_0) ^ ((fiEnable && (6419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1283_0 <=( _mesh_2_8_io_out_valid_0) ^ ((fiEnable && (6420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1284_0 <=( _mesh_3_8_io_out_valid_0) ^ ((fiEnable && (6421 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1285_0 <=( _mesh_4_8_io_out_valid_0) ^ ((fiEnable && (6422 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1286_0 <=( _mesh_5_8_io_out_valid_0) ^ ((fiEnable && (6423 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1287_0 <=( _mesh_6_8_io_out_valid_0) ^ ((fiEnable && (6424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1288_0 <=( _mesh_7_8_io_out_valid_0) ^ ((fiEnable && (6425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1289_0 <=( _mesh_8_8_io_out_valid_0) ^ ((fiEnable && (6426 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1290_0 <=( _mesh_9_8_io_out_valid_0) ^ ((fiEnable && (6427 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1291_0 <=( _mesh_10_8_io_out_valid_0) ^ ((fiEnable && (6428 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1292_0 <=( _mesh_11_8_io_out_valid_0) ^ ((fiEnable && (6429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1293_0 <=( _mesh_12_8_io_out_valid_0) ^ ((fiEnable && (6430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1294_0 <=( _mesh_13_8_io_out_valid_0) ^ ((fiEnable && (6431 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1295_0 <=( _mesh_14_8_io_out_valid_0) ^ ((fiEnable && (6432 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1296_0 <=( _mesh_15_8_io_out_valid_0) ^ ((fiEnable && (6433 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1297_0 <=( _mesh_16_8_io_out_valid_0) ^ ((fiEnable && (6434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1298_0 <=( _mesh_17_8_io_out_valid_0) ^ ((fiEnable && (6435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1299_0 <=( _mesh_18_8_io_out_valid_0) ^ ((fiEnable && (6436 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1300_0 <=( _mesh_19_8_io_out_valid_0) ^ ((fiEnable && (6437 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1301_0 <=( _mesh_20_8_io_out_valid_0) ^ ((fiEnable && (6438 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1302_0 <=( _mesh_21_8_io_out_valid_0) ^ ((fiEnable && (6439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1303_0 <=( _mesh_22_8_io_out_valid_0) ^ ((fiEnable && (6440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1304_0 <=( _mesh_23_8_io_out_valid_0) ^ ((fiEnable && (6441 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1305_0 <=( _mesh_24_8_io_out_valid_0) ^ ((fiEnable && (6442 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1306_0 <=( _mesh_25_8_io_out_valid_0) ^ ((fiEnable && (6443 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1307_0 <=( _mesh_26_8_io_out_valid_0) ^ ((fiEnable && (6444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1308_0 <=( _mesh_27_8_io_out_valid_0) ^ ((fiEnable && (6445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1309_0 <=( _mesh_28_8_io_out_valid_0) ^ ((fiEnable && (6446 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1310_0 <=( _mesh_29_8_io_out_valid_0) ^ ((fiEnable && (6447 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1311_0 <=( _mesh_30_8_io_out_valid_0) ^ ((fiEnable && (6448 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1312_0 <=( io_in_valid_9_0) ^ ((fiEnable && (6449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1313_0 <=( _mesh_0_9_io_out_valid_0) ^ ((fiEnable && (6450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1314_0 <=( _mesh_1_9_io_out_valid_0) ^ ((fiEnable && (6451 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1315_0 <=( _mesh_2_9_io_out_valid_0) ^ ((fiEnable && (6452 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1316_0 <=( _mesh_3_9_io_out_valid_0) ^ ((fiEnable && (6453 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1317_0 <=( _mesh_4_9_io_out_valid_0) ^ ((fiEnable && (6454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1318_0 <=( _mesh_5_9_io_out_valid_0) ^ ((fiEnable && (6455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1319_0 <=( _mesh_6_9_io_out_valid_0) ^ ((fiEnable && (6456 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1320_0 <=( _mesh_7_9_io_out_valid_0) ^ ((fiEnable && (6457 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1321_0 <=( _mesh_8_9_io_out_valid_0) ^ ((fiEnable && (6458 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1322_0 <=( _mesh_9_9_io_out_valid_0) ^ ((fiEnable && (6459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1323_0 <=( _mesh_10_9_io_out_valid_0) ^ ((fiEnable && (6460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1324_0 <=( _mesh_11_9_io_out_valid_0) ^ ((fiEnable && (6461 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1325_0 <=( _mesh_12_9_io_out_valid_0) ^ ((fiEnable && (6462 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1326_0 <=( _mesh_13_9_io_out_valid_0) ^ ((fiEnable && (6463 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1327_0 <=( _mesh_14_9_io_out_valid_0) ^ ((fiEnable && (6464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1328_0 <=( _mesh_15_9_io_out_valid_0) ^ ((fiEnable && (6465 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1329_0 <=( _mesh_16_9_io_out_valid_0) ^ ((fiEnable && (6466 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1330_0 <=( _mesh_17_9_io_out_valid_0) ^ ((fiEnable && (6467 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1331_0 <=( _mesh_18_9_io_out_valid_0) ^ ((fiEnable && (6468 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1332_0 <=( _mesh_19_9_io_out_valid_0) ^ ((fiEnable && (6469 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1333_0 <=( _mesh_20_9_io_out_valid_0) ^ ((fiEnable && (6470 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1334_0 <=( _mesh_21_9_io_out_valid_0) ^ ((fiEnable && (6471 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1335_0 <=( _mesh_22_9_io_out_valid_0) ^ ((fiEnable && (6472 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1336_0 <=( _mesh_23_9_io_out_valid_0) ^ ((fiEnable && (6473 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1337_0 <=( _mesh_24_9_io_out_valid_0) ^ ((fiEnable && (6474 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1338_0 <=( _mesh_25_9_io_out_valid_0) ^ ((fiEnable && (6475 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1339_0 <=( _mesh_26_9_io_out_valid_0) ^ ((fiEnable && (6476 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1340_0 <=( _mesh_27_9_io_out_valid_0) ^ ((fiEnable && (6477 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1341_0 <=( _mesh_28_9_io_out_valid_0) ^ ((fiEnable && (6478 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1342_0 <=( _mesh_29_9_io_out_valid_0) ^ ((fiEnable && (6479 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1343_0 <=( _mesh_30_9_io_out_valid_0) ^ ((fiEnable && (6480 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1344_0 <=( io_in_valid_10_0) ^ ((fiEnable && (6481 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1345_0 <=( _mesh_0_10_io_out_valid_0) ^ ((fiEnable && (6482 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1346_0 <=( _mesh_1_10_io_out_valid_0) ^ ((fiEnable && (6483 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1347_0 <=( _mesh_2_10_io_out_valid_0) ^ ((fiEnable && (6484 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1348_0 <=( _mesh_3_10_io_out_valid_0) ^ ((fiEnable && (6485 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1349_0 <=( _mesh_4_10_io_out_valid_0) ^ ((fiEnable && (6486 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1350_0 <=( _mesh_5_10_io_out_valid_0) ^ ((fiEnable && (6487 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1351_0 <=( _mesh_6_10_io_out_valid_0) ^ ((fiEnable && (6488 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1352_0 <=( _mesh_7_10_io_out_valid_0) ^ ((fiEnable && (6489 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1353_0 <=( _mesh_8_10_io_out_valid_0) ^ ((fiEnable && (6490 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1354_0 <=( _mesh_9_10_io_out_valid_0) ^ ((fiEnable && (6491 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1355_0 <=( _mesh_10_10_io_out_valid_0) ^ ((fiEnable && (6492 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1356_0 <=( _mesh_11_10_io_out_valid_0) ^ ((fiEnable && (6493 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1357_0 <=( _mesh_12_10_io_out_valid_0) ^ ((fiEnable && (6494 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1358_0 <=( _mesh_13_10_io_out_valid_0) ^ ((fiEnable && (6495 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1359_0 <=( _mesh_14_10_io_out_valid_0) ^ ((fiEnable && (6496 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1360_0 <=( _mesh_15_10_io_out_valid_0) ^ ((fiEnable && (6497 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1361_0 <=( _mesh_16_10_io_out_valid_0) ^ ((fiEnable && (6498 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1362_0 <=( _mesh_17_10_io_out_valid_0) ^ ((fiEnable && (6499 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1363_0 <=( _mesh_18_10_io_out_valid_0) ^ ((fiEnable && (6500 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1364_0 <=( _mesh_19_10_io_out_valid_0) ^ ((fiEnable && (6501 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1365_0 <=( _mesh_20_10_io_out_valid_0) ^ ((fiEnable && (6502 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1366_0 <=( _mesh_21_10_io_out_valid_0) ^ ((fiEnable && (6503 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1367_0 <=( _mesh_22_10_io_out_valid_0) ^ ((fiEnable && (6504 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1368_0 <=( _mesh_23_10_io_out_valid_0) ^ ((fiEnable && (6505 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1369_0 <=( _mesh_24_10_io_out_valid_0) ^ ((fiEnable && (6506 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1370_0 <=( _mesh_25_10_io_out_valid_0) ^ ((fiEnable && (6507 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1371_0 <=( _mesh_26_10_io_out_valid_0) ^ ((fiEnable && (6508 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1372_0 <=( _mesh_27_10_io_out_valid_0) ^ ((fiEnable && (6509 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1373_0 <=( _mesh_28_10_io_out_valid_0) ^ ((fiEnable && (6510 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1374_0 <=( _mesh_29_10_io_out_valid_0) ^ ((fiEnable && (6511 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1375_0 <=( _mesh_30_10_io_out_valid_0) ^ ((fiEnable && (6512 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1376_0 <=( io_in_valid_11_0) ^ ((fiEnable && (6513 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1377_0 <=( _mesh_0_11_io_out_valid_0) ^ ((fiEnable && (6514 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1378_0 <=( _mesh_1_11_io_out_valid_0) ^ ((fiEnable && (6515 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1379_0 <=( _mesh_2_11_io_out_valid_0) ^ ((fiEnable && (6516 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1380_0 <=( _mesh_3_11_io_out_valid_0) ^ ((fiEnable && (6517 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1381_0 <=( _mesh_4_11_io_out_valid_0) ^ ((fiEnable && (6518 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1382_0 <=( _mesh_5_11_io_out_valid_0) ^ ((fiEnable && (6519 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1383_0 <=( _mesh_6_11_io_out_valid_0) ^ ((fiEnable && (6520 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1384_0 <=( _mesh_7_11_io_out_valid_0) ^ ((fiEnable && (6521 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1385_0 <=( _mesh_8_11_io_out_valid_0) ^ ((fiEnable && (6522 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1386_0 <=( _mesh_9_11_io_out_valid_0) ^ ((fiEnable && (6523 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1387_0 <=( _mesh_10_11_io_out_valid_0) ^ ((fiEnable && (6524 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1388_0 <=( _mesh_11_11_io_out_valid_0) ^ ((fiEnable && (6525 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1389_0 <=( _mesh_12_11_io_out_valid_0) ^ ((fiEnable && (6526 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1390_0 <=( _mesh_13_11_io_out_valid_0) ^ ((fiEnable && (6527 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1391_0 <=( _mesh_14_11_io_out_valid_0) ^ ((fiEnable && (6528 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1392_0 <=( _mesh_15_11_io_out_valid_0) ^ ((fiEnable && (6529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1393_0 <=( _mesh_16_11_io_out_valid_0) ^ ((fiEnable && (6530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1394_0 <=( _mesh_17_11_io_out_valid_0) ^ ((fiEnable && (6531 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1395_0 <=( _mesh_18_11_io_out_valid_0) ^ ((fiEnable && (6532 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1396_0 <=( _mesh_19_11_io_out_valid_0) ^ ((fiEnable && (6533 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1397_0 <=( _mesh_20_11_io_out_valid_0) ^ ((fiEnable && (6534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1398_0 <=( _mesh_21_11_io_out_valid_0) ^ ((fiEnable && (6535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1399_0 <=( _mesh_22_11_io_out_valid_0) ^ ((fiEnable && (6536 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1400_0 <=( _mesh_23_11_io_out_valid_0) ^ ((fiEnable && (6537 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1401_0 <=( _mesh_24_11_io_out_valid_0) ^ ((fiEnable && (6538 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1402_0 <=( _mesh_25_11_io_out_valid_0) ^ ((fiEnable && (6539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1403_0 <=( _mesh_26_11_io_out_valid_0) ^ ((fiEnable && (6540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1404_0 <=( _mesh_27_11_io_out_valid_0) ^ ((fiEnable && (6541 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1405_0 <=( _mesh_28_11_io_out_valid_0) ^ ((fiEnable && (6542 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1406_0 <=( _mesh_29_11_io_out_valid_0) ^ ((fiEnable && (6543 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1407_0 <=( _mesh_30_11_io_out_valid_0) ^ ((fiEnable && (6544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1408_0 <=( io_in_valid_12_0) ^ ((fiEnable && (6545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1409_0 <=( _mesh_0_12_io_out_valid_0) ^ ((fiEnable && (6546 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1410_0 <=( _mesh_1_12_io_out_valid_0) ^ ((fiEnable && (6547 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1411_0 <=( _mesh_2_12_io_out_valid_0) ^ ((fiEnable && (6548 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1412_0 <=( _mesh_3_12_io_out_valid_0) ^ ((fiEnable && (6549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1413_0 <=( _mesh_4_12_io_out_valid_0) ^ ((fiEnable && (6550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1414_0 <=( _mesh_5_12_io_out_valid_0) ^ ((fiEnable && (6551 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1415_0 <=( _mesh_6_12_io_out_valid_0) ^ ((fiEnable && (6552 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1416_0 <=( _mesh_7_12_io_out_valid_0) ^ ((fiEnable && (6553 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1417_0 <=( _mesh_8_12_io_out_valid_0) ^ ((fiEnable && (6554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1418_0 <=( _mesh_9_12_io_out_valid_0) ^ ((fiEnable && (6555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1419_0 <=( _mesh_10_12_io_out_valid_0) ^ ((fiEnable && (6556 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1420_0 <=( _mesh_11_12_io_out_valid_0) ^ ((fiEnable && (6557 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1421_0 <=( _mesh_12_12_io_out_valid_0) ^ ((fiEnable && (6558 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1422_0 <=( _mesh_13_12_io_out_valid_0) ^ ((fiEnable && (6559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1423_0 <=( _mesh_14_12_io_out_valid_0) ^ ((fiEnable && (6560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1424_0 <=( _mesh_15_12_io_out_valid_0) ^ ((fiEnable && (6561 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1425_0 <=( _mesh_16_12_io_out_valid_0) ^ ((fiEnable && (6562 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1426_0 <=( _mesh_17_12_io_out_valid_0) ^ ((fiEnable && (6563 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1427_0 <=( _mesh_18_12_io_out_valid_0) ^ ((fiEnable && (6564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1428_0 <=( _mesh_19_12_io_out_valid_0) ^ ((fiEnable && (6565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1429_0 <=( _mesh_20_12_io_out_valid_0) ^ ((fiEnable && (6566 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1430_0 <=( _mesh_21_12_io_out_valid_0) ^ ((fiEnable && (6567 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1431_0 <=( _mesh_22_12_io_out_valid_0) ^ ((fiEnable && (6568 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1432_0 <=( _mesh_23_12_io_out_valid_0) ^ ((fiEnable && (6569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1433_0 <=( _mesh_24_12_io_out_valid_0) ^ ((fiEnable && (6570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1434_0 <=( _mesh_25_12_io_out_valid_0) ^ ((fiEnable && (6571 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1435_0 <=( _mesh_26_12_io_out_valid_0) ^ ((fiEnable && (6572 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1436_0 <=( _mesh_27_12_io_out_valid_0) ^ ((fiEnable && (6573 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1437_0 <=( _mesh_28_12_io_out_valid_0) ^ ((fiEnable && (6574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1438_0 <=( _mesh_29_12_io_out_valid_0) ^ ((fiEnable && (6575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1439_0 <=( _mesh_30_12_io_out_valid_0) ^ ((fiEnable && (6576 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1440_0 <=( io_in_valid_13_0) ^ ((fiEnable && (6577 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1441_0 <=( _mesh_0_13_io_out_valid_0) ^ ((fiEnable && (6578 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1442_0 <=( _mesh_1_13_io_out_valid_0) ^ ((fiEnable && (6579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1443_0 <=( _mesh_2_13_io_out_valid_0) ^ ((fiEnable && (6580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1444_0 <=( _mesh_3_13_io_out_valid_0) ^ ((fiEnable && (6581 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1445_0 <=( _mesh_4_13_io_out_valid_0) ^ ((fiEnable && (6582 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1446_0 <=( _mesh_5_13_io_out_valid_0) ^ ((fiEnable && (6583 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1447_0 <=( _mesh_6_13_io_out_valid_0) ^ ((fiEnable && (6584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1448_0 <=( _mesh_7_13_io_out_valid_0) ^ ((fiEnable && (6585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1449_0 <=( _mesh_8_13_io_out_valid_0) ^ ((fiEnable && (6586 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1450_0 <=( _mesh_9_13_io_out_valid_0) ^ ((fiEnable && (6587 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1451_0 <=( _mesh_10_13_io_out_valid_0) ^ ((fiEnable && (6588 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1452_0 <=( _mesh_11_13_io_out_valid_0) ^ ((fiEnable && (6589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1453_0 <=( _mesh_12_13_io_out_valid_0) ^ ((fiEnable && (6590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1454_0 <=( _mesh_13_13_io_out_valid_0) ^ ((fiEnable && (6591 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1455_0 <=( _mesh_14_13_io_out_valid_0) ^ ((fiEnable && (6592 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1456_0 <=( _mesh_15_13_io_out_valid_0) ^ ((fiEnable && (6593 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1457_0 <=( _mesh_16_13_io_out_valid_0) ^ ((fiEnable && (6594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1458_0 <=( _mesh_17_13_io_out_valid_0) ^ ((fiEnable && (6595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1459_0 <=( _mesh_18_13_io_out_valid_0) ^ ((fiEnable && (6596 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1460_0 <=( _mesh_19_13_io_out_valid_0) ^ ((fiEnable && (6597 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1461_0 <=( _mesh_20_13_io_out_valid_0) ^ ((fiEnable && (6598 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1462_0 <=( _mesh_21_13_io_out_valid_0) ^ ((fiEnable && (6599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1463_0 <=( _mesh_22_13_io_out_valid_0) ^ ((fiEnable && (6600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1464_0 <=( _mesh_23_13_io_out_valid_0) ^ ((fiEnable && (6601 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1465_0 <=( _mesh_24_13_io_out_valid_0) ^ ((fiEnable && (6602 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1466_0 <=( _mesh_25_13_io_out_valid_0) ^ ((fiEnable && (6603 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1467_0 <=( _mesh_26_13_io_out_valid_0) ^ ((fiEnable && (6604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1468_0 <=( _mesh_27_13_io_out_valid_0) ^ ((fiEnable && (6605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1469_0 <=( _mesh_28_13_io_out_valid_0) ^ ((fiEnable && (6606 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1470_0 <=( _mesh_29_13_io_out_valid_0) ^ ((fiEnable && (6607 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1471_0 <=( _mesh_30_13_io_out_valid_0) ^ ((fiEnable && (6608 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1472_0 <=( io_in_valid_14_0) ^ ((fiEnable && (6609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1473_0 <=( _mesh_0_14_io_out_valid_0) ^ ((fiEnable && (6610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1474_0 <=( _mesh_1_14_io_out_valid_0) ^ ((fiEnable && (6611 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1475_0 <=( _mesh_2_14_io_out_valid_0) ^ ((fiEnable && (6612 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1476_0 <=( _mesh_3_14_io_out_valid_0) ^ ((fiEnable && (6613 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1477_0 <=( _mesh_4_14_io_out_valid_0) ^ ((fiEnable && (6614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1478_0 <=( _mesh_5_14_io_out_valid_0) ^ ((fiEnable && (6615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1479_0 <=( _mesh_6_14_io_out_valid_0) ^ ((fiEnable && (6616 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1480_0 <=( _mesh_7_14_io_out_valid_0) ^ ((fiEnable && (6617 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1481_0 <=( _mesh_8_14_io_out_valid_0) ^ ((fiEnable && (6618 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1482_0 <=( _mesh_9_14_io_out_valid_0) ^ ((fiEnable && (6619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1483_0 <=( _mesh_10_14_io_out_valid_0) ^ ((fiEnable && (6620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1484_0 <=( _mesh_11_14_io_out_valid_0) ^ ((fiEnable && (6621 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1485_0 <=( _mesh_12_14_io_out_valid_0) ^ ((fiEnable && (6622 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1486_0 <=( _mesh_13_14_io_out_valid_0) ^ ((fiEnable && (6623 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1487_0 <=( _mesh_14_14_io_out_valid_0) ^ ((fiEnable && (6624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1488_0 <=( _mesh_15_14_io_out_valid_0) ^ ((fiEnable && (6625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1489_0 <=( _mesh_16_14_io_out_valid_0) ^ ((fiEnable && (6626 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1490_0 <=( _mesh_17_14_io_out_valid_0) ^ ((fiEnable && (6627 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1491_0 <=( _mesh_18_14_io_out_valid_0) ^ ((fiEnable && (6628 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1492_0 <=( _mesh_19_14_io_out_valid_0) ^ ((fiEnable && (6629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1493_0 <=( _mesh_20_14_io_out_valid_0) ^ ((fiEnable && (6630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1494_0 <=( _mesh_21_14_io_out_valid_0) ^ ((fiEnable && (6631 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1495_0 <=( _mesh_22_14_io_out_valid_0) ^ ((fiEnable && (6632 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1496_0 <=( _mesh_23_14_io_out_valid_0) ^ ((fiEnable && (6633 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1497_0 <=( _mesh_24_14_io_out_valid_0) ^ ((fiEnable && (6634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1498_0 <=( _mesh_25_14_io_out_valid_0) ^ ((fiEnable && (6635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1499_0 <=( _mesh_26_14_io_out_valid_0) ^ ((fiEnable && (6636 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1500_0 <=( _mesh_27_14_io_out_valid_0) ^ ((fiEnable && (6637 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1501_0 <=( _mesh_28_14_io_out_valid_0) ^ ((fiEnable && (6638 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1502_0 <=( _mesh_29_14_io_out_valid_0) ^ ((fiEnable && (6639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1503_0 <=( _mesh_30_14_io_out_valid_0) ^ ((fiEnable && (6640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1504_0 <=( io_in_valid_15_0) ^ ((fiEnable && (6641 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1505_0 <=( _mesh_0_15_io_out_valid_0) ^ ((fiEnable && (6642 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1506_0 <=( _mesh_1_15_io_out_valid_0) ^ ((fiEnable && (6643 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1507_0 <=( _mesh_2_15_io_out_valid_0) ^ ((fiEnable && (6644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1508_0 <=( _mesh_3_15_io_out_valid_0) ^ ((fiEnable && (6645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1509_0 <=( _mesh_4_15_io_out_valid_0) ^ ((fiEnable && (6646 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1510_0 <=( _mesh_5_15_io_out_valid_0) ^ ((fiEnable && (6647 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1511_0 <=( _mesh_6_15_io_out_valid_0) ^ ((fiEnable && (6648 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1512_0 <=( _mesh_7_15_io_out_valid_0) ^ ((fiEnable && (6649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1513_0 <=( _mesh_8_15_io_out_valid_0) ^ ((fiEnable && (6650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1514_0 <=( _mesh_9_15_io_out_valid_0) ^ ((fiEnable && (6651 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1515_0 <=( _mesh_10_15_io_out_valid_0) ^ ((fiEnable && (6652 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1516_0 <=( _mesh_11_15_io_out_valid_0) ^ ((fiEnable && (6653 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1517_0 <=( _mesh_12_15_io_out_valid_0) ^ ((fiEnable && (6654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1518_0 <=( _mesh_13_15_io_out_valid_0) ^ ((fiEnable && (6655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1519_0 <=( _mesh_14_15_io_out_valid_0) ^ ((fiEnable && (6656 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1520_0 <=( _mesh_15_15_io_out_valid_0) ^ ((fiEnable && (6657 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1521_0 <=( _mesh_16_15_io_out_valid_0) ^ ((fiEnable && (6658 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1522_0 <=( _mesh_17_15_io_out_valid_0) ^ ((fiEnable && (6659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1523_0 <=( _mesh_18_15_io_out_valid_0) ^ ((fiEnable && (6660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1524_0 <=( _mesh_19_15_io_out_valid_0) ^ ((fiEnable && (6661 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1525_0 <=( _mesh_20_15_io_out_valid_0) ^ ((fiEnable && (6662 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1526_0 <=( _mesh_21_15_io_out_valid_0) ^ ((fiEnable && (6663 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1527_0 <=( _mesh_22_15_io_out_valid_0) ^ ((fiEnable && (6664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1528_0 <=( _mesh_23_15_io_out_valid_0) ^ ((fiEnable && (6665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1529_0 <=( _mesh_24_15_io_out_valid_0) ^ ((fiEnable && (6666 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1530_0 <=( _mesh_25_15_io_out_valid_0) ^ ((fiEnable && (6667 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1531_0 <=( _mesh_26_15_io_out_valid_0) ^ ((fiEnable && (6668 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1532_0 <=( _mesh_27_15_io_out_valid_0) ^ ((fiEnable && (6669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1533_0 <=( _mesh_28_15_io_out_valid_0) ^ ((fiEnable && (6670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1534_0 <=( _mesh_29_15_io_out_valid_0) ^ ((fiEnable && (6671 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1535_0 <=( _mesh_30_15_io_out_valid_0) ^ ((fiEnable && (6672 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1536_0 <=( io_in_valid_16_0) ^ ((fiEnable && (6673 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1537_0 <=( _mesh_0_16_io_out_valid_0) ^ ((fiEnable && (6674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1538_0 <=( _mesh_1_16_io_out_valid_0) ^ ((fiEnable && (6675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1539_0 <=( _mesh_2_16_io_out_valid_0) ^ ((fiEnable && (6676 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1540_0 <=( _mesh_3_16_io_out_valid_0) ^ ((fiEnable && (6677 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1541_0 <=( _mesh_4_16_io_out_valid_0) ^ ((fiEnable && (6678 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1542_0 <=( _mesh_5_16_io_out_valid_0) ^ ((fiEnable && (6679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1543_0 <=( _mesh_6_16_io_out_valid_0) ^ ((fiEnable && (6680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1544_0 <=( _mesh_7_16_io_out_valid_0) ^ ((fiEnable && (6681 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1545_0 <=( _mesh_8_16_io_out_valid_0) ^ ((fiEnable && (6682 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1546_0 <=( _mesh_9_16_io_out_valid_0) ^ ((fiEnable && (6683 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1547_0 <=( _mesh_10_16_io_out_valid_0) ^ ((fiEnable && (6684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1548_0 <=( _mesh_11_16_io_out_valid_0) ^ ((fiEnable && (6685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1549_0 <=( _mesh_12_16_io_out_valid_0) ^ ((fiEnable && (6686 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1550_0 <=( _mesh_13_16_io_out_valid_0) ^ ((fiEnable && (6687 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1551_0 <=( _mesh_14_16_io_out_valid_0) ^ ((fiEnable && (6688 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1552_0 <=( _mesh_15_16_io_out_valid_0) ^ ((fiEnable && (6689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1553_0 <=( _mesh_16_16_io_out_valid_0) ^ ((fiEnable && (6690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1554_0 <=( _mesh_17_16_io_out_valid_0) ^ ((fiEnable && (6691 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1555_0 <=( _mesh_18_16_io_out_valid_0) ^ ((fiEnable && (6692 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1556_0 <=( _mesh_19_16_io_out_valid_0) ^ ((fiEnable && (6693 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1557_0 <=( _mesh_20_16_io_out_valid_0) ^ ((fiEnable && (6694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1558_0 <=( _mesh_21_16_io_out_valid_0) ^ ((fiEnable && (6695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1559_0 <=( _mesh_22_16_io_out_valid_0) ^ ((fiEnable && (6696 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1560_0 <=( _mesh_23_16_io_out_valid_0) ^ ((fiEnable && (6697 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1561_0 <=( _mesh_24_16_io_out_valid_0) ^ ((fiEnable && (6698 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1562_0 <=( _mesh_25_16_io_out_valid_0) ^ ((fiEnable && (6699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1563_0 <=( _mesh_26_16_io_out_valid_0) ^ ((fiEnable && (6700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1564_0 <=( _mesh_27_16_io_out_valid_0) ^ ((fiEnable && (6701 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1565_0 <=( _mesh_28_16_io_out_valid_0) ^ ((fiEnable && (6702 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1566_0 <=( _mesh_29_16_io_out_valid_0) ^ ((fiEnable && (6703 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1567_0 <=( _mesh_30_16_io_out_valid_0) ^ ((fiEnable && (6704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1568_0 <=( io_in_valid_17_0) ^ ((fiEnable && (6705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1569_0 <=( _mesh_0_17_io_out_valid_0) ^ ((fiEnable && (6706 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1570_0 <=( _mesh_1_17_io_out_valid_0) ^ ((fiEnable && (6707 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1571_0 <=( _mesh_2_17_io_out_valid_0) ^ ((fiEnable && (6708 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1572_0 <=( _mesh_3_17_io_out_valid_0) ^ ((fiEnable && (6709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1573_0 <=( _mesh_4_17_io_out_valid_0) ^ ((fiEnable && (6710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1574_0 <=( _mesh_5_17_io_out_valid_0) ^ ((fiEnable && (6711 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1575_0 <=( _mesh_6_17_io_out_valid_0) ^ ((fiEnable && (6712 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1576_0 <=( _mesh_7_17_io_out_valid_0) ^ ((fiEnable && (6713 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1577_0 <=( _mesh_8_17_io_out_valid_0) ^ ((fiEnable && (6714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1578_0 <=( _mesh_9_17_io_out_valid_0) ^ ((fiEnable && (6715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1579_0 <=( _mesh_10_17_io_out_valid_0) ^ ((fiEnable && (6716 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1580_0 <=( _mesh_11_17_io_out_valid_0) ^ ((fiEnable && (6717 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1581_0 <=( _mesh_12_17_io_out_valid_0) ^ ((fiEnable && (6718 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1582_0 <=( _mesh_13_17_io_out_valid_0) ^ ((fiEnable && (6719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1583_0 <=( _mesh_14_17_io_out_valid_0) ^ ((fiEnable && (6720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1584_0 <=( _mesh_15_17_io_out_valid_0) ^ ((fiEnable && (6721 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1585_0 <=( _mesh_16_17_io_out_valid_0) ^ ((fiEnable && (6722 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1586_0 <=( _mesh_17_17_io_out_valid_0) ^ ((fiEnable && (6723 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1587_0 <=( _mesh_18_17_io_out_valid_0) ^ ((fiEnable && (6724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1588_0 <=( _mesh_19_17_io_out_valid_0) ^ ((fiEnable && (6725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1589_0 <=( _mesh_20_17_io_out_valid_0) ^ ((fiEnable && (6726 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1590_0 <=( _mesh_21_17_io_out_valid_0) ^ ((fiEnable && (6727 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1591_0 <=( _mesh_22_17_io_out_valid_0) ^ ((fiEnable && (6728 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1592_0 <=( _mesh_23_17_io_out_valid_0) ^ ((fiEnable && (6729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1593_0 <=( _mesh_24_17_io_out_valid_0) ^ ((fiEnable && (6730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1594_0 <=( _mesh_25_17_io_out_valid_0) ^ ((fiEnable && (6731 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1595_0 <=( _mesh_26_17_io_out_valid_0) ^ ((fiEnable && (6732 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1596_0 <=( _mesh_27_17_io_out_valid_0) ^ ((fiEnable && (6733 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1597_0 <=( _mesh_28_17_io_out_valid_0) ^ ((fiEnable && (6734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1598_0 <=( _mesh_29_17_io_out_valid_0) ^ ((fiEnable && (6735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1599_0 <=( _mesh_30_17_io_out_valid_0) ^ ((fiEnable && (6736 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1600_0 <=( io_in_valid_18_0) ^ ((fiEnable && (6737 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1601_0 <=( _mesh_0_18_io_out_valid_0) ^ ((fiEnable && (6738 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1602_0 <=( _mesh_1_18_io_out_valid_0) ^ ((fiEnable && (6739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1603_0 <=( _mesh_2_18_io_out_valid_0) ^ ((fiEnable && (6740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1604_0 <=( _mesh_3_18_io_out_valid_0) ^ ((fiEnable && (6741 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1605_0 <=( _mesh_4_18_io_out_valid_0) ^ ((fiEnable && (6742 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1606_0 <=( _mesh_5_18_io_out_valid_0) ^ ((fiEnable && (6743 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1607_0 <=( _mesh_6_18_io_out_valid_0) ^ ((fiEnable && (6744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1608_0 <=( _mesh_7_18_io_out_valid_0) ^ ((fiEnable && (6745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1609_0 <=( _mesh_8_18_io_out_valid_0) ^ ((fiEnable && (6746 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1610_0 <=( _mesh_9_18_io_out_valid_0) ^ ((fiEnable && (6747 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1611_0 <=( _mesh_10_18_io_out_valid_0) ^ ((fiEnable && (6748 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1612_0 <=( _mesh_11_18_io_out_valid_0) ^ ((fiEnable && (6749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1613_0 <=( _mesh_12_18_io_out_valid_0) ^ ((fiEnable && (6750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1614_0 <=( _mesh_13_18_io_out_valid_0) ^ ((fiEnable && (6751 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1615_0 <=( _mesh_14_18_io_out_valid_0) ^ ((fiEnable && (6752 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1616_0 <=( _mesh_15_18_io_out_valid_0) ^ ((fiEnable && (6753 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1617_0 <=( _mesh_16_18_io_out_valid_0) ^ ((fiEnable && (6754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1618_0 <=( _mesh_17_18_io_out_valid_0) ^ ((fiEnable && (6755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1619_0 <=( _mesh_18_18_io_out_valid_0) ^ ((fiEnable && (6756 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1620_0 <=( _mesh_19_18_io_out_valid_0) ^ ((fiEnable && (6757 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1621_0 <=( _mesh_20_18_io_out_valid_0) ^ ((fiEnable && (6758 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1622_0 <=( _mesh_21_18_io_out_valid_0) ^ ((fiEnable && (6759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1623_0 <=( _mesh_22_18_io_out_valid_0) ^ ((fiEnable && (6760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1624_0 <=( _mesh_23_18_io_out_valid_0) ^ ((fiEnable && (6761 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1625_0 <=( _mesh_24_18_io_out_valid_0) ^ ((fiEnable && (6762 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1626_0 <=( _mesh_25_18_io_out_valid_0) ^ ((fiEnable && (6763 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1627_0 <=( _mesh_26_18_io_out_valid_0) ^ ((fiEnable && (6764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1628_0 <=( _mesh_27_18_io_out_valid_0) ^ ((fiEnable && (6765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1629_0 <=( _mesh_28_18_io_out_valid_0) ^ ((fiEnable && (6766 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1630_0 <=( _mesh_29_18_io_out_valid_0) ^ ((fiEnable && (6767 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1631_0 <=( _mesh_30_18_io_out_valid_0) ^ ((fiEnable && (6768 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1632_0 <=( io_in_valid_19_0) ^ ((fiEnable && (6769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1633_0 <=( _mesh_0_19_io_out_valid_0) ^ ((fiEnable && (6770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1634_0 <=( _mesh_1_19_io_out_valid_0) ^ ((fiEnable && (6771 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1635_0 <=( _mesh_2_19_io_out_valid_0) ^ ((fiEnable && (6772 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1636_0 <=( _mesh_3_19_io_out_valid_0) ^ ((fiEnable && (6773 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1637_0 <=( _mesh_4_19_io_out_valid_0) ^ ((fiEnable && (6774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1638_0 <=( _mesh_5_19_io_out_valid_0) ^ ((fiEnable && (6775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1639_0 <=( _mesh_6_19_io_out_valid_0) ^ ((fiEnable && (6776 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1640_0 <=( _mesh_7_19_io_out_valid_0) ^ ((fiEnable && (6777 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1641_0 <=( _mesh_8_19_io_out_valid_0) ^ ((fiEnable && (6778 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1642_0 <=( _mesh_9_19_io_out_valid_0) ^ ((fiEnable && (6779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1643_0 <=( _mesh_10_19_io_out_valid_0) ^ ((fiEnable && (6780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1644_0 <=( _mesh_11_19_io_out_valid_0) ^ ((fiEnable && (6781 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1645_0 <=( _mesh_12_19_io_out_valid_0) ^ ((fiEnable && (6782 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1646_0 <=( _mesh_13_19_io_out_valid_0) ^ ((fiEnable && (6783 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1647_0 <=( _mesh_14_19_io_out_valid_0) ^ ((fiEnable && (6784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1648_0 <=( _mesh_15_19_io_out_valid_0) ^ ((fiEnable && (6785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1649_0 <=( _mesh_16_19_io_out_valid_0) ^ ((fiEnable && (6786 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1650_0 <=( _mesh_17_19_io_out_valid_0) ^ ((fiEnable && (6787 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1651_0 <=( _mesh_18_19_io_out_valid_0) ^ ((fiEnable && (6788 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1652_0 <=( _mesh_19_19_io_out_valid_0) ^ ((fiEnable && (6789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1653_0 <=( _mesh_20_19_io_out_valid_0) ^ ((fiEnable && (6790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1654_0 <=( _mesh_21_19_io_out_valid_0) ^ ((fiEnable && (6791 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1655_0 <=( _mesh_22_19_io_out_valid_0) ^ ((fiEnable && (6792 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1656_0 <=( _mesh_23_19_io_out_valid_0) ^ ((fiEnable && (6793 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1657_0 <=( _mesh_24_19_io_out_valid_0) ^ ((fiEnable && (6794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1658_0 <=( _mesh_25_19_io_out_valid_0) ^ ((fiEnable && (6795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1659_0 <=( _mesh_26_19_io_out_valid_0) ^ ((fiEnable && (6796 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1660_0 <=( _mesh_27_19_io_out_valid_0) ^ ((fiEnable && (6797 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1661_0 <=( _mesh_28_19_io_out_valid_0) ^ ((fiEnable && (6798 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1662_0 <=( _mesh_29_19_io_out_valid_0) ^ ((fiEnable && (6799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1663_0 <=( _mesh_30_19_io_out_valid_0) ^ ((fiEnable && (6800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1664_0 <=( io_in_valid_20_0) ^ ((fiEnable && (6801 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1665_0 <=( _mesh_0_20_io_out_valid_0) ^ ((fiEnable && (6802 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1666_0 <=( _mesh_1_20_io_out_valid_0) ^ ((fiEnable && (6803 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1667_0 <=( _mesh_2_20_io_out_valid_0) ^ ((fiEnable && (6804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1668_0 <=( _mesh_3_20_io_out_valid_0) ^ ((fiEnable && (6805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1669_0 <=( _mesh_4_20_io_out_valid_0) ^ ((fiEnable && (6806 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1670_0 <=( _mesh_5_20_io_out_valid_0) ^ ((fiEnable && (6807 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1671_0 <=( _mesh_6_20_io_out_valid_0) ^ ((fiEnable && (6808 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1672_0 <=( _mesh_7_20_io_out_valid_0) ^ ((fiEnable && (6809 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1673_0 <=( _mesh_8_20_io_out_valid_0) ^ ((fiEnable && (6810 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1674_0 <=( _mesh_9_20_io_out_valid_0) ^ ((fiEnable && (6811 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1675_0 <=( _mesh_10_20_io_out_valid_0) ^ ((fiEnable && (6812 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1676_0 <=( _mesh_11_20_io_out_valid_0) ^ ((fiEnable && (6813 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1677_0 <=( _mesh_12_20_io_out_valid_0) ^ ((fiEnable && (6814 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1678_0 <=( _mesh_13_20_io_out_valid_0) ^ ((fiEnable && (6815 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1679_0 <=( _mesh_14_20_io_out_valid_0) ^ ((fiEnable && (6816 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1680_0 <=( _mesh_15_20_io_out_valid_0) ^ ((fiEnable && (6817 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1681_0 <=( _mesh_16_20_io_out_valid_0) ^ ((fiEnable && (6818 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1682_0 <=( _mesh_17_20_io_out_valid_0) ^ ((fiEnable && (6819 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1683_0 <=( _mesh_18_20_io_out_valid_0) ^ ((fiEnable && (6820 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1684_0 <=( _mesh_19_20_io_out_valid_0) ^ ((fiEnable && (6821 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1685_0 <=( _mesh_20_20_io_out_valid_0) ^ ((fiEnable && (6822 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1686_0 <=( _mesh_21_20_io_out_valid_0) ^ ((fiEnable && (6823 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1687_0 <=( _mesh_22_20_io_out_valid_0) ^ ((fiEnable && (6824 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1688_0 <=( _mesh_23_20_io_out_valid_0) ^ ((fiEnable && (6825 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1689_0 <=( _mesh_24_20_io_out_valid_0) ^ ((fiEnable && (6826 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1690_0 <=( _mesh_25_20_io_out_valid_0) ^ ((fiEnable && (6827 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1691_0 <=( _mesh_26_20_io_out_valid_0) ^ ((fiEnable && (6828 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1692_0 <=( _mesh_27_20_io_out_valid_0) ^ ((fiEnable && (6829 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1693_0 <=( _mesh_28_20_io_out_valid_0) ^ ((fiEnable && (6830 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1694_0 <=( _mesh_29_20_io_out_valid_0) ^ ((fiEnable && (6831 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1695_0 <=( _mesh_30_20_io_out_valid_0) ^ ((fiEnable && (6832 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1696_0 <=( io_in_valid_21_0) ^ ((fiEnable && (6833 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1697_0 <=( _mesh_0_21_io_out_valid_0) ^ ((fiEnable && (6834 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1698_0 <=( _mesh_1_21_io_out_valid_0) ^ ((fiEnable && (6835 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1699_0 <=( _mesh_2_21_io_out_valid_0) ^ ((fiEnable && (6836 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1700_0 <=( _mesh_3_21_io_out_valid_0) ^ ((fiEnable && (6837 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1701_0 <=( _mesh_4_21_io_out_valid_0) ^ ((fiEnable && (6838 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1702_0 <=( _mesh_5_21_io_out_valid_0) ^ ((fiEnable && (6839 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1703_0 <=( _mesh_6_21_io_out_valid_0) ^ ((fiEnable && (6840 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1704_0 <=( _mesh_7_21_io_out_valid_0) ^ ((fiEnable && (6841 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1705_0 <=( _mesh_8_21_io_out_valid_0) ^ ((fiEnable && (6842 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1706_0 <=( _mesh_9_21_io_out_valid_0) ^ ((fiEnable && (6843 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1707_0 <=( _mesh_10_21_io_out_valid_0) ^ ((fiEnable && (6844 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1708_0 <=( _mesh_11_21_io_out_valid_0) ^ ((fiEnable && (6845 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1709_0 <=( _mesh_12_21_io_out_valid_0) ^ ((fiEnable && (6846 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1710_0 <=( _mesh_13_21_io_out_valid_0) ^ ((fiEnable && (6847 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1711_0 <=( _mesh_14_21_io_out_valid_0) ^ ((fiEnable && (6848 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1712_0 <=( _mesh_15_21_io_out_valid_0) ^ ((fiEnable && (6849 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1713_0 <=( _mesh_16_21_io_out_valid_0) ^ ((fiEnable && (6850 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1714_0 <=( _mesh_17_21_io_out_valid_0) ^ ((fiEnable && (6851 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1715_0 <=( _mesh_18_21_io_out_valid_0) ^ ((fiEnable && (6852 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1716_0 <=( _mesh_19_21_io_out_valid_0) ^ ((fiEnable && (6853 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1717_0 <=( _mesh_20_21_io_out_valid_0) ^ ((fiEnable && (6854 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1718_0 <=( _mesh_21_21_io_out_valid_0) ^ ((fiEnable && (6855 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1719_0 <=( _mesh_22_21_io_out_valid_0) ^ ((fiEnable && (6856 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1720_0 <=( _mesh_23_21_io_out_valid_0) ^ ((fiEnable && (6857 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1721_0 <=( _mesh_24_21_io_out_valid_0) ^ ((fiEnable && (6858 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1722_0 <=( _mesh_25_21_io_out_valid_0) ^ ((fiEnable && (6859 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1723_0 <=( _mesh_26_21_io_out_valid_0) ^ ((fiEnable && (6860 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1724_0 <=( _mesh_27_21_io_out_valid_0) ^ ((fiEnable && (6861 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1725_0 <=( _mesh_28_21_io_out_valid_0) ^ ((fiEnable && (6862 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1726_0 <=( _mesh_29_21_io_out_valid_0) ^ ((fiEnable && (6863 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1727_0 <=( _mesh_30_21_io_out_valid_0) ^ ((fiEnable && (6864 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1728_0 <=( io_in_valid_22_0) ^ ((fiEnable && (6865 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1729_0 <=( _mesh_0_22_io_out_valid_0) ^ ((fiEnable && (6866 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1730_0 <=( _mesh_1_22_io_out_valid_0) ^ ((fiEnable && (6867 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1731_0 <=( _mesh_2_22_io_out_valid_0) ^ ((fiEnable && (6868 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1732_0 <=( _mesh_3_22_io_out_valid_0) ^ ((fiEnable && (6869 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1733_0 <=( _mesh_4_22_io_out_valid_0) ^ ((fiEnable && (6870 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1734_0 <=( _mesh_5_22_io_out_valid_0) ^ ((fiEnable && (6871 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1735_0 <=( _mesh_6_22_io_out_valid_0) ^ ((fiEnable && (6872 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1736_0 <=( _mesh_7_22_io_out_valid_0) ^ ((fiEnable && (6873 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1737_0 <=( _mesh_8_22_io_out_valid_0) ^ ((fiEnable && (6874 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1738_0 <=( _mesh_9_22_io_out_valid_0) ^ ((fiEnable && (6875 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1739_0 <=( _mesh_10_22_io_out_valid_0) ^ ((fiEnable && (6876 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1740_0 <=( _mesh_11_22_io_out_valid_0) ^ ((fiEnable && (6877 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1741_0 <=( _mesh_12_22_io_out_valid_0) ^ ((fiEnable && (6878 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1742_0 <=( _mesh_13_22_io_out_valid_0) ^ ((fiEnable && (6879 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1743_0 <=( _mesh_14_22_io_out_valid_0) ^ ((fiEnable && (6880 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1744_0 <=( _mesh_15_22_io_out_valid_0) ^ ((fiEnable && (6881 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1745_0 <=( _mesh_16_22_io_out_valid_0) ^ ((fiEnable && (6882 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1746_0 <=( _mesh_17_22_io_out_valid_0) ^ ((fiEnable && (6883 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1747_0 <=( _mesh_18_22_io_out_valid_0) ^ ((fiEnable && (6884 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1748_0 <=( _mesh_19_22_io_out_valid_0) ^ ((fiEnable && (6885 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1749_0 <=( _mesh_20_22_io_out_valid_0) ^ ((fiEnable && (6886 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1750_0 <=( _mesh_21_22_io_out_valid_0) ^ ((fiEnable && (6887 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1751_0 <=( _mesh_22_22_io_out_valid_0) ^ ((fiEnable && (6888 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1752_0 <=( _mesh_23_22_io_out_valid_0) ^ ((fiEnable && (6889 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1753_0 <=( _mesh_24_22_io_out_valid_0) ^ ((fiEnable && (6890 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1754_0 <=( _mesh_25_22_io_out_valid_0) ^ ((fiEnable && (6891 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1755_0 <=( _mesh_26_22_io_out_valid_0) ^ ((fiEnable && (6892 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1756_0 <=( _mesh_27_22_io_out_valid_0) ^ ((fiEnable && (6893 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1757_0 <=( _mesh_28_22_io_out_valid_0) ^ ((fiEnable && (6894 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1758_0 <=( _mesh_29_22_io_out_valid_0) ^ ((fiEnable && (6895 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1759_0 <=( _mesh_30_22_io_out_valid_0) ^ ((fiEnable && (6896 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1760_0 <=( io_in_valid_23_0) ^ ((fiEnable && (6897 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1761_0 <=( _mesh_0_23_io_out_valid_0) ^ ((fiEnable && (6898 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1762_0 <=( _mesh_1_23_io_out_valid_0) ^ ((fiEnable && (6899 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1763_0 <=( _mesh_2_23_io_out_valid_0) ^ ((fiEnable && (6900 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1764_0 <=( _mesh_3_23_io_out_valid_0) ^ ((fiEnable && (6901 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1765_0 <=( _mesh_4_23_io_out_valid_0) ^ ((fiEnable && (6902 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1766_0 <=( _mesh_5_23_io_out_valid_0) ^ ((fiEnable && (6903 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1767_0 <=( _mesh_6_23_io_out_valid_0) ^ ((fiEnable && (6904 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1768_0 <=( _mesh_7_23_io_out_valid_0) ^ ((fiEnable && (6905 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1769_0 <=( _mesh_8_23_io_out_valid_0) ^ ((fiEnable && (6906 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1770_0 <=( _mesh_9_23_io_out_valid_0) ^ ((fiEnable && (6907 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1771_0 <=( _mesh_10_23_io_out_valid_0) ^ ((fiEnable && (6908 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1772_0 <=( _mesh_11_23_io_out_valid_0) ^ ((fiEnable && (6909 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1773_0 <=( _mesh_12_23_io_out_valid_0) ^ ((fiEnable && (6910 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1774_0 <=( _mesh_13_23_io_out_valid_0) ^ ((fiEnable && (6911 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1775_0 <=( _mesh_14_23_io_out_valid_0) ^ ((fiEnable && (6912 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1776_0 <=( _mesh_15_23_io_out_valid_0) ^ ((fiEnable && (6913 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1777_0 <=( _mesh_16_23_io_out_valid_0) ^ ((fiEnable && (6914 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1778_0 <=( _mesh_17_23_io_out_valid_0) ^ ((fiEnable && (6915 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1779_0 <=( _mesh_18_23_io_out_valid_0) ^ ((fiEnable && (6916 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1780_0 <=( _mesh_19_23_io_out_valid_0) ^ ((fiEnable && (6917 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1781_0 <=( _mesh_20_23_io_out_valid_0) ^ ((fiEnable && (6918 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1782_0 <=( _mesh_21_23_io_out_valid_0) ^ ((fiEnable && (6919 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1783_0 <=( _mesh_22_23_io_out_valid_0) ^ ((fiEnable && (6920 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1784_0 <=( _mesh_23_23_io_out_valid_0) ^ ((fiEnable && (6921 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1785_0 <=( _mesh_24_23_io_out_valid_0) ^ ((fiEnable && (6922 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1786_0 <=( _mesh_25_23_io_out_valid_0) ^ ((fiEnable && (6923 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1787_0 <=( _mesh_26_23_io_out_valid_0) ^ ((fiEnable && (6924 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1788_0 <=( _mesh_27_23_io_out_valid_0) ^ ((fiEnable && (6925 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1789_0 <=( _mesh_28_23_io_out_valid_0) ^ ((fiEnable && (6926 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1790_0 <=( _mesh_29_23_io_out_valid_0) ^ ((fiEnable && (6927 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1791_0 <=( _mesh_30_23_io_out_valid_0) ^ ((fiEnable && (6928 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1792_0 <=( io_in_valid_24_0) ^ ((fiEnable && (6929 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1793_0 <=( _mesh_0_24_io_out_valid_0) ^ ((fiEnable && (6930 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1794_0 <=( _mesh_1_24_io_out_valid_0) ^ ((fiEnable && (6931 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1795_0 <=( _mesh_2_24_io_out_valid_0) ^ ((fiEnable && (6932 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1796_0 <=( _mesh_3_24_io_out_valid_0) ^ ((fiEnable && (6933 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1797_0 <=( _mesh_4_24_io_out_valid_0) ^ ((fiEnable && (6934 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1798_0 <=( _mesh_5_24_io_out_valid_0) ^ ((fiEnable && (6935 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1799_0 <=( _mesh_6_24_io_out_valid_0) ^ ((fiEnable && (6936 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1800_0 <=( _mesh_7_24_io_out_valid_0) ^ ((fiEnable && (6937 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1801_0 <=( _mesh_8_24_io_out_valid_0) ^ ((fiEnable && (6938 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1802_0 <=( _mesh_9_24_io_out_valid_0) ^ ((fiEnable && (6939 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1803_0 <=( _mesh_10_24_io_out_valid_0) ^ ((fiEnable && (6940 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1804_0 <=( _mesh_11_24_io_out_valid_0) ^ ((fiEnable && (6941 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1805_0 <=( _mesh_12_24_io_out_valid_0) ^ ((fiEnable && (6942 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1806_0 <=( _mesh_13_24_io_out_valid_0) ^ ((fiEnable && (6943 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1807_0 <=( _mesh_14_24_io_out_valid_0) ^ ((fiEnable && (6944 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1808_0 <=( _mesh_15_24_io_out_valid_0) ^ ((fiEnable && (6945 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1809_0 <=( _mesh_16_24_io_out_valid_0) ^ ((fiEnable && (6946 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1810_0 <=( _mesh_17_24_io_out_valid_0) ^ ((fiEnable && (6947 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1811_0 <=( _mesh_18_24_io_out_valid_0) ^ ((fiEnable && (6948 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1812_0 <=( _mesh_19_24_io_out_valid_0) ^ ((fiEnable && (6949 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1813_0 <=( _mesh_20_24_io_out_valid_0) ^ ((fiEnable && (6950 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1814_0 <=( _mesh_21_24_io_out_valid_0) ^ ((fiEnable && (6951 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1815_0 <=( _mesh_22_24_io_out_valid_0) ^ ((fiEnable && (6952 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1816_0 <=( _mesh_23_24_io_out_valid_0) ^ ((fiEnable && (6953 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1817_0 <=( _mesh_24_24_io_out_valid_0) ^ ((fiEnable && (6954 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1818_0 <=( _mesh_25_24_io_out_valid_0) ^ ((fiEnable && (6955 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1819_0 <=( _mesh_26_24_io_out_valid_0) ^ ((fiEnable && (6956 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1820_0 <=( _mesh_27_24_io_out_valid_0) ^ ((fiEnable && (6957 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1821_0 <=( _mesh_28_24_io_out_valid_0) ^ ((fiEnable && (6958 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1822_0 <=( _mesh_29_24_io_out_valid_0) ^ ((fiEnable && (6959 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1823_0 <=( _mesh_30_24_io_out_valid_0) ^ ((fiEnable && (6960 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1824_0 <=( io_in_valid_25_0) ^ ((fiEnable && (6961 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1825_0 <=( _mesh_0_25_io_out_valid_0) ^ ((fiEnable && (6962 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1826_0 <=( _mesh_1_25_io_out_valid_0) ^ ((fiEnable && (6963 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1827_0 <=( _mesh_2_25_io_out_valid_0) ^ ((fiEnable && (6964 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1828_0 <=( _mesh_3_25_io_out_valid_0) ^ ((fiEnable && (6965 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1829_0 <=( _mesh_4_25_io_out_valid_0) ^ ((fiEnable && (6966 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1830_0 <=( _mesh_5_25_io_out_valid_0) ^ ((fiEnable && (6967 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1831_0 <=( _mesh_6_25_io_out_valid_0) ^ ((fiEnable && (6968 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1832_0 <=( _mesh_7_25_io_out_valid_0) ^ ((fiEnable && (6969 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1833_0 <=( _mesh_8_25_io_out_valid_0) ^ ((fiEnable && (6970 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1834_0 <=( _mesh_9_25_io_out_valid_0) ^ ((fiEnable && (6971 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1835_0 <=( _mesh_10_25_io_out_valid_0) ^ ((fiEnable && (6972 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1836_0 <=( _mesh_11_25_io_out_valid_0) ^ ((fiEnable && (6973 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1837_0 <=( _mesh_12_25_io_out_valid_0) ^ ((fiEnable && (6974 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1838_0 <=( _mesh_13_25_io_out_valid_0) ^ ((fiEnable && (6975 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1839_0 <=( _mesh_14_25_io_out_valid_0) ^ ((fiEnable && (6976 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1840_0 <=( _mesh_15_25_io_out_valid_0) ^ ((fiEnable && (6977 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1841_0 <=( _mesh_16_25_io_out_valid_0) ^ ((fiEnable && (6978 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1842_0 <=( _mesh_17_25_io_out_valid_0) ^ ((fiEnable && (6979 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1843_0 <=( _mesh_18_25_io_out_valid_0) ^ ((fiEnable && (6980 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1844_0 <=( _mesh_19_25_io_out_valid_0) ^ ((fiEnable && (6981 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1845_0 <=( _mesh_20_25_io_out_valid_0) ^ ((fiEnable && (6982 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1846_0 <=( _mesh_21_25_io_out_valid_0) ^ ((fiEnable && (6983 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1847_0 <=( _mesh_22_25_io_out_valid_0) ^ ((fiEnable && (6984 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1848_0 <=( _mesh_23_25_io_out_valid_0) ^ ((fiEnable && (6985 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1849_0 <=( _mesh_24_25_io_out_valid_0) ^ ((fiEnable && (6986 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1850_0 <=( _mesh_25_25_io_out_valid_0) ^ ((fiEnable && (6987 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1851_0 <=( _mesh_26_25_io_out_valid_0) ^ ((fiEnable && (6988 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1852_0 <=( _mesh_27_25_io_out_valid_0) ^ ((fiEnable && (6989 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1853_0 <=( _mesh_28_25_io_out_valid_0) ^ ((fiEnable && (6990 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1854_0 <=( _mesh_29_25_io_out_valid_0) ^ ((fiEnable && (6991 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1855_0 <=( _mesh_30_25_io_out_valid_0) ^ ((fiEnable && (6992 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1856_0 <=( io_in_valid_26_0) ^ ((fiEnable && (6993 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1857_0 <=( _mesh_0_26_io_out_valid_0) ^ ((fiEnable && (6994 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1858_0 <=( _mesh_1_26_io_out_valid_0) ^ ((fiEnable && (6995 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1859_0 <=( _mesh_2_26_io_out_valid_0) ^ ((fiEnable && (6996 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1860_0 <=( _mesh_3_26_io_out_valid_0) ^ ((fiEnable && (6997 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1861_0 <=( _mesh_4_26_io_out_valid_0) ^ ((fiEnable && (6998 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1862_0 <=( _mesh_5_26_io_out_valid_0) ^ ((fiEnable && (6999 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1863_0 <=( _mesh_6_26_io_out_valid_0) ^ ((fiEnable && (7000 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1864_0 <=( _mesh_7_26_io_out_valid_0) ^ ((fiEnable && (7001 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1865_0 <=( _mesh_8_26_io_out_valid_0) ^ ((fiEnable && (7002 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1866_0 <=( _mesh_9_26_io_out_valid_0) ^ ((fiEnable && (7003 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1867_0 <=( _mesh_10_26_io_out_valid_0) ^ ((fiEnable && (7004 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1868_0 <=( _mesh_11_26_io_out_valid_0) ^ ((fiEnable && (7005 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1869_0 <=( _mesh_12_26_io_out_valid_0) ^ ((fiEnable && (7006 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1870_0 <=( _mesh_13_26_io_out_valid_0) ^ ((fiEnable && (7007 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1871_0 <=( _mesh_14_26_io_out_valid_0) ^ ((fiEnable && (7008 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1872_0 <=( _mesh_15_26_io_out_valid_0) ^ ((fiEnable && (7009 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1873_0 <=( _mesh_16_26_io_out_valid_0) ^ ((fiEnable && (7010 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1874_0 <=( _mesh_17_26_io_out_valid_0) ^ ((fiEnable && (7011 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1875_0 <=( _mesh_18_26_io_out_valid_0) ^ ((fiEnable && (7012 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1876_0 <=( _mesh_19_26_io_out_valid_0) ^ ((fiEnable && (7013 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1877_0 <=( _mesh_20_26_io_out_valid_0) ^ ((fiEnable && (7014 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1878_0 <=( _mesh_21_26_io_out_valid_0) ^ ((fiEnable && (7015 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1879_0 <=( _mesh_22_26_io_out_valid_0) ^ ((fiEnable && (7016 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1880_0 <=( _mesh_23_26_io_out_valid_0) ^ ((fiEnable && (7017 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1881_0 <=( _mesh_24_26_io_out_valid_0) ^ ((fiEnable && (7018 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1882_0 <=( _mesh_25_26_io_out_valid_0) ^ ((fiEnable && (7019 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1883_0 <=( _mesh_26_26_io_out_valid_0) ^ ((fiEnable && (7020 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1884_0 <=( _mesh_27_26_io_out_valid_0) ^ ((fiEnable && (7021 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1885_0 <=( _mesh_28_26_io_out_valid_0) ^ ((fiEnable && (7022 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1886_0 <=( _mesh_29_26_io_out_valid_0) ^ ((fiEnable && (7023 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1887_0 <=( _mesh_30_26_io_out_valid_0) ^ ((fiEnable && (7024 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1888_0 <=( io_in_valid_27_0) ^ ((fiEnable && (7025 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1889_0 <=( _mesh_0_27_io_out_valid_0) ^ ((fiEnable && (7026 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1890_0 <=( _mesh_1_27_io_out_valid_0) ^ ((fiEnable && (7027 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1891_0 <=( _mesh_2_27_io_out_valid_0) ^ ((fiEnable && (7028 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1892_0 <=( _mesh_3_27_io_out_valid_0) ^ ((fiEnable && (7029 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1893_0 <=( _mesh_4_27_io_out_valid_0) ^ ((fiEnable && (7030 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1894_0 <=( _mesh_5_27_io_out_valid_0) ^ ((fiEnable && (7031 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1895_0 <=( _mesh_6_27_io_out_valid_0) ^ ((fiEnable && (7032 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1896_0 <=( _mesh_7_27_io_out_valid_0) ^ ((fiEnable && (7033 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1897_0 <=( _mesh_8_27_io_out_valid_0) ^ ((fiEnable && (7034 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1898_0 <=( _mesh_9_27_io_out_valid_0) ^ ((fiEnable && (7035 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1899_0 <=( _mesh_10_27_io_out_valid_0) ^ ((fiEnable && (7036 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1900_0 <=( _mesh_11_27_io_out_valid_0) ^ ((fiEnable && (7037 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1901_0 <=( _mesh_12_27_io_out_valid_0) ^ ((fiEnable && (7038 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1902_0 <=( _mesh_13_27_io_out_valid_0) ^ ((fiEnable && (7039 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1903_0 <=( _mesh_14_27_io_out_valid_0) ^ ((fiEnable && (7040 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1904_0 <=( _mesh_15_27_io_out_valid_0) ^ ((fiEnable && (7041 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1905_0 <=( _mesh_16_27_io_out_valid_0) ^ ((fiEnable && (7042 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1906_0 <=( _mesh_17_27_io_out_valid_0) ^ ((fiEnable && (7043 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1907_0 <=( _mesh_18_27_io_out_valid_0) ^ ((fiEnable && (7044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1908_0 <=( _mesh_19_27_io_out_valid_0) ^ ((fiEnable && (7045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1909_0 <=( _mesh_20_27_io_out_valid_0) ^ ((fiEnable && (7046 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1910_0 <=( _mesh_21_27_io_out_valid_0) ^ ((fiEnable && (7047 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1911_0 <=( _mesh_22_27_io_out_valid_0) ^ ((fiEnable && (7048 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1912_0 <=( _mesh_23_27_io_out_valid_0) ^ ((fiEnable && (7049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1913_0 <=( _mesh_24_27_io_out_valid_0) ^ ((fiEnable && (7050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1914_0 <=( _mesh_25_27_io_out_valid_0) ^ ((fiEnable && (7051 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1915_0 <=( _mesh_26_27_io_out_valid_0) ^ ((fiEnable && (7052 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1916_0 <=( _mesh_27_27_io_out_valid_0) ^ ((fiEnable && (7053 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1917_0 <=( _mesh_28_27_io_out_valid_0) ^ ((fiEnable && (7054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1918_0 <=( _mesh_29_27_io_out_valid_0) ^ ((fiEnable && (7055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1919_0 <=( _mesh_30_27_io_out_valid_0) ^ ((fiEnable && (7056 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1920_0 <=( io_in_valid_28_0) ^ ((fiEnable && (7057 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1921_0 <=( _mesh_0_28_io_out_valid_0) ^ ((fiEnable && (7058 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1922_0 <=( _mesh_1_28_io_out_valid_0) ^ ((fiEnable && (7059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1923_0 <=( _mesh_2_28_io_out_valid_0) ^ ((fiEnable && (7060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1924_0 <=( _mesh_3_28_io_out_valid_0) ^ ((fiEnable && (7061 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1925_0 <=( _mesh_4_28_io_out_valid_0) ^ ((fiEnable && (7062 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1926_0 <=( _mesh_5_28_io_out_valid_0) ^ ((fiEnable && (7063 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1927_0 <=( _mesh_6_28_io_out_valid_0) ^ ((fiEnable && (7064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1928_0 <=( _mesh_7_28_io_out_valid_0) ^ ((fiEnable && (7065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1929_0 <=( _mesh_8_28_io_out_valid_0) ^ ((fiEnable && (7066 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1930_0 <=( _mesh_9_28_io_out_valid_0) ^ ((fiEnable && (7067 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1931_0 <=( _mesh_10_28_io_out_valid_0) ^ ((fiEnable && (7068 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1932_0 <=( _mesh_11_28_io_out_valid_0) ^ ((fiEnable && (7069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1933_0 <=( _mesh_12_28_io_out_valid_0) ^ ((fiEnable && (7070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1934_0 <=( _mesh_13_28_io_out_valid_0) ^ ((fiEnable && (7071 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1935_0 <=( _mesh_14_28_io_out_valid_0) ^ ((fiEnable && (7072 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1936_0 <=( _mesh_15_28_io_out_valid_0) ^ ((fiEnable && (7073 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1937_0 <=( _mesh_16_28_io_out_valid_0) ^ ((fiEnable && (7074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1938_0 <=( _mesh_17_28_io_out_valid_0) ^ ((fiEnable && (7075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1939_0 <=( _mesh_18_28_io_out_valid_0) ^ ((fiEnable && (7076 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1940_0 <=( _mesh_19_28_io_out_valid_0) ^ ((fiEnable && (7077 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1941_0 <=( _mesh_20_28_io_out_valid_0) ^ ((fiEnable && (7078 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1942_0 <=( _mesh_21_28_io_out_valid_0) ^ ((fiEnable && (7079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1943_0 <=( _mesh_22_28_io_out_valid_0) ^ ((fiEnable && (7080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1944_0 <=( _mesh_23_28_io_out_valid_0) ^ ((fiEnable && (7081 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1945_0 <=( _mesh_24_28_io_out_valid_0) ^ ((fiEnable && (7082 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1946_0 <=( _mesh_25_28_io_out_valid_0) ^ ((fiEnable && (7083 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1947_0 <=( _mesh_26_28_io_out_valid_0) ^ ((fiEnable && (7084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1948_0 <=( _mesh_27_28_io_out_valid_0) ^ ((fiEnable && (7085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1949_0 <=( _mesh_28_28_io_out_valid_0) ^ ((fiEnable && (7086 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1950_0 <=( _mesh_29_28_io_out_valid_0) ^ ((fiEnable && (7087 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1951_0 <=( _mesh_30_28_io_out_valid_0) ^ ((fiEnable && (7088 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1952_0 <=( io_in_valid_29_0) ^ ((fiEnable && (7089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1953_0 <=( _mesh_0_29_io_out_valid_0) ^ ((fiEnable && (7090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1954_0 <=( _mesh_1_29_io_out_valid_0) ^ ((fiEnable && (7091 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1955_0 <=( _mesh_2_29_io_out_valid_0) ^ ((fiEnable && (7092 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1956_0 <=( _mesh_3_29_io_out_valid_0) ^ ((fiEnable && (7093 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1957_0 <=( _mesh_4_29_io_out_valid_0) ^ ((fiEnable && (7094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1958_0 <=( _mesh_5_29_io_out_valid_0) ^ ((fiEnable && (7095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1959_0 <=( _mesh_6_29_io_out_valid_0) ^ ((fiEnable && (7096 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1960_0 <=( _mesh_7_29_io_out_valid_0) ^ ((fiEnable && (7097 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1961_0 <=( _mesh_8_29_io_out_valid_0) ^ ((fiEnable && (7098 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1962_0 <=( _mesh_9_29_io_out_valid_0) ^ ((fiEnable && (7099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1963_0 <=( _mesh_10_29_io_out_valid_0) ^ ((fiEnable && (7100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1964_0 <=( _mesh_11_29_io_out_valid_0) ^ ((fiEnable && (7101 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1965_0 <=( _mesh_12_29_io_out_valid_0) ^ ((fiEnable && (7102 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1966_0 <=( _mesh_13_29_io_out_valid_0) ^ ((fiEnable && (7103 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1967_0 <=( _mesh_14_29_io_out_valid_0) ^ ((fiEnable && (7104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1968_0 <=( _mesh_15_29_io_out_valid_0) ^ ((fiEnable && (7105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1969_0 <=( _mesh_16_29_io_out_valid_0) ^ ((fiEnable && (7106 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1970_0 <=( _mesh_17_29_io_out_valid_0) ^ ((fiEnable && (7107 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1971_0 <=( _mesh_18_29_io_out_valid_0) ^ ((fiEnable && (7108 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1972_0 <=( _mesh_19_29_io_out_valid_0) ^ ((fiEnable && (7109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1973_0 <=( _mesh_20_29_io_out_valid_0) ^ ((fiEnable && (7110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1974_0 <=( _mesh_21_29_io_out_valid_0) ^ ((fiEnable && (7111 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1975_0 <=( _mesh_22_29_io_out_valid_0) ^ ((fiEnable && (7112 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1976_0 <=( _mesh_23_29_io_out_valid_0) ^ ((fiEnable && (7113 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1977_0 <=( _mesh_24_29_io_out_valid_0) ^ ((fiEnable && (7114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1978_0 <=( _mesh_25_29_io_out_valid_0) ^ ((fiEnable && (7115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1979_0 <=( _mesh_26_29_io_out_valid_0) ^ ((fiEnable && (7116 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1980_0 <=( _mesh_27_29_io_out_valid_0) ^ ((fiEnable && (7117 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1981_0 <=( _mesh_28_29_io_out_valid_0) ^ ((fiEnable && (7118 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1982_0 <=( _mesh_29_29_io_out_valid_0) ^ ((fiEnable && (7119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1983_0 <=( _mesh_30_29_io_out_valid_0) ^ ((fiEnable && (7120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1984_0 <=( io_in_valid_30_0) ^ ((fiEnable && (7121 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1985_0 <=( _mesh_0_30_io_out_valid_0) ^ ((fiEnable && (7122 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1986_0 <=( _mesh_1_30_io_out_valid_0) ^ ((fiEnable && (7123 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1987_0 <=( _mesh_2_30_io_out_valid_0) ^ ((fiEnable && (7124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1988_0 <=( _mesh_3_30_io_out_valid_0) ^ ((fiEnable && (7125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1989_0 <=( _mesh_4_30_io_out_valid_0) ^ ((fiEnable && (7126 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1990_0 <=( _mesh_5_30_io_out_valid_0) ^ ((fiEnable && (7127 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1991_0 <=( _mesh_6_30_io_out_valid_0) ^ ((fiEnable && (7128 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1992_0 <=( _mesh_7_30_io_out_valid_0) ^ ((fiEnable && (7129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1993_0 <=( _mesh_8_30_io_out_valid_0) ^ ((fiEnable && (7130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1994_0 <=( _mesh_9_30_io_out_valid_0) ^ ((fiEnable && (7131 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1995_0 <=( _mesh_10_30_io_out_valid_0) ^ ((fiEnable && (7132 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1996_0 <=( _mesh_11_30_io_out_valid_0) ^ ((fiEnable && (7133 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1997_0 <=( _mesh_12_30_io_out_valid_0) ^ ((fiEnable && (7134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1998_0 <=( _mesh_13_30_io_out_valid_0) ^ ((fiEnable && (7135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_1999_0 <=( _mesh_14_30_io_out_valid_0) ^ ((fiEnable && (7136 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2000_0 <=( _mesh_15_30_io_out_valid_0) ^ ((fiEnable && (7137 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2001_0 <=( _mesh_16_30_io_out_valid_0) ^ ((fiEnable && (7138 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2002_0 <=( _mesh_17_30_io_out_valid_0) ^ ((fiEnable && (7139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2003_0 <=( _mesh_18_30_io_out_valid_0) ^ ((fiEnable && (7140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2004_0 <=( _mesh_19_30_io_out_valid_0) ^ ((fiEnable && (7141 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2005_0 <=( _mesh_20_30_io_out_valid_0) ^ ((fiEnable && (7142 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2006_0 <=( _mesh_21_30_io_out_valid_0) ^ ((fiEnable && (7143 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2007_0 <=( _mesh_22_30_io_out_valid_0) ^ ((fiEnable && (7144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2008_0 <=( _mesh_23_30_io_out_valid_0) ^ ((fiEnable && (7145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2009_0 <=( _mesh_24_30_io_out_valid_0) ^ ((fiEnable && (7146 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2010_0 <=( _mesh_25_30_io_out_valid_0) ^ ((fiEnable && (7147 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2011_0 <=( _mesh_26_30_io_out_valid_0) ^ ((fiEnable && (7148 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2012_0 <=( _mesh_27_30_io_out_valid_0) ^ ((fiEnable && (7149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2013_0 <=( _mesh_28_30_io_out_valid_0) ^ ((fiEnable && (7150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2014_0 <=( _mesh_29_30_io_out_valid_0) ^ ((fiEnable && (7151 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2015_0 <=( _mesh_30_30_io_out_valid_0) ^ ((fiEnable && (7152 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2016_0 <=( io_in_valid_31_0) ^ ((fiEnable && (7153 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2017_0 <=( _mesh_0_31_io_out_valid_0) ^ ((fiEnable && (7154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2018_0 <=( _mesh_1_31_io_out_valid_0) ^ ((fiEnable && (7155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2019_0 <=( _mesh_2_31_io_out_valid_0) ^ ((fiEnable && (7156 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2020_0 <=( _mesh_3_31_io_out_valid_0) ^ ((fiEnable && (7157 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2021_0 <=( _mesh_4_31_io_out_valid_0) ^ ((fiEnable && (7158 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2022_0 <=( _mesh_5_31_io_out_valid_0) ^ ((fiEnable && (7159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2023_0 <=( _mesh_6_31_io_out_valid_0) ^ ((fiEnable && (7160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2024_0 <=( _mesh_7_31_io_out_valid_0) ^ ((fiEnable && (7161 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2025_0 <=( _mesh_8_31_io_out_valid_0) ^ ((fiEnable && (7162 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2026_0 <=( _mesh_9_31_io_out_valid_0) ^ ((fiEnable && (7163 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2027_0 <=( _mesh_10_31_io_out_valid_0) ^ ((fiEnable && (7164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2028_0 <=( _mesh_11_31_io_out_valid_0) ^ ((fiEnable && (7165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2029_0 <=( _mesh_12_31_io_out_valid_0) ^ ((fiEnable && (7166 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2030_0 <=( _mesh_13_31_io_out_valid_0) ^ ((fiEnable && (7167 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2031_0 <=( _mesh_14_31_io_out_valid_0) ^ ((fiEnable && (7168 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2032_0 <=( _mesh_15_31_io_out_valid_0) ^ ((fiEnable && (7169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2033_0 <=( _mesh_16_31_io_out_valid_0) ^ ((fiEnable && (7170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2034_0 <=( _mesh_17_31_io_out_valid_0) ^ ((fiEnable && (7171 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2035_0 <=( _mesh_18_31_io_out_valid_0) ^ ((fiEnable && (7172 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2036_0 <=( _mesh_19_31_io_out_valid_0) ^ ((fiEnable && (7173 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2037_0 <=( _mesh_20_31_io_out_valid_0) ^ ((fiEnable && (7174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2038_0 <=( _mesh_21_31_io_out_valid_0) ^ ((fiEnable && (7175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2039_0 <=( _mesh_22_31_io_out_valid_0) ^ ((fiEnable && (7176 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2040_0 <=( _mesh_23_31_io_out_valid_0) ^ ((fiEnable && (7177 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2041_0 <=( _mesh_24_31_io_out_valid_0) ^ ((fiEnable && (7178 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2042_0 <=( _mesh_25_31_io_out_valid_0) ^ ((fiEnable && (7179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2043_0 <=( _mesh_26_31_io_out_valid_0) ^ ((fiEnable && (7180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2044_0 <=( _mesh_27_31_io_out_valid_0) ^ ((fiEnable && (7181 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2045_0 <=( _mesh_28_31_io_out_valid_0) ^ ((fiEnable && (7182 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2046_0 <=( _mesh_29_31_io_out_valid_0) ^ ((fiEnable && (7183 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2047_0 <=( _mesh_30_31_io_out_valid_0) ^ ((fiEnable && (7184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_2048_0 <=( io_in_id_0_0) ^ ((fiEnable && (7185 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2049_0 <=( _mesh_0_0_io_out_id_0) ^ ((fiEnable && (7186 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2050_0 <=( _mesh_1_0_io_out_id_0) ^ ((fiEnable && (7187 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2051_0 <=( _mesh_2_0_io_out_id_0) ^ ((fiEnable && (7188 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2052_0 <=( _mesh_3_0_io_out_id_0) ^ ((fiEnable && (7189 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2053_0 <=( _mesh_4_0_io_out_id_0) ^ ((fiEnable && (7190 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2054_0 <=( _mesh_5_0_io_out_id_0) ^ ((fiEnable && (7191 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2055_0 <=( _mesh_6_0_io_out_id_0) ^ ((fiEnable && (7192 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2056_0 <=( _mesh_7_0_io_out_id_0) ^ ((fiEnable && (7193 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2057_0 <=( _mesh_8_0_io_out_id_0) ^ ((fiEnable && (7194 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2058_0 <=( _mesh_9_0_io_out_id_0) ^ ((fiEnable && (7195 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2059_0 <=( _mesh_10_0_io_out_id_0) ^ ((fiEnable && (7196 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2060_0 <=( _mesh_11_0_io_out_id_0) ^ ((fiEnable && (7197 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2061_0 <=( _mesh_12_0_io_out_id_0) ^ ((fiEnable && (7198 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2062_0 <=( _mesh_13_0_io_out_id_0) ^ ((fiEnable && (7199 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2063_0 <=( _mesh_14_0_io_out_id_0) ^ ((fiEnable && (7200 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2064_0 <=( _mesh_15_0_io_out_id_0) ^ ((fiEnable && (7201 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2065_0 <=( _mesh_16_0_io_out_id_0) ^ ((fiEnable && (7202 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2066_0 <=( _mesh_17_0_io_out_id_0) ^ ((fiEnable && (7203 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2067_0 <=( _mesh_18_0_io_out_id_0) ^ ((fiEnable && (7204 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2068_0 <=( _mesh_19_0_io_out_id_0) ^ ((fiEnable && (7205 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2069_0 <=( _mesh_20_0_io_out_id_0) ^ ((fiEnable && (7206 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2070_0 <=( _mesh_21_0_io_out_id_0) ^ ((fiEnable && (7207 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2071_0 <=( _mesh_22_0_io_out_id_0) ^ ((fiEnable && (7208 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2072_0 <=( _mesh_23_0_io_out_id_0) ^ ((fiEnable && (7209 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2073_0 <=( _mesh_24_0_io_out_id_0) ^ ((fiEnable && (7210 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2074_0 <=( _mesh_25_0_io_out_id_0) ^ ((fiEnable && (7211 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2075_0 <=( _mesh_26_0_io_out_id_0) ^ ((fiEnable && (7212 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2076_0 <=( _mesh_27_0_io_out_id_0) ^ ((fiEnable && (7213 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2077_0 <=( _mesh_28_0_io_out_id_0) ^ ((fiEnable && (7214 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2078_0 <=( _mesh_29_0_io_out_id_0) ^ ((fiEnable && (7215 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2079_0 <=( _mesh_30_0_io_out_id_0) ^ ((fiEnable && (7216 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2080_0 <=( io_in_id_1_0) ^ ((fiEnable && (7217 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2081_0 <=( _mesh_0_1_io_out_id_0) ^ ((fiEnable && (7218 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2082_0 <=( _mesh_1_1_io_out_id_0) ^ ((fiEnable && (7219 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2083_0 <=( _mesh_2_1_io_out_id_0) ^ ((fiEnable && (7220 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2084_0 <=( _mesh_3_1_io_out_id_0) ^ ((fiEnable && (7221 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2085_0 <=( _mesh_4_1_io_out_id_0) ^ ((fiEnable && (7222 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2086_0 <=( _mesh_5_1_io_out_id_0) ^ ((fiEnable && (7223 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2087_0 <=( _mesh_6_1_io_out_id_0) ^ ((fiEnable && (7224 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2088_0 <=( _mesh_7_1_io_out_id_0) ^ ((fiEnable && (7225 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2089_0 <=( _mesh_8_1_io_out_id_0) ^ ((fiEnable && (7226 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2090_0 <=( _mesh_9_1_io_out_id_0) ^ ((fiEnable && (7227 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2091_0 <=( _mesh_10_1_io_out_id_0) ^ ((fiEnable && (7228 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2092_0 <=( _mesh_11_1_io_out_id_0) ^ ((fiEnable && (7229 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2093_0 <=( _mesh_12_1_io_out_id_0) ^ ((fiEnable && (7230 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2094_0 <=( _mesh_13_1_io_out_id_0) ^ ((fiEnable && (7231 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2095_0 <=( _mesh_14_1_io_out_id_0) ^ ((fiEnable && (7232 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2096_0 <=( _mesh_15_1_io_out_id_0) ^ ((fiEnable && (7233 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2097_0 <=( _mesh_16_1_io_out_id_0) ^ ((fiEnable && (7234 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2098_0 <=( _mesh_17_1_io_out_id_0) ^ ((fiEnable && (7235 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2099_0 <=( _mesh_18_1_io_out_id_0) ^ ((fiEnable && (7236 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2100_0 <=( _mesh_19_1_io_out_id_0) ^ ((fiEnable && (7237 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2101_0 <=( _mesh_20_1_io_out_id_0) ^ ((fiEnable && (7238 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2102_0 <=( _mesh_21_1_io_out_id_0) ^ ((fiEnable && (7239 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2103_0 <=( _mesh_22_1_io_out_id_0) ^ ((fiEnable && (7240 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2104_0 <=( _mesh_23_1_io_out_id_0) ^ ((fiEnable && (7241 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2105_0 <=( _mesh_24_1_io_out_id_0) ^ ((fiEnable && (7242 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2106_0 <=( _mesh_25_1_io_out_id_0) ^ ((fiEnable && (7243 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2107_0 <=( _mesh_26_1_io_out_id_0) ^ ((fiEnable && (7244 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2108_0 <=( _mesh_27_1_io_out_id_0) ^ ((fiEnable && (7245 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2109_0 <=( _mesh_28_1_io_out_id_0) ^ ((fiEnable && (7246 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2110_0 <=( _mesh_29_1_io_out_id_0) ^ ((fiEnable && (7247 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2111_0 <=( _mesh_30_1_io_out_id_0) ^ ((fiEnable && (7248 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2112_0 <=( io_in_id_2_0) ^ ((fiEnable && (7249 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2113_0 <=( _mesh_0_2_io_out_id_0) ^ ((fiEnable && (7250 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2114_0 <=( _mesh_1_2_io_out_id_0) ^ ((fiEnable && (7251 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2115_0 <=( _mesh_2_2_io_out_id_0) ^ ((fiEnable && (7252 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2116_0 <=( _mesh_3_2_io_out_id_0) ^ ((fiEnable && (7253 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2117_0 <=( _mesh_4_2_io_out_id_0) ^ ((fiEnable && (7254 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2118_0 <=( _mesh_5_2_io_out_id_0) ^ ((fiEnable && (7255 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2119_0 <=( _mesh_6_2_io_out_id_0) ^ ((fiEnable && (7256 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2120_0 <=( _mesh_7_2_io_out_id_0) ^ ((fiEnable && (7257 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2121_0 <=( _mesh_8_2_io_out_id_0) ^ ((fiEnable && (7258 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2122_0 <=( _mesh_9_2_io_out_id_0) ^ ((fiEnable && (7259 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2123_0 <=( _mesh_10_2_io_out_id_0) ^ ((fiEnable && (7260 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2124_0 <=( _mesh_11_2_io_out_id_0) ^ ((fiEnable && (7261 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2125_0 <=( _mesh_12_2_io_out_id_0) ^ ((fiEnable && (7262 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2126_0 <=( _mesh_13_2_io_out_id_0) ^ ((fiEnable && (7263 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2127_0 <=( _mesh_14_2_io_out_id_0) ^ ((fiEnable && (7264 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2128_0 <=( _mesh_15_2_io_out_id_0) ^ ((fiEnable && (7265 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2129_0 <=( _mesh_16_2_io_out_id_0) ^ ((fiEnable && (7266 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2130_0 <=( _mesh_17_2_io_out_id_0) ^ ((fiEnable && (7267 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2131_0 <=( _mesh_18_2_io_out_id_0) ^ ((fiEnable && (7268 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2132_0 <=( _mesh_19_2_io_out_id_0) ^ ((fiEnable && (7269 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2133_0 <=( _mesh_20_2_io_out_id_0) ^ ((fiEnable && (7270 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2134_0 <=( _mesh_21_2_io_out_id_0) ^ ((fiEnable && (7271 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2135_0 <=( _mesh_22_2_io_out_id_0) ^ ((fiEnable && (7272 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2136_0 <=( _mesh_23_2_io_out_id_0) ^ ((fiEnable && (7273 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2137_0 <=( _mesh_24_2_io_out_id_0) ^ ((fiEnable && (7274 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2138_0 <=( _mesh_25_2_io_out_id_0) ^ ((fiEnable && (7275 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2139_0 <=( _mesh_26_2_io_out_id_0) ^ ((fiEnable && (7276 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2140_0 <=( _mesh_27_2_io_out_id_0) ^ ((fiEnable && (7277 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2141_0 <=( _mesh_28_2_io_out_id_0) ^ ((fiEnable && (7278 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2142_0 <=( _mesh_29_2_io_out_id_0) ^ ((fiEnable && (7279 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2143_0 <=( _mesh_30_2_io_out_id_0) ^ ((fiEnable && (7280 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2144_0 <=( io_in_id_3_0) ^ ((fiEnable && (7281 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2145_0 <=( _mesh_0_3_io_out_id_0) ^ ((fiEnable && (7282 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2146_0 <=( _mesh_1_3_io_out_id_0) ^ ((fiEnable && (7283 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2147_0 <=( _mesh_2_3_io_out_id_0) ^ ((fiEnable && (7284 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2148_0 <=( _mesh_3_3_io_out_id_0) ^ ((fiEnable && (7285 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2149_0 <=( _mesh_4_3_io_out_id_0) ^ ((fiEnable && (7286 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2150_0 <=( _mesh_5_3_io_out_id_0) ^ ((fiEnable && (7287 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2151_0 <=( _mesh_6_3_io_out_id_0) ^ ((fiEnable && (7288 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2152_0 <=( _mesh_7_3_io_out_id_0) ^ ((fiEnable && (7289 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2153_0 <=( _mesh_8_3_io_out_id_0) ^ ((fiEnable && (7290 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2154_0 <=( _mesh_9_3_io_out_id_0) ^ ((fiEnable && (7291 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2155_0 <=( _mesh_10_3_io_out_id_0) ^ ((fiEnable && (7292 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2156_0 <=( _mesh_11_3_io_out_id_0) ^ ((fiEnable && (7293 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2157_0 <=( _mesh_12_3_io_out_id_0) ^ ((fiEnable && (7294 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2158_0 <=( _mesh_13_3_io_out_id_0) ^ ((fiEnable && (7295 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2159_0 <=( _mesh_14_3_io_out_id_0) ^ ((fiEnable && (7296 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2160_0 <=( _mesh_15_3_io_out_id_0) ^ ((fiEnable && (7297 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2161_0 <=( _mesh_16_3_io_out_id_0) ^ ((fiEnable && (7298 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2162_0 <=( _mesh_17_3_io_out_id_0) ^ ((fiEnable && (7299 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2163_0 <=( _mesh_18_3_io_out_id_0) ^ ((fiEnable && (7300 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2164_0 <=( _mesh_19_3_io_out_id_0) ^ ((fiEnable && (7301 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2165_0 <=( _mesh_20_3_io_out_id_0) ^ ((fiEnable && (7302 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2166_0 <=( _mesh_21_3_io_out_id_0) ^ ((fiEnable && (7303 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2167_0 <=( _mesh_22_3_io_out_id_0) ^ ((fiEnable && (7304 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2168_0 <=( _mesh_23_3_io_out_id_0) ^ ((fiEnable && (7305 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2169_0 <=( _mesh_24_3_io_out_id_0) ^ ((fiEnable && (7306 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2170_0 <=( _mesh_25_3_io_out_id_0) ^ ((fiEnable && (7307 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2171_0 <=( _mesh_26_3_io_out_id_0) ^ ((fiEnable && (7308 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2172_0 <=( _mesh_27_3_io_out_id_0) ^ ((fiEnable && (7309 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2173_0 <=( _mesh_28_3_io_out_id_0) ^ ((fiEnable && (7310 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2174_0 <=( _mesh_29_3_io_out_id_0) ^ ((fiEnable && (7311 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2175_0 <=( _mesh_30_3_io_out_id_0) ^ ((fiEnable && (7312 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2176_0 <=( io_in_id_4_0) ^ ((fiEnable && (7313 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2177_0 <=( _mesh_0_4_io_out_id_0) ^ ((fiEnable && (7314 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2178_0 <=( _mesh_1_4_io_out_id_0) ^ ((fiEnable && (7315 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2179_0 <=( _mesh_2_4_io_out_id_0) ^ ((fiEnable && (7316 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2180_0 <=( _mesh_3_4_io_out_id_0) ^ ((fiEnable && (7317 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2181_0 <=( _mesh_4_4_io_out_id_0) ^ ((fiEnable && (7318 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2182_0 <=( _mesh_5_4_io_out_id_0) ^ ((fiEnable && (7319 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2183_0 <=( _mesh_6_4_io_out_id_0) ^ ((fiEnable && (7320 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2184_0 <=( _mesh_7_4_io_out_id_0) ^ ((fiEnable && (7321 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2185_0 <=( _mesh_8_4_io_out_id_0) ^ ((fiEnable && (7322 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2186_0 <=( _mesh_9_4_io_out_id_0) ^ ((fiEnable && (7323 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2187_0 <=( _mesh_10_4_io_out_id_0) ^ ((fiEnable && (7324 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2188_0 <=( _mesh_11_4_io_out_id_0) ^ ((fiEnable && (7325 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2189_0 <=( _mesh_12_4_io_out_id_0) ^ ((fiEnable && (7326 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2190_0 <=( _mesh_13_4_io_out_id_0) ^ ((fiEnable && (7327 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2191_0 <=( _mesh_14_4_io_out_id_0) ^ ((fiEnable && (7328 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2192_0 <=( _mesh_15_4_io_out_id_0) ^ ((fiEnable && (7329 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2193_0 <=( _mesh_16_4_io_out_id_0) ^ ((fiEnable && (7330 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2194_0 <=( _mesh_17_4_io_out_id_0) ^ ((fiEnable && (7331 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2195_0 <=( _mesh_18_4_io_out_id_0) ^ ((fiEnable && (7332 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2196_0 <=( _mesh_19_4_io_out_id_0) ^ ((fiEnable && (7333 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2197_0 <=( _mesh_20_4_io_out_id_0) ^ ((fiEnable && (7334 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2198_0 <=( _mesh_21_4_io_out_id_0) ^ ((fiEnable && (7335 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2199_0 <=( _mesh_22_4_io_out_id_0) ^ ((fiEnable && (7336 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2200_0 <=( _mesh_23_4_io_out_id_0) ^ ((fiEnable && (7337 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2201_0 <=( _mesh_24_4_io_out_id_0) ^ ((fiEnable && (7338 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2202_0 <=( _mesh_25_4_io_out_id_0) ^ ((fiEnable && (7339 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2203_0 <=( _mesh_26_4_io_out_id_0) ^ ((fiEnable && (7340 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2204_0 <=( _mesh_27_4_io_out_id_0) ^ ((fiEnable && (7341 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2205_0 <=( _mesh_28_4_io_out_id_0) ^ ((fiEnable && (7342 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2206_0 <=( _mesh_29_4_io_out_id_0) ^ ((fiEnable && (7343 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2207_0 <=( _mesh_30_4_io_out_id_0) ^ ((fiEnable && (7344 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2208_0 <=( io_in_id_5_0) ^ ((fiEnable && (7345 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2209_0 <=( _mesh_0_5_io_out_id_0) ^ ((fiEnable && (7346 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2210_0 <=( _mesh_1_5_io_out_id_0) ^ ((fiEnable && (7347 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2211_0 <=( _mesh_2_5_io_out_id_0) ^ ((fiEnable && (7348 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2212_0 <=( _mesh_3_5_io_out_id_0) ^ ((fiEnable && (7349 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2213_0 <=( _mesh_4_5_io_out_id_0) ^ ((fiEnable && (7350 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2214_0 <=( _mesh_5_5_io_out_id_0) ^ ((fiEnable && (7351 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2215_0 <=( _mesh_6_5_io_out_id_0) ^ ((fiEnable && (7352 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2216_0 <=( _mesh_7_5_io_out_id_0) ^ ((fiEnable && (7353 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2217_0 <=( _mesh_8_5_io_out_id_0) ^ ((fiEnable && (7354 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2218_0 <=( _mesh_9_5_io_out_id_0) ^ ((fiEnable && (7355 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2219_0 <=( _mesh_10_5_io_out_id_0) ^ ((fiEnable && (7356 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2220_0 <=( _mesh_11_5_io_out_id_0) ^ ((fiEnable && (7357 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2221_0 <=( _mesh_12_5_io_out_id_0) ^ ((fiEnable && (7358 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2222_0 <=( _mesh_13_5_io_out_id_0) ^ ((fiEnable && (7359 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2223_0 <=( _mesh_14_5_io_out_id_0) ^ ((fiEnable && (7360 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2224_0 <=( _mesh_15_5_io_out_id_0) ^ ((fiEnable && (7361 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2225_0 <=( _mesh_16_5_io_out_id_0) ^ ((fiEnable && (7362 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2226_0 <=( _mesh_17_5_io_out_id_0) ^ ((fiEnable && (7363 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2227_0 <=( _mesh_18_5_io_out_id_0) ^ ((fiEnable && (7364 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2228_0 <=( _mesh_19_5_io_out_id_0) ^ ((fiEnable && (7365 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2229_0 <=( _mesh_20_5_io_out_id_0) ^ ((fiEnable && (7366 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2230_0 <=( _mesh_21_5_io_out_id_0) ^ ((fiEnable && (7367 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2231_0 <=( _mesh_22_5_io_out_id_0) ^ ((fiEnable && (7368 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2232_0 <=( _mesh_23_5_io_out_id_0) ^ ((fiEnable && (7369 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2233_0 <=( _mesh_24_5_io_out_id_0) ^ ((fiEnable && (7370 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2234_0 <=( _mesh_25_5_io_out_id_0) ^ ((fiEnable && (7371 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2235_0 <=( _mesh_26_5_io_out_id_0) ^ ((fiEnable && (7372 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2236_0 <=( _mesh_27_5_io_out_id_0) ^ ((fiEnable && (7373 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2237_0 <=( _mesh_28_5_io_out_id_0) ^ ((fiEnable && (7374 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2238_0 <=( _mesh_29_5_io_out_id_0) ^ ((fiEnable && (7375 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2239_0 <=( _mesh_30_5_io_out_id_0) ^ ((fiEnable && (7376 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2240_0 <=( io_in_id_6_0) ^ ((fiEnable && (7377 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2241_0 <=( _mesh_0_6_io_out_id_0) ^ ((fiEnable && (7378 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2242_0 <=( _mesh_1_6_io_out_id_0) ^ ((fiEnable && (7379 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2243_0 <=( _mesh_2_6_io_out_id_0) ^ ((fiEnable && (7380 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2244_0 <=( _mesh_3_6_io_out_id_0) ^ ((fiEnable && (7381 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2245_0 <=( _mesh_4_6_io_out_id_0) ^ ((fiEnable && (7382 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2246_0 <=( _mesh_5_6_io_out_id_0) ^ ((fiEnable && (7383 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2247_0 <=( _mesh_6_6_io_out_id_0) ^ ((fiEnable && (7384 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2248_0 <=( _mesh_7_6_io_out_id_0) ^ ((fiEnable && (7385 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2249_0 <=( _mesh_8_6_io_out_id_0) ^ ((fiEnable && (7386 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2250_0 <=( _mesh_9_6_io_out_id_0) ^ ((fiEnable && (7387 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2251_0 <=( _mesh_10_6_io_out_id_0) ^ ((fiEnable && (7388 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2252_0 <=( _mesh_11_6_io_out_id_0) ^ ((fiEnable && (7389 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2253_0 <=( _mesh_12_6_io_out_id_0) ^ ((fiEnable && (7390 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2254_0 <=( _mesh_13_6_io_out_id_0) ^ ((fiEnable && (7391 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2255_0 <=( _mesh_14_6_io_out_id_0) ^ ((fiEnable && (7392 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2256_0 <=( _mesh_15_6_io_out_id_0) ^ ((fiEnable && (7393 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2257_0 <=( _mesh_16_6_io_out_id_0) ^ ((fiEnable && (7394 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2258_0 <=( _mesh_17_6_io_out_id_0) ^ ((fiEnable && (7395 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2259_0 <=( _mesh_18_6_io_out_id_0) ^ ((fiEnable && (7396 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2260_0 <=( _mesh_19_6_io_out_id_0) ^ ((fiEnable && (7397 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2261_0 <=( _mesh_20_6_io_out_id_0) ^ ((fiEnable && (7398 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2262_0 <=( _mesh_21_6_io_out_id_0) ^ ((fiEnable && (7399 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2263_0 <=( _mesh_22_6_io_out_id_0) ^ ((fiEnable && (7400 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2264_0 <=( _mesh_23_6_io_out_id_0) ^ ((fiEnable && (7401 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2265_0 <=( _mesh_24_6_io_out_id_0) ^ ((fiEnable && (7402 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2266_0 <=( _mesh_25_6_io_out_id_0) ^ ((fiEnable && (7403 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2267_0 <=( _mesh_26_6_io_out_id_0) ^ ((fiEnable && (7404 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2268_0 <=( _mesh_27_6_io_out_id_0) ^ ((fiEnable && (7405 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2269_0 <=( _mesh_28_6_io_out_id_0) ^ ((fiEnable && (7406 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2270_0 <=( _mesh_29_6_io_out_id_0) ^ ((fiEnable && (7407 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2271_0 <=( _mesh_30_6_io_out_id_0) ^ ((fiEnable && (7408 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2272_0 <=( io_in_id_7_0) ^ ((fiEnable && (7409 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2273_0 <=( _mesh_0_7_io_out_id_0) ^ ((fiEnable && (7410 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2274_0 <=( _mesh_1_7_io_out_id_0) ^ ((fiEnable && (7411 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2275_0 <=( _mesh_2_7_io_out_id_0) ^ ((fiEnable && (7412 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2276_0 <=( _mesh_3_7_io_out_id_0) ^ ((fiEnable && (7413 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2277_0 <=( _mesh_4_7_io_out_id_0) ^ ((fiEnable && (7414 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2278_0 <=( _mesh_5_7_io_out_id_0) ^ ((fiEnable && (7415 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2279_0 <=( _mesh_6_7_io_out_id_0) ^ ((fiEnable && (7416 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2280_0 <=( _mesh_7_7_io_out_id_0) ^ ((fiEnable && (7417 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2281_0 <=( _mesh_8_7_io_out_id_0) ^ ((fiEnable && (7418 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2282_0 <=( _mesh_9_7_io_out_id_0) ^ ((fiEnable && (7419 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2283_0 <=( _mesh_10_7_io_out_id_0) ^ ((fiEnable && (7420 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2284_0 <=( _mesh_11_7_io_out_id_0) ^ ((fiEnable && (7421 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2285_0 <=( _mesh_12_7_io_out_id_0) ^ ((fiEnable && (7422 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2286_0 <=( _mesh_13_7_io_out_id_0) ^ ((fiEnable && (7423 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2287_0 <=( _mesh_14_7_io_out_id_0) ^ ((fiEnable && (7424 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2288_0 <=( _mesh_15_7_io_out_id_0) ^ ((fiEnable && (7425 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2289_0 <=( _mesh_16_7_io_out_id_0) ^ ((fiEnable && (7426 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2290_0 <=( _mesh_17_7_io_out_id_0) ^ ((fiEnable && (7427 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2291_0 <=( _mesh_18_7_io_out_id_0) ^ ((fiEnable && (7428 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2292_0 <=( _mesh_19_7_io_out_id_0) ^ ((fiEnable && (7429 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2293_0 <=( _mesh_20_7_io_out_id_0) ^ ((fiEnable && (7430 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2294_0 <=( _mesh_21_7_io_out_id_0) ^ ((fiEnable && (7431 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2295_0 <=( _mesh_22_7_io_out_id_0) ^ ((fiEnable && (7432 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2296_0 <=( _mesh_23_7_io_out_id_0) ^ ((fiEnable && (7433 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2297_0 <=( _mesh_24_7_io_out_id_0) ^ ((fiEnable && (7434 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2298_0 <=( _mesh_25_7_io_out_id_0) ^ ((fiEnable && (7435 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2299_0 <=( _mesh_26_7_io_out_id_0) ^ ((fiEnable && (7436 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2300_0 <=( _mesh_27_7_io_out_id_0) ^ ((fiEnable && (7437 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2301_0 <=( _mesh_28_7_io_out_id_0) ^ ((fiEnable && (7438 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2302_0 <=( _mesh_29_7_io_out_id_0) ^ ((fiEnable && (7439 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2303_0 <=( _mesh_30_7_io_out_id_0) ^ ((fiEnable && (7440 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2304_0 <=( io_in_id_8_0) ^ ((fiEnable && (7441 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2305_0 <=( _mesh_0_8_io_out_id_0) ^ ((fiEnable && (7442 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2306_0 <=( _mesh_1_8_io_out_id_0) ^ ((fiEnable && (7443 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2307_0 <=( _mesh_2_8_io_out_id_0) ^ ((fiEnable && (7444 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2308_0 <=( _mesh_3_8_io_out_id_0) ^ ((fiEnable && (7445 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2309_0 <=( _mesh_4_8_io_out_id_0) ^ ((fiEnable && (7446 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2310_0 <=( _mesh_5_8_io_out_id_0) ^ ((fiEnable && (7447 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2311_0 <=( _mesh_6_8_io_out_id_0) ^ ((fiEnable && (7448 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2312_0 <=( _mesh_7_8_io_out_id_0) ^ ((fiEnable && (7449 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2313_0 <=( _mesh_8_8_io_out_id_0) ^ ((fiEnable && (7450 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2314_0 <=( _mesh_9_8_io_out_id_0) ^ ((fiEnable && (7451 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2315_0 <=( _mesh_10_8_io_out_id_0) ^ ((fiEnable && (7452 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2316_0 <=( _mesh_11_8_io_out_id_0) ^ ((fiEnable && (7453 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2317_0 <=( _mesh_12_8_io_out_id_0) ^ ((fiEnable && (7454 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2318_0 <=( _mesh_13_8_io_out_id_0) ^ ((fiEnable && (7455 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2319_0 <=( _mesh_14_8_io_out_id_0) ^ ((fiEnable && (7456 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2320_0 <=( _mesh_15_8_io_out_id_0) ^ ((fiEnable && (7457 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2321_0 <=( _mesh_16_8_io_out_id_0) ^ ((fiEnable && (7458 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2322_0 <=( _mesh_17_8_io_out_id_0) ^ ((fiEnable && (7459 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2323_0 <=( _mesh_18_8_io_out_id_0) ^ ((fiEnable && (7460 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2324_0 <=( _mesh_19_8_io_out_id_0) ^ ((fiEnable && (7461 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2325_0 <=( _mesh_20_8_io_out_id_0) ^ ((fiEnable && (7462 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2326_0 <=( _mesh_21_8_io_out_id_0) ^ ((fiEnable && (7463 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2327_0 <=( _mesh_22_8_io_out_id_0) ^ ((fiEnable && (7464 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2328_0 <=( _mesh_23_8_io_out_id_0) ^ ((fiEnable && (7465 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2329_0 <=( _mesh_24_8_io_out_id_0) ^ ((fiEnable && (7466 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2330_0 <=( _mesh_25_8_io_out_id_0) ^ ((fiEnable && (7467 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2331_0 <=( _mesh_26_8_io_out_id_0) ^ ((fiEnable && (7468 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2332_0 <=( _mesh_27_8_io_out_id_0) ^ ((fiEnable && (7469 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2333_0 <=( _mesh_28_8_io_out_id_0) ^ ((fiEnable && (7470 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2334_0 <=( _mesh_29_8_io_out_id_0) ^ ((fiEnable && (7471 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2335_0 <=( _mesh_30_8_io_out_id_0) ^ ((fiEnable && (7472 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2336_0 <=( io_in_id_9_0) ^ ((fiEnable && (7473 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2337_0 <=( _mesh_0_9_io_out_id_0) ^ ((fiEnable && (7474 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2338_0 <=( _mesh_1_9_io_out_id_0) ^ ((fiEnable && (7475 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2339_0 <=( _mesh_2_9_io_out_id_0) ^ ((fiEnable && (7476 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2340_0 <=( _mesh_3_9_io_out_id_0) ^ ((fiEnable && (7477 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2341_0 <=( _mesh_4_9_io_out_id_0) ^ ((fiEnable && (7478 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2342_0 <=( _mesh_5_9_io_out_id_0) ^ ((fiEnable && (7479 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2343_0 <=( _mesh_6_9_io_out_id_0) ^ ((fiEnable && (7480 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2344_0 <=( _mesh_7_9_io_out_id_0) ^ ((fiEnable && (7481 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2345_0 <=( _mesh_8_9_io_out_id_0) ^ ((fiEnable && (7482 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2346_0 <=( _mesh_9_9_io_out_id_0) ^ ((fiEnable && (7483 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2347_0 <=( _mesh_10_9_io_out_id_0) ^ ((fiEnable && (7484 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2348_0 <=( _mesh_11_9_io_out_id_0) ^ ((fiEnable && (7485 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2349_0 <=( _mesh_12_9_io_out_id_0) ^ ((fiEnable && (7486 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2350_0 <=( _mesh_13_9_io_out_id_0) ^ ((fiEnable && (7487 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2351_0 <=( _mesh_14_9_io_out_id_0) ^ ((fiEnable && (7488 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2352_0 <=( _mesh_15_9_io_out_id_0) ^ ((fiEnable && (7489 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2353_0 <=( _mesh_16_9_io_out_id_0) ^ ((fiEnable && (7490 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2354_0 <=( _mesh_17_9_io_out_id_0) ^ ((fiEnable && (7491 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2355_0 <=( _mesh_18_9_io_out_id_0) ^ ((fiEnable && (7492 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2356_0 <=( _mesh_19_9_io_out_id_0) ^ ((fiEnable && (7493 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2357_0 <=( _mesh_20_9_io_out_id_0) ^ ((fiEnable && (7494 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2358_0 <=( _mesh_21_9_io_out_id_0) ^ ((fiEnable && (7495 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2359_0 <=( _mesh_22_9_io_out_id_0) ^ ((fiEnable && (7496 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2360_0 <=( _mesh_23_9_io_out_id_0) ^ ((fiEnable && (7497 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2361_0 <=( _mesh_24_9_io_out_id_0) ^ ((fiEnable && (7498 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2362_0 <=( _mesh_25_9_io_out_id_0) ^ ((fiEnable && (7499 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2363_0 <=( _mesh_26_9_io_out_id_0) ^ ((fiEnable && (7500 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2364_0 <=( _mesh_27_9_io_out_id_0) ^ ((fiEnable && (7501 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2365_0 <=( _mesh_28_9_io_out_id_0) ^ ((fiEnable && (7502 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2366_0 <=( _mesh_29_9_io_out_id_0) ^ ((fiEnable && (7503 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2367_0 <=( _mesh_30_9_io_out_id_0) ^ ((fiEnable && (7504 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2368_0 <=( io_in_id_10_0) ^ ((fiEnable && (7505 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2369_0 <=( _mesh_0_10_io_out_id_0) ^ ((fiEnable && (7506 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2370_0 <=( _mesh_1_10_io_out_id_0) ^ ((fiEnable && (7507 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2371_0 <=( _mesh_2_10_io_out_id_0) ^ ((fiEnable && (7508 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2372_0 <=( _mesh_3_10_io_out_id_0) ^ ((fiEnable && (7509 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2373_0 <=( _mesh_4_10_io_out_id_0) ^ ((fiEnable && (7510 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2374_0 <=( _mesh_5_10_io_out_id_0) ^ ((fiEnable && (7511 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2375_0 <=( _mesh_6_10_io_out_id_0) ^ ((fiEnable && (7512 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2376_0 <=( _mesh_7_10_io_out_id_0) ^ ((fiEnable && (7513 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2377_0 <=( _mesh_8_10_io_out_id_0) ^ ((fiEnable && (7514 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2378_0 <=( _mesh_9_10_io_out_id_0) ^ ((fiEnable && (7515 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2379_0 <=( _mesh_10_10_io_out_id_0) ^ ((fiEnable && (7516 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2380_0 <=( _mesh_11_10_io_out_id_0) ^ ((fiEnable && (7517 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2381_0 <=( _mesh_12_10_io_out_id_0) ^ ((fiEnable && (7518 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2382_0 <=( _mesh_13_10_io_out_id_0) ^ ((fiEnable && (7519 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2383_0 <=( _mesh_14_10_io_out_id_0) ^ ((fiEnable && (7520 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2384_0 <=( _mesh_15_10_io_out_id_0) ^ ((fiEnable && (7521 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2385_0 <=( _mesh_16_10_io_out_id_0) ^ ((fiEnable && (7522 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2386_0 <=( _mesh_17_10_io_out_id_0) ^ ((fiEnable && (7523 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2387_0 <=( _mesh_18_10_io_out_id_0) ^ ((fiEnable && (7524 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2388_0 <=( _mesh_19_10_io_out_id_0) ^ ((fiEnable && (7525 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2389_0 <=( _mesh_20_10_io_out_id_0) ^ ((fiEnable && (7526 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2390_0 <=( _mesh_21_10_io_out_id_0) ^ ((fiEnable && (7527 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2391_0 <=( _mesh_22_10_io_out_id_0) ^ ((fiEnable && (7528 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2392_0 <=( _mesh_23_10_io_out_id_0) ^ ((fiEnable && (7529 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2393_0 <=( _mesh_24_10_io_out_id_0) ^ ((fiEnable && (7530 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2394_0 <=( _mesh_25_10_io_out_id_0) ^ ((fiEnable && (7531 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2395_0 <=( _mesh_26_10_io_out_id_0) ^ ((fiEnable && (7532 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2396_0 <=( _mesh_27_10_io_out_id_0) ^ ((fiEnable && (7533 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2397_0 <=( _mesh_28_10_io_out_id_0) ^ ((fiEnable && (7534 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2398_0 <=( _mesh_29_10_io_out_id_0) ^ ((fiEnable && (7535 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2399_0 <=( _mesh_30_10_io_out_id_0) ^ ((fiEnable && (7536 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2400_0 <=( io_in_id_11_0) ^ ((fiEnable && (7537 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2401_0 <=( _mesh_0_11_io_out_id_0) ^ ((fiEnable && (7538 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2402_0 <=( _mesh_1_11_io_out_id_0) ^ ((fiEnable && (7539 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2403_0 <=( _mesh_2_11_io_out_id_0) ^ ((fiEnable && (7540 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2404_0 <=( _mesh_3_11_io_out_id_0) ^ ((fiEnable && (7541 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2405_0 <=( _mesh_4_11_io_out_id_0) ^ ((fiEnable && (7542 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2406_0 <=( _mesh_5_11_io_out_id_0) ^ ((fiEnable && (7543 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2407_0 <=( _mesh_6_11_io_out_id_0) ^ ((fiEnable && (7544 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2408_0 <=( _mesh_7_11_io_out_id_0) ^ ((fiEnable && (7545 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2409_0 <=( _mesh_8_11_io_out_id_0) ^ ((fiEnable && (7546 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2410_0 <=( _mesh_9_11_io_out_id_0) ^ ((fiEnable && (7547 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2411_0 <=( _mesh_10_11_io_out_id_0) ^ ((fiEnable && (7548 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2412_0 <=( _mesh_11_11_io_out_id_0) ^ ((fiEnable && (7549 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2413_0 <=( _mesh_12_11_io_out_id_0) ^ ((fiEnable && (7550 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2414_0 <=( _mesh_13_11_io_out_id_0) ^ ((fiEnable && (7551 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2415_0 <=( _mesh_14_11_io_out_id_0) ^ ((fiEnable && (7552 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2416_0 <=( _mesh_15_11_io_out_id_0) ^ ((fiEnable && (7553 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2417_0 <=( _mesh_16_11_io_out_id_0) ^ ((fiEnable && (7554 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2418_0 <=( _mesh_17_11_io_out_id_0) ^ ((fiEnable && (7555 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2419_0 <=( _mesh_18_11_io_out_id_0) ^ ((fiEnable && (7556 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2420_0 <=( _mesh_19_11_io_out_id_0) ^ ((fiEnable && (7557 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2421_0 <=( _mesh_20_11_io_out_id_0) ^ ((fiEnable && (7558 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2422_0 <=( _mesh_21_11_io_out_id_0) ^ ((fiEnable && (7559 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2423_0 <=( _mesh_22_11_io_out_id_0) ^ ((fiEnable && (7560 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2424_0 <=( _mesh_23_11_io_out_id_0) ^ ((fiEnable && (7561 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2425_0 <=( _mesh_24_11_io_out_id_0) ^ ((fiEnable && (7562 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2426_0 <=( _mesh_25_11_io_out_id_0) ^ ((fiEnable && (7563 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2427_0 <=( _mesh_26_11_io_out_id_0) ^ ((fiEnable && (7564 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2428_0 <=( _mesh_27_11_io_out_id_0) ^ ((fiEnable && (7565 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2429_0 <=( _mesh_28_11_io_out_id_0) ^ ((fiEnable && (7566 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2430_0 <=( _mesh_29_11_io_out_id_0) ^ ((fiEnable && (7567 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2431_0 <=( _mesh_30_11_io_out_id_0) ^ ((fiEnable && (7568 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2432_0 <=( io_in_id_12_0) ^ ((fiEnable && (7569 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2433_0 <=( _mesh_0_12_io_out_id_0) ^ ((fiEnable && (7570 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2434_0 <=( _mesh_1_12_io_out_id_0) ^ ((fiEnable && (7571 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2435_0 <=( _mesh_2_12_io_out_id_0) ^ ((fiEnable && (7572 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2436_0 <=( _mesh_3_12_io_out_id_0) ^ ((fiEnable && (7573 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2437_0 <=( _mesh_4_12_io_out_id_0) ^ ((fiEnable && (7574 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2438_0 <=( _mesh_5_12_io_out_id_0) ^ ((fiEnable && (7575 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2439_0 <=( _mesh_6_12_io_out_id_0) ^ ((fiEnable && (7576 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2440_0 <=( _mesh_7_12_io_out_id_0) ^ ((fiEnable && (7577 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2441_0 <=( _mesh_8_12_io_out_id_0) ^ ((fiEnable && (7578 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2442_0 <=( _mesh_9_12_io_out_id_0) ^ ((fiEnable && (7579 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2443_0 <=( _mesh_10_12_io_out_id_0) ^ ((fiEnable && (7580 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2444_0 <=( _mesh_11_12_io_out_id_0) ^ ((fiEnable && (7581 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2445_0 <=( _mesh_12_12_io_out_id_0) ^ ((fiEnable && (7582 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2446_0 <=( _mesh_13_12_io_out_id_0) ^ ((fiEnable && (7583 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2447_0 <=( _mesh_14_12_io_out_id_0) ^ ((fiEnable && (7584 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2448_0 <=( _mesh_15_12_io_out_id_0) ^ ((fiEnable && (7585 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2449_0 <=( _mesh_16_12_io_out_id_0) ^ ((fiEnable && (7586 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2450_0 <=( _mesh_17_12_io_out_id_0) ^ ((fiEnable && (7587 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2451_0 <=( _mesh_18_12_io_out_id_0) ^ ((fiEnable && (7588 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2452_0 <=( _mesh_19_12_io_out_id_0) ^ ((fiEnable && (7589 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2453_0 <=( _mesh_20_12_io_out_id_0) ^ ((fiEnable && (7590 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2454_0 <=( _mesh_21_12_io_out_id_0) ^ ((fiEnable && (7591 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2455_0 <=( _mesh_22_12_io_out_id_0) ^ ((fiEnable && (7592 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2456_0 <=( _mesh_23_12_io_out_id_0) ^ ((fiEnable && (7593 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2457_0 <=( _mesh_24_12_io_out_id_0) ^ ((fiEnable && (7594 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2458_0 <=( _mesh_25_12_io_out_id_0) ^ ((fiEnable && (7595 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2459_0 <=( _mesh_26_12_io_out_id_0) ^ ((fiEnable && (7596 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2460_0 <=( _mesh_27_12_io_out_id_0) ^ ((fiEnable && (7597 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2461_0 <=( _mesh_28_12_io_out_id_0) ^ ((fiEnable && (7598 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2462_0 <=( _mesh_29_12_io_out_id_0) ^ ((fiEnable && (7599 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2463_0 <=( _mesh_30_12_io_out_id_0) ^ ((fiEnable && (7600 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2464_0 <=( io_in_id_13_0) ^ ((fiEnable && (7601 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2465_0 <=( _mesh_0_13_io_out_id_0) ^ ((fiEnable && (7602 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2466_0 <=( _mesh_1_13_io_out_id_0) ^ ((fiEnable && (7603 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2467_0 <=( _mesh_2_13_io_out_id_0) ^ ((fiEnable && (7604 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2468_0 <=( _mesh_3_13_io_out_id_0) ^ ((fiEnable && (7605 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2469_0 <=( _mesh_4_13_io_out_id_0) ^ ((fiEnable && (7606 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2470_0 <=( _mesh_5_13_io_out_id_0) ^ ((fiEnable && (7607 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2471_0 <=( _mesh_6_13_io_out_id_0) ^ ((fiEnable && (7608 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2472_0 <=( _mesh_7_13_io_out_id_0) ^ ((fiEnable && (7609 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2473_0 <=( _mesh_8_13_io_out_id_0) ^ ((fiEnable && (7610 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2474_0 <=( _mesh_9_13_io_out_id_0) ^ ((fiEnable && (7611 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2475_0 <=( _mesh_10_13_io_out_id_0) ^ ((fiEnable && (7612 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2476_0 <=( _mesh_11_13_io_out_id_0) ^ ((fiEnable && (7613 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2477_0 <=( _mesh_12_13_io_out_id_0) ^ ((fiEnable && (7614 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2478_0 <=( _mesh_13_13_io_out_id_0) ^ ((fiEnable && (7615 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2479_0 <=( _mesh_14_13_io_out_id_0) ^ ((fiEnable && (7616 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2480_0 <=( _mesh_15_13_io_out_id_0) ^ ((fiEnable && (7617 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2481_0 <=( _mesh_16_13_io_out_id_0) ^ ((fiEnable && (7618 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2482_0 <=( _mesh_17_13_io_out_id_0) ^ ((fiEnable && (7619 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2483_0 <=( _mesh_18_13_io_out_id_0) ^ ((fiEnable && (7620 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2484_0 <=( _mesh_19_13_io_out_id_0) ^ ((fiEnable && (7621 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2485_0 <=( _mesh_20_13_io_out_id_0) ^ ((fiEnable && (7622 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2486_0 <=( _mesh_21_13_io_out_id_0) ^ ((fiEnable && (7623 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2487_0 <=( _mesh_22_13_io_out_id_0) ^ ((fiEnable && (7624 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2488_0 <=( _mesh_23_13_io_out_id_0) ^ ((fiEnable && (7625 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2489_0 <=( _mesh_24_13_io_out_id_0) ^ ((fiEnable && (7626 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2490_0 <=( _mesh_25_13_io_out_id_0) ^ ((fiEnable && (7627 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2491_0 <=( _mesh_26_13_io_out_id_0) ^ ((fiEnable && (7628 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2492_0 <=( _mesh_27_13_io_out_id_0) ^ ((fiEnable && (7629 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2493_0 <=( _mesh_28_13_io_out_id_0) ^ ((fiEnable && (7630 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2494_0 <=( _mesh_29_13_io_out_id_0) ^ ((fiEnable && (7631 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2495_0 <=( _mesh_30_13_io_out_id_0) ^ ((fiEnable && (7632 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2496_0 <=( io_in_id_14_0) ^ ((fiEnable && (7633 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2497_0 <=( _mesh_0_14_io_out_id_0) ^ ((fiEnable && (7634 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2498_0 <=( _mesh_1_14_io_out_id_0) ^ ((fiEnable && (7635 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2499_0 <=( _mesh_2_14_io_out_id_0) ^ ((fiEnable && (7636 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2500_0 <=( _mesh_3_14_io_out_id_0) ^ ((fiEnable && (7637 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2501_0 <=( _mesh_4_14_io_out_id_0) ^ ((fiEnable && (7638 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2502_0 <=( _mesh_5_14_io_out_id_0) ^ ((fiEnable && (7639 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2503_0 <=( _mesh_6_14_io_out_id_0) ^ ((fiEnable && (7640 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2504_0 <=( _mesh_7_14_io_out_id_0) ^ ((fiEnable && (7641 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2505_0 <=( _mesh_8_14_io_out_id_0) ^ ((fiEnable && (7642 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2506_0 <=( _mesh_9_14_io_out_id_0) ^ ((fiEnable && (7643 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2507_0 <=( _mesh_10_14_io_out_id_0) ^ ((fiEnable && (7644 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2508_0 <=( _mesh_11_14_io_out_id_0) ^ ((fiEnable && (7645 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2509_0 <=( _mesh_12_14_io_out_id_0) ^ ((fiEnable && (7646 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2510_0 <=( _mesh_13_14_io_out_id_0) ^ ((fiEnable && (7647 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2511_0 <=( _mesh_14_14_io_out_id_0) ^ ((fiEnable && (7648 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2512_0 <=( _mesh_15_14_io_out_id_0) ^ ((fiEnable && (7649 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2513_0 <=( _mesh_16_14_io_out_id_0) ^ ((fiEnable && (7650 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2514_0 <=( _mesh_17_14_io_out_id_0) ^ ((fiEnable && (7651 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2515_0 <=( _mesh_18_14_io_out_id_0) ^ ((fiEnable && (7652 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2516_0 <=( _mesh_19_14_io_out_id_0) ^ ((fiEnable && (7653 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2517_0 <=( _mesh_20_14_io_out_id_0) ^ ((fiEnable && (7654 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2518_0 <=( _mesh_21_14_io_out_id_0) ^ ((fiEnable && (7655 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2519_0 <=( _mesh_22_14_io_out_id_0) ^ ((fiEnable && (7656 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2520_0 <=( _mesh_23_14_io_out_id_0) ^ ((fiEnable && (7657 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2521_0 <=( _mesh_24_14_io_out_id_0) ^ ((fiEnable && (7658 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2522_0 <=( _mesh_25_14_io_out_id_0) ^ ((fiEnable && (7659 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2523_0 <=( _mesh_26_14_io_out_id_0) ^ ((fiEnable && (7660 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2524_0 <=( _mesh_27_14_io_out_id_0) ^ ((fiEnable && (7661 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2525_0 <=( _mesh_28_14_io_out_id_0) ^ ((fiEnable && (7662 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2526_0 <=( _mesh_29_14_io_out_id_0) ^ ((fiEnable && (7663 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2527_0 <=( _mesh_30_14_io_out_id_0) ^ ((fiEnable && (7664 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2528_0 <=( io_in_id_15_0) ^ ((fiEnable && (7665 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2529_0 <=( _mesh_0_15_io_out_id_0) ^ ((fiEnable && (7666 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2530_0 <=( _mesh_1_15_io_out_id_0) ^ ((fiEnable && (7667 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2531_0 <=( _mesh_2_15_io_out_id_0) ^ ((fiEnable && (7668 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2532_0 <=( _mesh_3_15_io_out_id_0) ^ ((fiEnable && (7669 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2533_0 <=( _mesh_4_15_io_out_id_0) ^ ((fiEnable && (7670 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2534_0 <=( _mesh_5_15_io_out_id_0) ^ ((fiEnable && (7671 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2535_0 <=( _mesh_6_15_io_out_id_0) ^ ((fiEnable && (7672 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2536_0 <=( _mesh_7_15_io_out_id_0) ^ ((fiEnable && (7673 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2537_0 <=( _mesh_8_15_io_out_id_0) ^ ((fiEnable && (7674 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2538_0 <=( _mesh_9_15_io_out_id_0) ^ ((fiEnable && (7675 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2539_0 <=( _mesh_10_15_io_out_id_0) ^ ((fiEnable && (7676 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2540_0 <=( _mesh_11_15_io_out_id_0) ^ ((fiEnable && (7677 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2541_0 <=( _mesh_12_15_io_out_id_0) ^ ((fiEnable && (7678 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2542_0 <=( _mesh_13_15_io_out_id_0) ^ ((fiEnable && (7679 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2543_0 <=( _mesh_14_15_io_out_id_0) ^ ((fiEnable && (7680 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2544_0 <=( _mesh_15_15_io_out_id_0) ^ ((fiEnable && (7681 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2545_0 <=( _mesh_16_15_io_out_id_0) ^ ((fiEnable && (7682 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2546_0 <=( _mesh_17_15_io_out_id_0) ^ ((fiEnable && (7683 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2547_0 <=( _mesh_18_15_io_out_id_0) ^ ((fiEnable && (7684 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2548_0 <=( _mesh_19_15_io_out_id_0) ^ ((fiEnable && (7685 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2549_0 <=( _mesh_20_15_io_out_id_0) ^ ((fiEnable && (7686 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2550_0 <=( _mesh_21_15_io_out_id_0) ^ ((fiEnable && (7687 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2551_0 <=( _mesh_22_15_io_out_id_0) ^ ((fiEnable && (7688 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2552_0 <=( _mesh_23_15_io_out_id_0) ^ ((fiEnable && (7689 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2553_0 <=( _mesh_24_15_io_out_id_0) ^ ((fiEnable && (7690 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2554_0 <=( _mesh_25_15_io_out_id_0) ^ ((fiEnable && (7691 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2555_0 <=( _mesh_26_15_io_out_id_0) ^ ((fiEnable && (7692 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2556_0 <=( _mesh_27_15_io_out_id_0) ^ ((fiEnable && (7693 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2557_0 <=( _mesh_28_15_io_out_id_0) ^ ((fiEnable && (7694 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2558_0 <=( _mesh_29_15_io_out_id_0) ^ ((fiEnable && (7695 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2559_0 <=( _mesh_30_15_io_out_id_0) ^ ((fiEnable && (7696 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2560_0 <=( io_in_id_16_0) ^ ((fiEnable && (7697 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2561_0 <=( _mesh_0_16_io_out_id_0) ^ ((fiEnable && (7698 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2562_0 <=( _mesh_1_16_io_out_id_0) ^ ((fiEnable && (7699 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2563_0 <=( _mesh_2_16_io_out_id_0) ^ ((fiEnable && (7700 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2564_0 <=( _mesh_3_16_io_out_id_0) ^ ((fiEnable && (7701 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2565_0 <=( _mesh_4_16_io_out_id_0) ^ ((fiEnable && (7702 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2566_0 <=( _mesh_5_16_io_out_id_0) ^ ((fiEnable && (7703 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2567_0 <=( _mesh_6_16_io_out_id_0) ^ ((fiEnable && (7704 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2568_0 <=( _mesh_7_16_io_out_id_0) ^ ((fiEnable && (7705 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2569_0 <=( _mesh_8_16_io_out_id_0) ^ ((fiEnable && (7706 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2570_0 <=( _mesh_9_16_io_out_id_0) ^ ((fiEnable && (7707 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2571_0 <=( _mesh_10_16_io_out_id_0) ^ ((fiEnable && (7708 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2572_0 <=( _mesh_11_16_io_out_id_0) ^ ((fiEnable && (7709 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2573_0 <=( _mesh_12_16_io_out_id_0) ^ ((fiEnable && (7710 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2574_0 <=( _mesh_13_16_io_out_id_0) ^ ((fiEnable && (7711 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2575_0 <=( _mesh_14_16_io_out_id_0) ^ ((fiEnable && (7712 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2576_0 <=( _mesh_15_16_io_out_id_0) ^ ((fiEnable && (7713 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2577_0 <=( _mesh_16_16_io_out_id_0) ^ ((fiEnable && (7714 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2578_0 <=( _mesh_17_16_io_out_id_0) ^ ((fiEnable && (7715 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2579_0 <=( _mesh_18_16_io_out_id_0) ^ ((fiEnable && (7716 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2580_0 <=( _mesh_19_16_io_out_id_0) ^ ((fiEnable && (7717 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2581_0 <=( _mesh_20_16_io_out_id_0) ^ ((fiEnable && (7718 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2582_0 <=( _mesh_21_16_io_out_id_0) ^ ((fiEnable && (7719 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2583_0 <=( _mesh_22_16_io_out_id_0) ^ ((fiEnable && (7720 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2584_0 <=( _mesh_23_16_io_out_id_0) ^ ((fiEnable && (7721 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2585_0 <=( _mesh_24_16_io_out_id_0) ^ ((fiEnable && (7722 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2586_0 <=( _mesh_25_16_io_out_id_0) ^ ((fiEnable && (7723 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2587_0 <=( _mesh_26_16_io_out_id_0) ^ ((fiEnable && (7724 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2588_0 <=( _mesh_27_16_io_out_id_0) ^ ((fiEnable && (7725 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2589_0 <=( _mesh_28_16_io_out_id_0) ^ ((fiEnable && (7726 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2590_0 <=( _mesh_29_16_io_out_id_0) ^ ((fiEnable && (7727 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2591_0 <=( _mesh_30_16_io_out_id_0) ^ ((fiEnable && (7728 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2592_0 <=( io_in_id_17_0) ^ ((fiEnable && (7729 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2593_0 <=( _mesh_0_17_io_out_id_0) ^ ((fiEnable && (7730 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2594_0 <=( _mesh_1_17_io_out_id_0) ^ ((fiEnable && (7731 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2595_0 <=( _mesh_2_17_io_out_id_0) ^ ((fiEnable && (7732 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2596_0 <=( _mesh_3_17_io_out_id_0) ^ ((fiEnable && (7733 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2597_0 <=( _mesh_4_17_io_out_id_0) ^ ((fiEnable && (7734 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2598_0 <=( _mesh_5_17_io_out_id_0) ^ ((fiEnable && (7735 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2599_0 <=( _mesh_6_17_io_out_id_0) ^ ((fiEnable && (7736 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2600_0 <=( _mesh_7_17_io_out_id_0) ^ ((fiEnable && (7737 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2601_0 <=( _mesh_8_17_io_out_id_0) ^ ((fiEnable && (7738 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2602_0 <=( _mesh_9_17_io_out_id_0) ^ ((fiEnable && (7739 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2603_0 <=( _mesh_10_17_io_out_id_0) ^ ((fiEnable && (7740 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2604_0 <=( _mesh_11_17_io_out_id_0) ^ ((fiEnable && (7741 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2605_0 <=( _mesh_12_17_io_out_id_0) ^ ((fiEnable && (7742 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2606_0 <=( _mesh_13_17_io_out_id_0) ^ ((fiEnable && (7743 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2607_0 <=( _mesh_14_17_io_out_id_0) ^ ((fiEnable && (7744 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2608_0 <=( _mesh_15_17_io_out_id_0) ^ ((fiEnable && (7745 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2609_0 <=( _mesh_16_17_io_out_id_0) ^ ((fiEnable && (7746 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2610_0 <=( _mesh_17_17_io_out_id_0) ^ ((fiEnable && (7747 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2611_0 <=( _mesh_18_17_io_out_id_0) ^ ((fiEnable && (7748 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2612_0 <=( _mesh_19_17_io_out_id_0) ^ ((fiEnable && (7749 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2613_0 <=( _mesh_20_17_io_out_id_0) ^ ((fiEnable && (7750 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2614_0 <=( _mesh_21_17_io_out_id_0) ^ ((fiEnable && (7751 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2615_0 <=( _mesh_22_17_io_out_id_0) ^ ((fiEnable && (7752 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2616_0 <=( _mesh_23_17_io_out_id_0) ^ ((fiEnable && (7753 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2617_0 <=( _mesh_24_17_io_out_id_0) ^ ((fiEnable && (7754 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2618_0 <=( _mesh_25_17_io_out_id_0) ^ ((fiEnable && (7755 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2619_0 <=( _mesh_26_17_io_out_id_0) ^ ((fiEnable && (7756 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2620_0 <=( _mesh_27_17_io_out_id_0) ^ ((fiEnable && (7757 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2621_0 <=( _mesh_28_17_io_out_id_0) ^ ((fiEnable && (7758 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2622_0 <=( _mesh_29_17_io_out_id_0) ^ ((fiEnable && (7759 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2623_0 <=( _mesh_30_17_io_out_id_0) ^ ((fiEnable && (7760 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2624_0 <=( io_in_id_18_0) ^ ((fiEnable && (7761 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2625_0 <=( _mesh_0_18_io_out_id_0) ^ ((fiEnable && (7762 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2626_0 <=( _mesh_1_18_io_out_id_0) ^ ((fiEnable && (7763 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2627_0 <=( _mesh_2_18_io_out_id_0) ^ ((fiEnable && (7764 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2628_0 <=( _mesh_3_18_io_out_id_0) ^ ((fiEnable && (7765 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2629_0 <=( _mesh_4_18_io_out_id_0) ^ ((fiEnable && (7766 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2630_0 <=( _mesh_5_18_io_out_id_0) ^ ((fiEnable && (7767 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2631_0 <=( _mesh_6_18_io_out_id_0) ^ ((fiEnable && (7768 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2632_0 <=( _mesh_7_18_io_out_id_0) ^ ((fiEnable && (7769 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2633_0 <=( _mesh_8_18_io_out_id_0) ^ ((fiEnable && (7770 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2634_0 <=( _mesh_9_18_io_out_id_0) ^ ((fiEnable && (7771 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2635_0 <=( _mesh_10_18_io_out_id_0) ^ ((fiEnable && (7772 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2636_0 <=( _mesh_11_18_io_out_id_0) ^ ((fiEnable && (7773 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2637_0 <=( _mesh_12_18_io_out_id_0) ^ ((fiEnable && (7774 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2638_0 <=( _mesh_13_18_io_out_id_0) ^ ((fiEnable && (7775 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2639_0 <=( _mesh_14_18_io_out_id_0) ^ ((fiEnable && (7776 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2640_0 <=( _mesh_15_18_io_out_id_0) ^ ((fiEnable && (7777 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2641_0 <=( _mesh_16_18_io_out_id_0) ^ ((fiEnable && (7778 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2642_0 <=( _mesh_17_18_io_out_id_0) ^ ((fiEnable && (7779 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2643_0 <=( _mesh_18_18_io_out_id_0) ^ ((fiEnable && (7780 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2644_0 <=( _mesh_19_18_io_out_id_0) ^ ((fiEnable && (7781 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2645_0 <=( _mesh_20_18_io_out_id_0) ^ ((fiEnable && (7782 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2646_0 <=( _mesh_21_18_io_out_id_0) ^ ((fiEnable && (7783 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2647_0 <=( _mesh_22_18_io_out_id_0) ^ ((fiEnable && (7784 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2648_0 <=( _mesh_23_18_io_out_id_0) ^ ((fiEnable && (7785 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2649_0 <=( _mesh_24_18_io_out_id_0) ^ ((fiEnable && (7786 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2650_0 <=( _mesh_25_18_io_out_id_0) ^ ((fiEnable && (7787 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2651_0 <=( _mesh_26_18_io_out_id_0) ^ ((fiEnable && (7788 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2652_0 <=( _mesh_27_18_io_out_id_0) ^ ((fiEnable && (7789 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2653_0 <=( _mesh_28_18_io_out_id_0) ^ ((fiEnable && (7790 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2654_0 <=( _mesh_29_18_io_out_id_0) ^ ((fiEnable && (7791 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2655_0 <=( _mesh_30_18_io_out_id_0) ^ ((fiEnable && (7792 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2656_0 <=( io_in_id_19_0) ^ ((fiEnable && (7793 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2657_0 <=( _mesh_0_19_io_out_id_0) ^ ((fiEnable && (7794 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2658_0 <=( _mesh_1_19_io_out_id_0) ^ ((fiEnable && (7795 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2659_0 <=( _mesh_2_19_io_out_id_0) ^ ((fiEnable && (7796 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2660_0 <=( _mesh_3_19_io_out_id_0) ^ ((fiEnable && (7797 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2661_0 <=( _mesh_4_19_io_out_id_0) ^ ((fiEnable && (7798 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2662_0 <=( _mesh_5_19_io_out_id_0) ^ ((fiEnable && (7799 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2663_0 <=( _mesh_6_19_io_out_id_0) ^ ((fiEnable && (7800 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2664_0 <=( _mesh_7_19_io_out_id_0) ^ ((fiEnable && (7801 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2665_0 <=( _mesh_8_19_io_out_id_0) ^ ((fiEnable && (7802 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2666_0 <=( _mesh_9_19_io_out_id_0) ^ ((fiEnable && (7803 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2667_0 <=( _mesh_10_19_io_out_id_0) ^ ((fiEnable && (7804 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2668_0 <=( _mesh_11_19_io_out_id_0) ^ ((fiEnable && (7805 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2669_0 <=( _mesh_12_19_io_out_id_0) ^ ((fiEnable && (7806 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2670_0 <=( _mesh_13_19_io_out_id_0) ^ ((fiEnable && (7807 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2671_0 <=( _mesh_14_19_io_out_id_0) ^ ((fiEnable && (7808 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2672_0 <=( _mesh_15_19_io_out_id_0) ^ ((fiEnable && (7809 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2673_0 <=( _mesh_16_19_io_out_id_0) ^ ((fiEnable && (7810 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2674_0 <=( _mesh_17_19_io_out_id_0) ^ ((fiEnable && (7811 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2675_0 <=( _mesh_18_19_io_out_id_0) ^ ((fiEnable && (7812 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2676_0 <=( _mesh_19_19_io_out_id_0) ^ ((fiEnable && (7813 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2677_0 <=( _mesh_20_19_io_out_id_0) ^ ((fiEnable && (7814 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2678_0 <=( _mesh_21_19_io_out_id_0) ^ ((fiEnable && (7815 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2679_0 <=( _mesh_22_19_io_out_id_0) ^ ((fiEnable && (7816 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2680_0 <=( _mesh_23_19_io_out_id_0) ^ ((fiEnable && (7817 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2681_0 <=( _mesh_24_19_io_out_id_0) ^ ((fiEnable && (7818 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2682_0 <=( _mesh_25_19_io_out_id_0) ^ ((fiEnable && (7819 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2683_0 <=( _mesh_26_19_io_out_id_0) ^ ((fiEnable && (7820 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2684_0 <=( _mesh_27_19_io_out_id_0) ^ ((fiEnable && (7821 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2685_0 <=( _mesh_28_19_io_out_id_0) ^ ((fiEnable && (7822 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2686_0 <=( _mesh_29_19_io_out_id_0) ^ ((fiEnable && (7823 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2687_0 <=( _mesh_30_19_io_out_id_0) ^ ((fiEnable && (7824 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2688_0 <=( io_in_id_20_0) ^ ((fiEnable && (7825 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2689_0 <=( _mesh_0_20_io_out_id_0) ^ ((fiEnable && (7826 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2690_0 <=( _mesh_1_20_io_out_id_0) ^ ((fiEnable && (7827 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2691_0 <=( _mesh_2_20_io_out_id_0) ^ ((fiEnable && (7828 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2692_0 <=( _mesh_3_20_io_out_id_0) ^ ((fiEnable && (7829 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2693_0 <=( _mesh_4_20_io_out_id_0) ^ ((fiEnable && (7830 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2694_0 <=( _mesh_5_20_io_out_id_0) ^ ((fiEnable && (7831 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2695_0 <=( _mesh_6_20_io_out_id_0) ^ ((fiEnable && (7832 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2696_0 <=( _mesh_7_20_io_out_id_0) ^ ((fiEnable && (7833 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2697_0 <=( _mesh_8_20_io_out_id_0) ^ ((fiEnable && (7834 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2698_0 <=( _mesh_9_20_io_out_id_0) ^ ((fiEnable && (7835 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2699_0 <=( _mesh_10_20_io_out_id_0) ^ ((fiEnable && (7836 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2700_0 <=( _mesh_11_20_io_out_id_0) ^ ((fiEnable && (7837 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2701_0 <=( _mesh_12_20_io_out_id_0) ^ ((fiEnable && (7838 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2702_0 <=( _mesh_13_20_io_out_id_0) ^ ((fiEnable && (7839 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2703_0 <=( _mesh_14_20_io_out_id_0) ^ ((fiEnable && (7840 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2704_0 <=( _mesh_15_20_io_out_id_0) ^ ((fiEnable && (7841 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2705_0 <=( _mesh_16_20_io_out_id_0) ^ ((fiEnable && (7842 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2706_0 <=( _mesh_17_20_io_out_id_0) ^ ((fiEnable && (7843 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2707_0 <=( _mesh_18_20_io_out_id_0) ^ ((fiEnable && (7844 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2708_0 <=( _mesh_19_20_io_out_id_0) ^ ((fiEnable && (7845 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2709_0 <=( _mesh_20_20_io_out_id_0) ^ ((fiEnable && (7846 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2710_0 <=( _mesh_21_20_io_out_id_0) ^ ((fiEnable && (7847 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2711_0 <=( _mesh_22_20_io_out_id_0) ^ ((fiEnable && (7848 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2712_0 <=( _mesh_23_20_io_out_id_0) ^ ((fiEnable && (7849 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2713_0 <=( _mesh_24_20_io_out_id_0) ^ ((fiEnable && (7850 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2714_0 <=( _mesh_25_20_io_out_id_0) ^ ((fiEnable && (7851 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2715_0 <=( _mesh_26_20_io_out_id_0) ^ ((fiEnable && (7852 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2716_0 <=( _mesh_27_20_io_out_id_0) ^ ((fiEnable && (7853 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2717_0 <=( _mesh_28_20_io_out_id_0) ^ ((fiEnable && (7854 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2718_0 <=( _mesh_29_20_io_out_id_0) ^ ((fiEnable && (7855 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2719_0 <=( _mesh_30_20_io_out_id_0) ^ ((fiEnable && (7856 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2720_0 <=( io_in_id_21_0) ^ ((fiEnable && (7857 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2721_0 <=( _mesh_0_21_io_out_id_0) ^ ((fiEnable && (7858 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2722_0 <=( _mesh_1_21_io_out_id_0) ^ ((fiEnable && (7859 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2723_0 <=( _mesh_2_21_io_out_id_0) ^ ((fiEnable && (7860 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2724_0 <=( _mesh_3_21_io_out_id_0) ^ ((fiEnable && (7861 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2725_0 <=( _mesh_4_21_io_out_id_0) ^ ((fiEnable && (7862 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2726_0 <=( _mesh_5_21_io_out_id_0) ^ ((fiEnable && (7863 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2727_0 <=( _mesh_6_21_io_out_id_0) ^ ((fiEnable && (7864 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2728_0 <=( _mesh_7_21_io_out_id_0) ^ ((fiEnable && (7865 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2729_0 <=( _mesh_8_21_io_out_id_0) ^ ((fiEnable && (7866 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2730_0 <=( _mesh_9_21_io_out_id_0) ^ ((fiEnable && (7867 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2731_0 <=( _mesh_10_21_io_out_id_0) ^ ((fiEnable && (7868 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2732_0 <=( _mesh_11_21_io_out_id_0) ^ ((fiEnable && (7869 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2733_0 <=( _mesh_12_21_io_out_id_0) ^ ((fiEnable && (7870 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2734_0 <=( _mesh_13_21_io_out_id_0) ^ ((fiEnable && (7871 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2735_0 <=( _mesh_14_21_io_out_id_0) ^ ((fiEnable && (7872 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2736_0 <=( _mesh_15_21_io_out_id_0) ^ ((fiEnable && (7873 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2737_0 <=( _mesh_16_21_io_out_id_0) ^ ((fiEnable && (7874 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2738_0 <=( _mesh_17_21_io_out_id_0) ^ ((fiEnable && (7875 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2739_0 <=( _mesh_18_21_io_out_id_0) ^ ((fiEnable && (7876 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2740_0 <=( _mesh_19_21_io_out_id_0) ^ ((fiEnable && (7877 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2741_0 <=( _mesh_20_21_io_out_id_0) ^ ((fiEnable && (7878 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2742_0 <=( _mesh_21_21_io_out_id_0) ^ ((fiEnable && (7879 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2743_0 <=( _mesh_22_21_io_out_id_0) ^ ((fiEnable && (7880 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2744_0 <=( _mesh_23_21_io_out_id_0) ^ ((fiEnable && (7881 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2745_0 <=( _mesh_24_21_io_out_id_0) ^ ((fiEnable && (7882 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2746_0 <=( _mesh_25_21_io_out_id_0) ^ ((fiEnable && (7883 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2747_0 <=( _mesh_26_21_io_out_id_0) ^ ((fiEnable && (7884 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2748_0 <=( _mesh_27_21_io_out_id_0) ^ ((fiEnable && (7885 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2749_0 <=( _mesh_28_21_io_out_id_0) ^ ((fiEnable && (7886 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2750_0 <=( _mesh_29_21_io_out_id_0) ^ ((fiEnable && (7887 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2751_0 <=( _mesh_30_21_io_out_id_0) ^ ((fiEnable && (7888 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2752_0 <=( io_in_id_22_0) ^ ((fiEnable && (7889 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2753_0 <=( _mesh_0_22_io_out_id_0) ^ ((fiEnable && (7890 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2754_0 <=( _mesh_1_22_io_out_id_0) ^ ((fiEnable && (7891 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2755_0 <=( _mesh_2_22_io_out_id_0) ^ ((fiEnable && (7892 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2756_0 <=( _mesh_3_22_io_out_id_0) ^ ((fiEnable && (7893 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2757_0 <=( _mesh_4_22_io_out_id_0) ^ ((fiEnable && (7894 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2758_0 <=( _mesh_5_22_io_out_id_0) ^ ((fiEnable && (7895 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2759_0 <=( _mesh_6_22_io_out_id_0) ^ ((fiEnable && (7896 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2760_0 <=( _mesh_7_22_io_out_id_0) ^ ((fiEnable && (7897 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2761_0 <=( _mesh_8_22_io_out_id_0) ^ ((fiEnable && (7898 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2762_0 <=( _mesh_9_22_io_out_id_0) ^ ((fiEnable && (7899 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2763_0 <=( _mesh_10_22_io_out_id_0) ^ ((fiEnable && (7900 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2764_0 <=( _mesh_11_22_io_out_id_0) ^ ((fiEnable && (7901 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2765_0 <=( _mesh_12_22_io_out_id_0) ^ ((fiEnable && (7902 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2766_0 <=( _mesh_13_22_io_out_id_0) ^ ((fiEnable && (7903 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2767_0 <=( _mesh_14_22_io_out_id_0) ^ ((fiEnable && (7904 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2768_0 <=( _mesh_15_22_io_out_id_0) ^ ((fiEnable && (7905 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2769_0 <=( _mesh_16_22_io_out_id_0) ^ ((fiEnable && (7906 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2770_0 <=( _mesh_17_22_io_out_id_0) ^ ((fiEnable && (7907 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2771_0 <=( _mesh_18_22_io_out_id_0) ^ ((fiEnable && (7908 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2772_0 <=( _mesh_19_22_io_out_id_0) ^ ((fiEnable && (7909 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2773_0 <=( _mesh_20_22_io_out_id_0) ^ ((fiEnable && (7910 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2774_0 <=( _mesh_21_22_io_out_id_0) ^ ((fiEnable && (7911 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2775_0 <=( _mesh_22_22_io_out_id_0) ^ ((fiEnable && (7912 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2776_0 <=( _mesh_23_22_io_out_id_0) ^ ((fiEnable && (7913 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2777_0 <=( _mesh_24_22_io_out_id_0) ^ ((fiEnable && (7914 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2778_0 <=( _mesh_25_22_io_out_id_0) ^ ((fiEnable && (7915 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2779_0 <=( _mesh_26_22_io_out_id_0) ^ ((fiEnable && (7916 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2780_0 <=( _mesh_27_22_io_out_id_0) ^ ((fiEnable && (7917 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2781_0 <=( _mesh_28_22_io_out_id_0) ^ ((fiEnable && (7918 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2782_0 <=( _mesh_29_22_io_out_id_0) ^ ((fiEnable && (7919 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2783_0 <=( _mesh_30_22_io_out_id_0) ^ ((fiEnable && (7920 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2784_0 <=( io_in_id_23_0) ^ ((fiEnable && (7921 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2785_0 <=( _mesh_0_23_io_out_id_0) ^ ((fiEnable && (7922 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2786_0 <=( _mesh_1_23_io_out_id_0) ^ ((fiEnable && (7923 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2787_0 <=( _mesh_2_23_io_out_id_0) ^ ((fiEnable && (7924 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2788_0 <=( _mesh_3_23_io_out_id_0) ^ ((fiEnable && (7925 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2789_0 <=( _mesh_4_23_io_out_id_0) ^ ((fiEnable && (7926 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2790_0 <=( _mesh_5_23_io_out_id_0) ^ ((fiEnable && (7927 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2791_0 <=( _mesh_6_23_io_out_id_0) ^ ((fiEnable && (7928 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2792_0 <=( _mesh_7_23_io_out_id_0) ^ ((fiEnable && (7929 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2793_0 <=( _mesh_8_23_io_out_id_0) ^ ((fiEnable && (7930 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2794_0 <=( _mesh_9_23_io_out_id_0) ^ ((fiEnable && (7931 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2795_0 <=( _mesh_10_23_io_out_id_0) ^ ((fiEnable && (7932 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2796_0 <=( _mesh_11_23_io_out_id_0) ^ ((fiEnable && (7933 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2797_0 <=( _mesh_12_23_io_out_id_0) ^ ((fiEnable && (7934 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2798_0 <=( _mesh_13_23_io_out_id_0) ^ ((fiEnable && (7935 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2799_0 <=( _mesh_14_23_io_out_id_0) ^ ((fiEnable && (7936 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2800_0 <=( _mesh_15_23_io_out_id_0) ^ ((fiEnable && (7937 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2801_0 <=( _mesh_16_23_io_out_id_0) ^ ((fiEnable && (7938 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2802_0 <=( _mesh_17_23_io_out_id_0) ^ ((fiEnable && (7939 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2803_0 <=( _mesh_18_23_io_out_id_0) ^ ((fiEnable && (7940 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2804_0 <=( _mesh_19_23_io_out_id_0) ^ ((fiEnable && (7941 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2805_0 <=( _mesh_20_23_io_out_id_0) ^ ((fiEnable && (7942 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2806_0 <=( _mesh_21_23_io_out_id_0) ^ ((fiEnable && (7943 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2807_0 <=( _mesh_22_23_io_out_id_0) ^ ((fiEnable && (7944 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2808_0 <=( _mesh_23_23_io_out_id_0) ^ ((fiEnable && (7945 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2809_0 <=( _mesh_24_23_io_out_id_0) ^ ((fiEnable && (7946 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2810_0 <=( _mesh_25_23_io_out_id_0) ^ ((fiEnable && (7947 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2811_0 <=( _mesh_26_23_io_out_id_0) ^ ((fiEnable && (7948 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2812_0 <=( _mesh_27_23_io_out_id_0) ^ ((fiEnable && (7949 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2813_0 <=( _mesh_28_23_io_out_id_0) ^ ((fiEnable && (7950 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2814_0 <=( _mesh_29_23_io_out_id_0) ^ ((fiEnable && (7951 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2815_0 <=( _mesh_30_23_io_out_id_0) ^ ((fiEnable && (7952 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2816_0 <=( io_in_id_24_0) ^ ((fiEnable && (7953 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2817_0 <=( _mesh_0_24_io_out_id_0) ^ ((fiEnable && (7954 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2818_0 <=( _mesh_1_24_io_out_id_0) ^ ((fiEnable && (7955 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2819_0 <=( _mesh_2_24_io_out_id_0) ^ ((fiEnable && (7956 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2820_0 <=( _mesh_3_24_io_out_id_0) ^ ((fiEnable && (7957 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2821_0 <=( _mesh_4_24_io_out_id_0) ^ ((fiEnable && (7958 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2822_0 <=( _mesh_5_24_io_out_id_0) ^ ((fiEnable && (7959 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2823_0 <=( _mesh_6_24_io_out_id_0) ^ ((fiEnable && (7960 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2824_0 <=( _mesh_7_24_io_out_id_0) ^ ((fiEnable && (7961 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2825_0 <=( _mesh_8_24_io_out_id_0) ^ ((fiEnable && (7962 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2826_0 <=( _mesh_9_24_io_out_id_0) ^ ((fiEnable && (7963 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2827_0 <=( _mesh_10_24_io_out_id_0) ^ ((fiEnable && (7964 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2828_0 <=( _mesh_11_24_io_out_id_0) ^ ((fiEnable && (7965 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2829_0 <=( _mesh_12_24_io_out_id_0) ^ ((fiEnable && (7966 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2830_0 <=( _mesh_13_24_io_out_id_0) ^ ((fiEnable && (7967 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2831_0 <=( _mesh_14_24_io_out_id_0) ^ ((fiEnable && (7968 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2832_0 <=( _mesh_15_24_io_out_id_0) ^ ((fiEnable && (7969 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2833_0 <=( _mesh_16_24_io_out_id_0) ^ ((fiEnable && (7970 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2834_0 <=( _mesh_17_24_io_out_id_0) ^ ((fiEnable && (7971 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2835_0 <=( _mesh_18_24_io_out_id_0) ^ ((fiEnable && (7972 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2836_0 <=( _mesh_19_24_io_out_id_0) ^ ((fiEnable && (7973 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2837_0 <=( _mesh_20_24_io_out_id_0) ^ ((fiEnable && (7974 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2838_0 <=( _mesh_21_24_io_out_id_0) ^ ((fiEnable && (7975 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2839_0 <=( _mesh_22_24_io_out_id_0) ^ ((fiEnable && (7976 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2840_0 <=( _mesh_23_24_io_out_id_0) ^ ((fiEnable && (7977 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2841_0 <=( _mesh_24_24_io_out_id_0) ^ ((fiEnable && (7978 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2842_0 <=( _mesh_25_24_io_out_id_0) ^ ((fiEnable && (7979 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2843_0 <=( _mesh_26_24_io_out_id_0) ^ ((fiEnable && (7980 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2844_0 <=( _mesh_27_24_io_out_id_0) ^ ((fiEnable && (7981 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2845_0 <=( _mesh_28_24_io_out_id_0) ^ ((fiEnable && (7982 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2846_0 <=( _mesh_29_24_io_out_id_0) ^ ((fiEnable && (7983 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2847_0 <=( _mesh_30_24_io_out_id_0) ^ ((fiEnable && (7984 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2848_0 <=( io_in_id_25_0) ^ ((fiEnable && (7985 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2849_0 <=( _mesh_0_25_io_out_id_0) ^ ((fiEnable && (7986 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2850_0 <=( _mesh_1_25_io_out_id_0) ^ ((fiEnable && (7987 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2851_0 <=( _mesh_2_25_io_out_id_0) ^ ((fiEnable && (7988 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2852_0 <=( _mesh_3_25_io_out_id_0) ^ ((fiEnable && (7989 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2853_0 <=( _mesh_4_25_io_out_id_0) ^ ((fiEnable && (7990 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2854_0 <=( _mesh_5_25_io_out_id_0) ^ ((fiEnable && (7991 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2855_0 <=( _mesh_6_25_io_out_id_0) ^ ((fiEnable && (7992 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2856_0 <=( _mesh_7_25_io_out_id_0) ^ ((fiEnable && (7993 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2857_0 <=( _mesh_8_25_io_out_id_0) ^ ((fiEnable && (7994 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2858_0 <=( _mesh_9_25_io_out_id_0) ^ ((fiEnable && (7995 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2859_0 <=( _mesh_10_25_io_out_id_0) ^ ((fiEnable && (7996 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2860_0 <=( _mesh_11_25_io_out_id_0) ^ ((fiEnable && (7997 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2861_0 <=( _mesh_12_25_io_out_id_0) ^ ((fiEnable && (7998 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2862_0 <=( _mesh_13_25_io_out_id_0) ^ ((fiEnable && (7999 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2863_0 <=( _mesh_14_25_io_out_id_0) ^ ((fiEnable && (8000 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2864_0 <=( _mesh_15_25_io_out_id_0) ^ ((fiEnable && (8001 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2865_0 <=( _mesh_16_25_io_out_id_0) ^ ((fiEnable && (8002 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2866_0 <=( _mesh_17_25_io_out_id_0) ^ ((fiEnable && (8003 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2867_0 <=( _mesh_18_25_io_out_id_0) ^ ((fiEnable && (8004 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2868_0 <=( _mesh_19_25_io_out_id_0) ^ ((fiEnable && (8005 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2869_0 <=( _mesh_20_25_io_out_id_0) ^ ((fiEnable && (8006 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2870_0 <=( _mesh_21_25_io_out_id_0) ^ ((fiEnable && (8007 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2871_0 <=( _mesh_22_25_io_out_id_0) ^ ((fiEnable && (8008 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2872_0 <=( _mesh_23_25_io_out_id_0) ^ ((fiEnable && (8009 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2873_0 <=( _mesh_24_25_io_out_id_0) ^ ((fiEnable && (8010 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2874_0 <=( _mesh_25_25_io_out_id_0) ^ ((fiEnable && (8011 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2875_0 <=( _mesh_26_25_io_out_id_0) ^ ((fiEnable && (8012 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2876_0 <=( _mesh_27_25_io_out_id_0) ^ ((fiEnable && (8013 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2877_0 <=( _mesh_28_25_io_out_id_0) ^ ((fiEnable && (8014 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2878_0 <=( _mesh_29_25_io_out_id_0) ^ ((fiEnable && (8015 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2879_0 <=( _mesh_30_25_io_out_id_0) ^ ((fiEnable && (8016 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2880_0 <=( io_in_id_26_0) ^ ((fiEnable && (8017 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2881_0 <=( _mesh_0_26_io_out_id_0) ^ ((fiEnable && (8018 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2882_0 <=( _mesh_1_26_io_out_id_0) ^ ((fiEnable && (8019 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2883_0 <=( _mesh_2_26_io_out_id_0) ^ ((fiEnable && (8020 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2884_0 <=( _mesh_3_26_io_out_id_0) ^ ((fiEnable && (8021 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2885_0 <=( _mesh_4_26_io_out_id_0) ^ ((fiEnable && (8022 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2886_0 <=( _mesh_5_26_io_out_id_0) ^ ((fiEnable && (8023 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2887_0 <=( _mesh_6_26_io_out_id_0) ^ ((fiEnable && (8024 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2888_0 <=( _mesh_7_26_io_out_id_0) ^ ((fiEnable && (8025 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2889_0 <=( _mesh_8_26_io_out_id_0) ^ ((fiEnable && (8026 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2890_0 <=( _mesh_9_26_io_out_id_0) ^ ((fiEnable && (8027 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2891_0 <=( _mesh_10_26_io_out_id_0) ^ ((fiEnable && (8028 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2892_0 <=( _mesh_11_26_io_out_id_0) ^ ((fiEnable && (8029 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2893_0 <=( _mesh_12_26_io_out_id_0) ^ ((fiEnable && (8030 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2894_0 <=( _mesh_13_26_io_out_id_0) ^ ((fiEnable && (8031 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2895_0 <=( _mesh_14_26_io_out_id_0) ^ ((fiEnable && (8032 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2896_0 <=( _mesh_15_26_io_out_id_0) ^ ((fiEnable && (8033 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2897_0 <=( _mesh_16_26_io_out_id_0) ^ ((fiEnable && (8034 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2898_0 <=( _mesh_17_26_io_out_id_0) ^ ((fiEnable && (8035 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2899_0 <=( _mesh_18_26_io_out_id_0) ^ ((fiEnable && (8036 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2900_0 <=( _mesh_19_26_io_out_id_0) ^ ((fiEnable && (8037 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2901_0 <=( _mesh_20_26_io_out_id_0) ^ ((fiEnable && (8038 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2902_0 <=( _mesh_21_26_io_out_id_0) ^ ((fiEnable && (8039 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2903_0 <=( _mesh_22_26_io_out_id_0) ^ ((fiEnable && (8040 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2904_0 <=( _mesh_23_26_io_out_id_0) ^ ((fiEnable && (8041 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2905_0 <=( _mesh_24_26_io_out_id_0) ^ ((fiEnable && (8042 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2906_0 <=( _mesh_25_26_io_out_id_0) ^ ((fiEnable && (8043 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2907_0 <=( _mesh_26_26_io_out_id_0) ^ ((fiEnable && (8044 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2908_0 <=( _mesh_27_26_io_out_id_0) ^ ((fiEnable && (8045 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2909_0 <=( _mesh_28_26_io_out_id_0) ^ ((fiEnable && (8046 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2910_0 <=( _mesh_29_26_io_out_id_0) ^ ((fiEnable && (8047 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2911_0 <=( _mesh_30_26_io_out_id_0) ^ ((fiEnable && (8048 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2912_0 <=( io_in_id_27_0) ^ ((fiEnable && (8049 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2913_0 <=( _mesh_0_27_io_out_id_0) ^ ((fiEnable && (8050 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2914_0 <=( _mesh_1_27_io_out_id_0) ^ ((fiEnable && (8051 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2915_0 <=( _mesh_2_27_io_out_id_0) ^ ((fiEnable && (8052 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2916_0 <=( _mesh_3_27_io_out_id_0) ^ ((fiEnable && (8053 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2917_0 <=( _mesh_4_27_io_out_id_0) ^ ((fiEnable && (8054 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2918_0 <=( _mesh_5_27_io_out_id_0) ^ ((fiEnable && (8055 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2919_0 <=( _mesh_6_27_io_out_id_0) ^ ((fiEnable && (8056 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2920_0 <=( _mesh_7_27_io_out_id_0) ^ ((fiEnable && (8057 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2921_0 <=( _mesh_8_27_io_out_id_0) ^ ((fiEnable && (8058 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2922_0 <=( _mesh_9_27_io_out_id_0) ^ ((fiEnable && (8059 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2923_0 <=( _mesh_10_27_io_out_id_0) ^ ((fiEnable && (8060 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2924_0 <=( _mesh_11_27_io_out_id_0) ^ ((fiEnable && (8061 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2925_0 <=( _mesh_12_27_io_out_id_0) ^ ((fiEnable && (8062 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2926_0 <=( _mesh_13_27_io_out_id_0) ^ ((fiEnable && (8063 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2927_0 <=( _mesh_14_27_io_out_id_0) ^ ((fiEnable && (8064 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2928_0 <=( _mesh_15_27_io_out_id_0) ^ ((fiEnable && (8065 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2929_0 <=( _mesh_16_27_io_out_id_0) ^ ((fiEnable && (8066 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2930_0 <=( _mesh_17_27_io_out_id_0) ^ ((fiEnable && (8067 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2931_0 <=( _mesh_18_27_io_out_id_0) ^ ((fiEnable && (8068 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2932_0 <=( _mesh_19_27_io_out_id_0) ^ ((fiEnable && (8069 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2933_0 <=( _mesh_20_27_io_out_id_0) ^ ((fiEnable && (8070 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2934_0 <=( _mesh_21_27_io_out_id_0) ^ ((fiEnable && (8071 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2935_0 <=( _mesh_22_27_io_out_id_0) ^ ((fiEnable && (8072 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2936_0 <=( _mesh_23_27_io_out_id_0) ^ ((fiEnable && (8073 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2937_0 <=( _mesh_24_27_io_out_id_0) ^ ((fiEnable && (8074 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2938_0 <=( _mesh_25_27_io_out_id_0) ^ ((fiEnable && (8075 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2939_0 <=( _mesh_26_27_io_out_id_0) ^ ((fiEnable && (8076 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2940_0 <=( _mesh_27_27_io_out_id_0) ^ ((fiEnable && (8077 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2941_0 <=( _mesh_28_27_io_out_id_0) ^ ((fiEnable && (8078 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2942_0 <=( _mesh_29_27_io_out_id_0) ^ ((fiEnable && (8079 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2943_0 <=( _mesh_30_27_io_out_id_0) ^ ((fiEnable && (8080 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2944_0 <=( io_in_id_28_0) ^ ((fiEnable && (8081 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2945_0 <=( _mesh_0_28_io_out_id_0) ^ ((fiEnable && (8082 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2946_0 <=( _mesh_1_28_io_out_id_0) ^ ((fiEnable && (8083 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2947_0 <=( _mesh_2_28_io_out_id_0) ^ ((fiEnable && (8084 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2948_0 <=( _mesh_3_28_io_out_id_0) ^ ((fiEnable && (8085 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2949_0 <=( _mesh_4_28_io_out_id_0) ^ ((fiEnable && (8086 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2950_0 <=( _mesh_5_28_io_out_id_0) ^ ((fiEnable && (8087 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2951_0 <=( _mesh_6_28_io_out_id_0) ^ ((fiEnable && (8088 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2952_0 <=( _mesh_7_28_io_out_id_0) ^ ((fiEnable && (8089 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2953_0 <=( _mesh_8_28_io_out_id_0) ^ ((fiEnable && (8090 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2954_0 <=( _mesh_9_28_io_out_id_0) ^ ((fiEnable && (8091 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2955_0 <=( _mesh_10_28_io_out_id_0) ^ ((fiEnable && (8092 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2956_0 <=( _mesh_11_28_io_out_id_0) ^ ((fiEnable && (8093 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2957_0 <=( _mesh_12_28_io_out_id_0) ^ ((fiEnable && (8094 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2958_0 <=( _mesh_13_28_io_out_id_0) ^ ((fiEnable && (8095 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2959_0 <=( _mesh_14_28_io_out_id_0) ^ ((fiEnable && (8096 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2960_0 <=( _mesh_15_28_io_out_id_0) ^ ((fiEnable && (8097 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2961_0 <=( _mesh_16_28_io_out_id_0) ^ ((fiEnable && (8098 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2962_0 <=( _mesh_17_28_io_out_id_0) ^ ((fiEnable && (8099 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2963_0 <=( _mesh_18_28_io_out_id_0) ^ ((fiEnable && (8100 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2964_0 <=( _mesh_19_28_io_out_id_0) ^ ((fiEnable && (8101 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2965_0 <=( _mesh_20_28_io_out_id_0) ^ ((fiEnable && (8102 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2966_0 <=( _mesh_21_28_io_out_id_0) ^ ((fiEnable && (8103 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2967_0 <=( _mesh_22_28_io_out_id_0) ^ ((fiEnable && (8104 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2968_0 <=( _mesh_23_28_io_out_id_0) ^ ((fiEnable && (8105 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2969_0 <=( _mesh_24_28_io_out_id_0) ^ ((fiEnable && (8106 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2970_0 <=( _mesh_25_28_io_out_id_0) ^ ((fiEnable && (8107 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2971_0 <=( _mesh_26_28_io_out_id_0) ^ ((fiEnable && (8108 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2972_0 <=( _mesh_27_28_io_out_id_0) ^ ((fiEnable && (8109 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2973_0 <=( _mesh_28_28_io_out_id_0) ^ ((fiEnable && (8110 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2974_0 <=( _mesh_29_28_io_out_id_0) ^ ((fiEnable && (8111 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2975_0 <=( _mesh_30_28_io_out_id_0) ^ ((fiEnable && (8112 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2976_0 <=( io_in_id_29_0) ^ ((fiEnable && (8113 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2977_0 <=( _mesh_0_29_io_out_id_0) ^ ((fiEnable && (8114 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2978_0 <=( _mesh_1_29_io_out_id_0) ^ ((fiEnable && (8115 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2979_0 <=( _mesh_2_29_io_out_id_0) ^ ((fiEnable && (8116 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2980_0 <=( _mesh_3_29_io_out_id_0) ^ ((fiEnable && (8117 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2981_0 <=( _mesh_4_29_io_out_id_0) ^ ((fiEnable && (8118 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2982_0 <=( _mesh_5_29_io_out_id_0) ^ ((fiEnable && (8119 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2983_0 <=( _mesh_6_29_io_out_id_0) ^ ((fiEnable && (8120 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2984_0 <=( _mesh_7_29_io_out_id_0) ^ ((fiEnable && (8121 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2985_0 <=( _mesh_8_29_io_out_id_0) ^ ((fiEnable && (8122 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2986_0 <=( _mesh_9_29_io_out_id_0) ^ ((fiEnable && (8123 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2987_0 <=( _mesh_10_29_io_out_id_0) ^ ((fiEnable && (8124 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2988_0 <=( _mesh_11_29_io_out_id_0) ^ ((fiEnable && (8125 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2989_0 <=( _mesh_12_29_io_out_id_0) ^ ((fiEnable && (8126 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2990_0 <=( _mesh_13_29_io_out_id_0) ^ ((fiEnable && (8127 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2991_0 <=( _mesh_14_29_io_out_id_0) ^ ((fiEnable && (8128 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2992_0 <=( _mesh_15_29_io_out_id_0) ^ ((fiEnable && (8129 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2993_0 <=( _mesh_16_29_io_out_id_0) ^ ((fiEnable && (8130 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2994_0 <=( _mesh_17_29_io_out_id_0) ^ ((fiEnable && (8131 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2995_0 <=( _mesh_18_29_io_out_id_0) ^ ((fiEnable && (8132 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2996_0 <=( _mesh_19_29_io_out_id_0) ^ ((fiEnable && (8133 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2997_0 <=( _mesh_20_29_io_out_id_0) ^ ((fiEnable && (8134 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2998_0 <=( _mesh_21_29_io_out_id_0) ^ ((fiEnable && (8135 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_2999_0 <=( _mesh_22_29_io_out_id_0) ^ ((fiEnable && (8136 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3000_0 <=( _mesh_23_29_io_out_id_0) ^ ((fiEnable && (8137 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3001_0 <=( _mesh_24_29_io_out_id_0) ^ ((fiEnable && (8138 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3002_0 <=( _mesh_25_29_io_out_id_0) ^ ((fiEnable && (8139 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3003_0 <=( _mesh_26_29_io_out_id_0) ^ ((fiEnable && (8140 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3004_0 <=( _mesh_27_29_io_out_id_0) ^ ((fiEnable && (8141 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3005_0 <=( _mesh_28_29_io_out_id_0) ^ ((fiEnable && (8142 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3006_0 <=( _mesh_29_29_io_out_id_0) ^ ((fiEnable && (8143 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3007_0 <=( _mesh_30_29_io_out_id_0) ^ ((fiEnable && (8144 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3008_0 <=( io_in_id_30_0) ^ ((fiEnable && (8145 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3009_0 <=( _mesh_0_30_io_out_id_0) ^ ((fiEnable && (8146 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3010_0 <=( _mesh_1_30_io_out_id_0) ^ ((fiEnable && (8147 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3011_0 <=( _mesh_2_30_io_out_id_0) ^ ((fiEnable && (8148 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3012_0 <=( _mesh_3_30_io_out_id_0) ^ ((fiEnable && (8149 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3013_0 <=( _mesh_4_30_io_out_id_0) ^ ((fiEnable && (8150 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3014_0 <=( _mesh_5_30_io_out_id_0) ^ ((fiEnable && (8151 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3015_0 <=( _mesh_6_30_io_out_id_0) ^ ((fiEnable && (8152 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3016_0 <=( _mesh_7_30_io_out_id_0) ^ ((fiEnable && (8153 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3017_0 <=( _mesh_8_30_io_out_id_0) ^ ((fiEnable && (8154 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3018_0 <=( _mesh_9_30_io_out_id_0) ^ ((fiEnable && (8155 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3019_0 <=( _mesh_10_30_io_out_id_0) ^ ((fiEnable && (8156 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3020_0 <=( _mesh_11_30_io_out_id_0) ^ ((fiEnable && (8157 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3021_0 <=( _mesh_12_30_io_out_id_0) ^ ((fiEnable && (8158 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3022_0 <=( _mesh_13_30_io_out_id_0) ^ ((fiEnable && (8159 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3023_0 <=( _mesh_14_30_io_out_id_0) ^ ((fiEnable && (8160 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3024_0 <=( _mesh_15_30_io_out_id_0) ^ ((fiEnable && (8161 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3025_0 <=( _mesh_16_30_io_out_id_0) ^ ((fiEnable && (8162 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3026_0 <=( _mesh_17_30_io_out_id_0) ^ ((fiEnable && (8163 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3027_0 <=( _mesh_18_30_io_out_id_0) ^ ((fiEnable && (8164 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3028_0 <=( _mesh_19_30_io_out_id_0) ^ ((fiEnable && (8165 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3029_0 <=( _mesh_20_30_io_out_id_0) ^ ((fiEnable && (8166 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3030_0 <=( _mesh_21_30_io_out_id_0) ^ ((fiEnable && (8167 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3031_0 <=( _mesh_22_30_io_out_id_0) ^ ((fiEnable && (8168 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3032_0 <=( _mesh_23_30_io_out_id_0) ^ ((fiEnable && (8169 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3033_0 <=( _mesh_24_30_io_out_id_0) ^ ((fiEnable && (8170 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3034_0 <=( _mesh_25_30_io_out_id_0) ^ ((fiEnable && (8171 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3035_0 <=( _mesh_26_30_io_out_id_0) ^ ((fiEnable && (8172 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3036_0 <=( _mesh_27_30_io_out_id_0) ^ ((fiEnable && (8173 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3037_0 <=( _mesh_28_30_io_out_id_0) ^ ((fiEnable && (8174 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3038_0 <=( _mesh_29_30_io_out_id_0) ^ ((fiEnable && (8175 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3039_0 <=( _mesh_30_30_io_out_id_0) ^ ((fiEnable && (8176 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3040_0 <=( io_in_id_31_0) ^ ((fiEnable && (8177 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3041_0 <=( _mesh_0_31_io_out_id_0) ^ ((fiEnable && (8178 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3042_0 <=( _mesh_1_31_io_out_id_0) ^ ((fiEnable && (8179 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3043_0 <=( _mesh_2_31_io_out_id_0) ^ ((fiEnable && (8180 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3044_0 <=( _mesh_3_31_io_out_id_0) ^ ((fiEnable && (8181 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3045_0 <=( _mesh_4_31_io_out_id_0) ^ ((fiEnable && (8182 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3046_0 <=( _mesh_5_31_io_out_id_0) ^ ((fiEnable && (8183 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3047_0 <=( _mesh_6_31_io_out_id_0) ^ ((fiEnable && (8184 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3048_0 <=( _mesh_7_31_io_out_id_0) ^ ((fiEnable && (8185 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3049_0 <=( _mesh_8_31_io_out_id_0) ^ ((fiEnable && (8186 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3050_0 <=( _mesh_9_31_io_out_id_0) ^ ((fiEnable && (8187 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3051_0 <=( _mesh_10_31_io_out_id_0) ^ ((fiEnable && (8188 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3052_0 <=( _mesh_11_31_io_out_id_0) ^ ((fiEnable && (8189 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3053_0 <=( _mesh_12_31_io_out_id_0) ^ ((fiEnable && (8190 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3054_0 <=( _mesh_13_31_io_out_id_0) ^ ((fiEnable && (8191 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3055_0 <=( _mesh_14_31_io_out_id_0) ^ ((fiEnable && (8192 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3056_0 <=( _mesh_15_31_io_out_id_0) ^ ((fiEnable && (8193 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3057_0 <=( _mesh_16_31_io_out_id_0) ^ ((fiEnable && (8194 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3058_0 <=( _mesh_17_31_io_out_id_0) ^ ((fiEnable && (8195 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3059_0 <=( _mesh_18_31_io_out_id_0) ^ ((fiEnable && (8196 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3060_0 <=( _mesh_19_31_io_out_id_0) ^ ((fiEnable && (8197 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3061_0 <=( _mesh_20_31_io_out_id_0) ^ ((fiEnable && (8198 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3062_0 <=( _mesh_21_31_io_out_id_0) ^ ((fiEnable && (8199 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3063_0 <=( _mesh_22_31_io_out_id_0) ^ ((fiEnable && (8200 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3064_0 <=( _mesh_23_31_io_out_id_0) ^ ((fiEnable && (8201 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3065_0 <=( _mesh_24_31_io_out_id_0) ^ ((fiEnable && (8202 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3066_0 <=( _mesh_25_31_io_out_id_0) ^ ((fiEnable && (8203 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3067_0 <=( _mesh_26_31_io_out_id_0) ^ ((fiEnable && (8204 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3068_0 <=( _mesh_27_31_io_out_id_0) ^ ((fiEnable && (8205 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3069_0 <=( _mesh_28_31_io_out_id_0) ^ ((fiEnable && (8206 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3070_0 <=( _mesh_29_31_io_out_id_0) ^ ((fiEnable && (8207 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3071_0 <=( _mesh_30_31_io_out_id_0) ^ ((fiEnable && (8208 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_3072_0 <=( io_in_last_0_0) ^ ((fiEnable && (8209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3073_0 <=( _mesh_0_0_io_out_last_0) ^ ((fiEnable && (8210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3074_0 <=( _mesh_1_0_io_out_last_0) ^ ((fiEnable && (8211 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3075_0 <=( _mesh_2_0_io_out_last_0) ^ ((fiEnable && (8212 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3076_0 <=( _mesh_3_0_io_out_last_0) ^ ((fiEnable && (8213 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3077_0 <=( _mesh_4_0_io_out_last_0) ^ ((fiEnable && (8214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3078_0 <=( _mesh_5_0_io_out_last_0) ^ ((fiEnable && (8215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3079_0 <=( _mesh_6_0_io_out_last_0) ^ ((fiEnable && (8216 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3080_0 <=( _mesh_7_0_io_out_last_0) ^ ((fiEnable && (8217 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3081_0 <=( _mesh_8_0_io_out_last_0) ^ ((fiEnable && (8218 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3082_0 <=( _mesh_9_0_io_out_last_0) ^ ((fiEnable && (8219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3083_0 <=( _mesh_10_0_io_out_last_0) ^ ((fiEnable && (8220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3084_0 <=( _mesh_11_0_io_out_last_0) ^ ((fiEnable && (8221 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3085_0 <=( _mesh_12_0_io_out_last_0) ^ ((fiEnable && (8222 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3086_0 <=( _mesh_13_0_io_out_last_0) ^ ((fiEnable && (8223 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3087_0 <=( _mesh_14_0_io_out_last_0) ^ ((fiEnable && (8224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3088_0 <=( _mesh_15_0_io_out_last_0) ^ ((fiEnable && (8225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3089_0 <=( _mesh_16_0_io_out_last_0) ^ ((fiEnable && (8226 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3090_0 <=( _mesh_17_0_io_out_last_0) ^ ((fiEnable && (8227 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3091_0 <=( _mesh_18_0_io_out_last_0) ^ ((fiEnable && (8228 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3092_0 <=( _mesh_19_0_io_out_last_0) ^ ((fiEnable && (8229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3093_0 <=( _mesh_20_0_io_out_last_0) ^ ((fiEnable && (8230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3094_0 <=( _mesh_21_0_io_out_last_0) ^ ((fiEnable && (8231 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3095_0 <=( _mesh_22_0_io_out_last_0) ^ ((fiEnable && (8232 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3096_0 <=( _mesh_23_0_io_out_last_0) ^ ((fiEnable && (8233 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3097_0 <=( _mesh_24_0_io_out_last_0) ^ ((fiEnable && (8234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3098_0 <=( _mesh_25_0_io_out_last_0) ^ ((fiEnable && (8235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3099_0 <=( _mesh_26_0_io_out_last_0) ^ ((fiEnable && (8236 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3100_0 <=( _mesh_27_0_io_out_last_0) ^ ((fiEnable && (8237 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3101_0 <=( _mesh_28_0_io_out_last_0) ^ ((fiEnable && (8238 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3102_0 <=( _mesh_29_0_io_out_last_0) ^ ((fiEnable && (8239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3103_0 <=( _mesh_30_0_io_out_last_0) ^ ((fiEnable && (8240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3104_0 <=( io_in_last_1_0) ^ ((fiEnable && (8241 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3105_0 <=( _mesh_0_1_io_out_last_0) ^ ((fiEnable && (8242 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3106_0 <=( _mesh_1_1_io_out_last_0) ^ ((fiEnable && (8243 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3107_0 <=( _mesh_2_1_io_out_last_0) ^ ((fiEnable && (8244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3108_0 <=( _mesh_3_1_io_out_last_0) ^ ((fiEnable && (8245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3109_0 <=( _mesh_4_1_io_out_last_0) ^ ((fiEnable && (8246 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3110_0 <=( _mesh_5_1_io_out_last_0) ^ ((fiEnable && (8247 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3111_0 <=( _mesh_6_1_io_out_last_0) ^ ((fiEnable && (8248 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3112_0 <=( _mesh_7_1_io_out_last_0) ^ ((fiEnable && (8249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3113_0 <=( _mesh_8_1_io_out_last_0) ^ ((fiEnable && (8250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3114_0 <=( _mesh_9_1_io_out_last_0) ^ ((fiEnable && (8251 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3115_0 <=( _mesh_10_1_io_out_last_0) ^ ((fiEnable && (8252 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3116_0 <=( _mesh_11_1_io_out_last_0) ^ ((fiEnable && (8253 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3117_0 <=( _mesh_12_1_io_out_last_0) ^ ((fiEnable && (8254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3118_0 <=( _mesh_13_1_io_out_last_0) ^ ((fiEnable && (8255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3119_0 <=( _mesh_14_1_io_out_last_0) ^ ((fiEnable && (8256 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3120_0 <=( _mesh_15_1_io_out_last_0) ^ ((fiEnable && (8257 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3121_0 <=( _mesh_16_1_io_out_last_0) ^ ((fiEnable && (8258 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3122_0 <=( _mesh_17_1_io_out_last_0) ^ ((fiEnable && (8259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3123_0 <=( _mesh_18_1_io_out_last_0) ^ ((fiEnable && (8260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3124_0 <=( _mesh_19_1_io_out_last_0) ^ ((fiEnable && (8261 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3125_0 <=( _mesh_20_1_io_out_last_0) ^ ((fiEnable && (8262 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3126_0 <=( _mesh_21_1_io_out_last_0) ^ ((fiEnable && (8263 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3127_0 <=( _mesh_22_1_io_out_last_0) ^ ((fiEnable && (8264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3128_0 <=( _mesh_23_1_io_out_last_0) ^ ((fiEnable && (8265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3129_0 <=( _mesh_24_1_io_out_last_0) ^ ((fiEnable && (8266 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3130_0 <=( _mesh_25_1_io_out_last_0) ^ ((fiEnable && (8267 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3131_0 <=( _mesh_26_1_io_out_last_0) ^ ((fiEnable && (8268 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3132_0 <=( _mesh_27_1_io_out_last_0) ^ ((fiEnable && (8269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3133_0 <=( _mesh_28_1_io_out_last_0) ^ ((fiEnable && (8270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3134_0 <=( _mesh_29_1_io_out_last_0) ^ ((fiEnable && (8271 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3135_0 <=( _mesh_30_1_io_out_last_0) ^ ((fiEnable && (8272 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3136_0 <=( io_in_last_2_0) ^ ((fiEnable && (8273 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3137_0 <=( _mesh_0_2_io_out_last_0) ^ ((fiEnable && (8274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3138_0 <=( _mesh_1_2_io_out_last_0) ^ ((fiEnable && (8275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3139_0 <=( _mesh_2_2_io_out_last_0) ^ ((fiEnable && (8276 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3140_0 <=( _mesh_3_2_io_out_last_0) ^ ((fiEnable && (8277 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3141_0 <=( _mesh_4_2_io_out_last_0) ^ ((fiEnable && (8278 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3142_0 <=( _mesh_5_2_io_out_last_0) ^ ((fiEnable && (8279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3143_0 <=( _mesh_6_2_io_out_last_0) ^ ((fiEnable && (8280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3144_0 <=( _mesh_7_2_io_out_last_0) ^ ((fiEnable && (8281 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3145_0 <=( _mesh_8_2_io_out_last_0) ^ ((fiEnable && (8282 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3146_0 <=( _mesh_9_2_io_out_last_0) ^ ((fiEnable && (8283 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3147_0 <=( _mesh_10_2_io_out_last_0) ^ ((fiEnable && (8284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3148_0 <=( _mesh_11_2_io_out_last_0) ^ ((fiEnable && (8285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3149_0 <=( _mesh_12_2_io_out_last_0) ^ ((fiEnable && (8286 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3150_0 <=( _mesh_13_2_io_out_last_0) ^ ((fiEnable && (8287 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3151_0 <=( _mesh_14_2_io_out_last_0) ^ ((fiEnable && (8288 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3152_0 <=( _mesh_15_2_io_out_last_0) ^ ((fiEnable && (8289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3153_0 <=( _mesh_16_2_io_out_last_0) ^ ((fiEnable && (8290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3154_0 <=( _mesh_17_2_io_out_last_0) ^ ((fiEnable && (8291 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3155_0 <=( _mesh_18_2_io_out_last_0) ^ ((fiEnable && (8292 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3156_0 <=( _mesh_19_2_io_out_last_0) ^ ((fiEnable && (8293 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3157_0 <=( _mesh_20_2_io_out_last_0) ^ ((fiEnable && (8294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3158_0 <=( _mesh_21_2_io_out_last_0) ^ ((fiEnable && (8295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3159_0 <=( _mesh_22_2_io_out_last_0) ^ ((fiEnable && (8296 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3160_0 <=( _mesh_23_2_io_out_last_0) ^ ((fiEnable && (8297 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3161_0 <=( _mesh_24_2_io_out_last_0) ^ ((fiEnable && (8298 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3162_0 <=( _mesh_25_2_io_out_last_0) ^ ((fiEnable && (8299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3163_0 <=( _mesh_26_2_io_out_last_0) ^ ((fiEnable && (8300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3164_0 <=( _mesh_27_2_io_out_last_0) ^ ((fiEnable && (8301 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3165_0 <=( _mesh_28_2_io_out_last_0) ^ ((fiEnable && (8302 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3166_0 <=( _mesh_29_2_io_out_last_0) ^ ((fiEnable && (8303 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3167_0 <=( _mesh_30_2_io_out_last_0) ^ ((fiEnable && (8304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3168_0 <=( io_in_last_3_0) ^ ((fiEnable && (8305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3169_0 <=( _mesh_0_3_io_out_last_0) ^ ((fiEnable && (8306 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3170_0 <=( _mesh_1_3_io_out_last_0) ^ ((fiEnable && (8307 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3171_0 <=( _mesh_2_3_io_out_last_0) ^ ((fiEnable && (8308 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3172_0 <=( _mesh_3_3_io_out_last_0) ^ ((fiEnable && (8309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3173_0 <=( _mesh_4_3_io_out_last_0) ^ ((fiEnable && (8310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3174_0 <=( _mesh_5_3_io_out_last_0) ^ ((fiEnable && (8311 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3175_0 <=( _mesh_6_3_io_out_last_0) ^ ((fiEnable && (8312 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3176_0 <=( _mesh_7_3_io_out_last_0) ^ ((fiEnable && (8313 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3177_0 <=( _mesh_8_3_io_out_last_0) ^ ((fiEnable && (8314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3178_0 <=( _mesh_9_3_io_out_last_0) ^ ((fiEnable && (8315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3179_0 <=( _mesh_10_3_io_out_last_0) ^ ((fiEnable && (8316 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3180_0 <=( _mesh_11_3_io_out_last_0) ^ ((fiEnable && (8317 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3181_0 <=( _mesh_12_3_io_out_last_0) ^ ((fiEnable && (8318 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3182_0 <=( _mesh_13_3_io_out_last_0) ^ ((fiEnable && (8319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3183_0 <=( _mesh_14_3_io_out_last_0) ^ ((fiEnable && (8320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3184_0 <=( _mesh_15_3_io_out_last_0) ^ ((fiEnable && (8321 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3185_0 <=( _mesh_16_3_io_out_last_0) ^ ((fiEnable && (8322 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3186_0 <=( _mesh_17_3_io_out_last_0) ^ ((fiEnable && (8323 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3187_0 <=( _mesh_18_3_io_out_last_0) ^ ((fiEnable && (8324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3188_0 <=( _mesh_19_3_io_out_last_0) ^ ((fiEnable && (8325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3189_0 <=( _mesh_20_3_io_out_last_0) ^ ((fiEnable && (8326 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3190_0 <=( _mesh_21_3_io_out_last_0) ^ ((fiEnable && (8327 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3191_0 <=( _mesh_22_3_io_out_last_0) ^ ((fiEnable && (8328 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3192_0 <=( _mesh_23_3_io_out_last_0) ^ ((fiEnable && (8329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3193_0 <=( _mesh_24_3_io_out_last_0) ^ ((fiEnable && (8330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3194_0 <=( _mesh_25_3_io_out_last_0) ^ ((fiEnable && (8331 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3195_0 <=( _mesh_26_3_io_out_last_0) ^ ((fiEnable && (8332 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3196_0 <=( _mesh_27_3_io_out_last_0) ^ ((fiEnable && (8333 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3197_0 <=( _mesh_28_3_io_out_last_0) ^ ((fiEnable && (8334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3198_0 <=( _mesh_29_3_io_out_last_0) ^ ((fiEnable && (8335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3199_0 <=( _mesh_30_3_io_out_last_0) ^ ((fiEnable && (8336 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3200_0 <=( io_in_last_4_0) ^ ((fiEnable && (8337 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3201_0 <=( _mesh_0_4_io_out_last_0) ^ ((fiEnable && (8338 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3202_0 <=( _mesh_1_4_io_out_last_0) ^ ((fiEnable && (8339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3203_0 <=( _mesh_2_4_io_out_last_0) ^ ((fiEnable && (8340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3204_0 <=( _mesh_3_4_io_out_last_0) ^ ((fiEnable && (8341 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3205_0 <=( _mesh_4_4_io_out_last_0) ^ ((fiEnable && (8342 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3206_0 <=( _mesh_5_4_io_out_last_0) ^ ((fiEnable && (8343 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3207_0 <=( _mesh_6_4_io_out_last_0) ^ ((fiEnable && (8344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3208_0 <=( _mesh_7_4_io_out_last_0) ^ ((fiEnable && (8345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3209_0 <=( _mesh_8_4_io_out_last_0) ^ ((fiEnable && (8346 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3210_0 <=( _mesh_9_4_io_out_last_0) ^ ((fiEnable && (8347 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3211_0 <=( _mesh_10_4_io_out_last_0) ^ ((fiEnable && (8348 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3212_0 <=( _mesh_11_4_io_out_last_0) ^ ((fiEnable && (8349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3213_0 <=( _mesh_12_4_io_out_last_0) ^ ((fiEnable && (8350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3214_0 <=( _mesh_13_4_io_out_last_0) ^ ((fiEnable && (8351 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3215_0 <=( _mesh_14_4_io_out_last_0) ^ ((fiEnable && (8352 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3216_0 <=( _mesh_15_4_io_out_last_0) ^ ((fiEnable && (8353 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3217_0 <=( _mesh_16_4_io_out_last_0) ^ ((fiEnable && (8354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3218_0 <=( _mesh_17_4_io_out_last_0) ^ ((fiEnable && (8355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3219_0 <=( _mesh_18_4_io_out_last_0) ^ ((fiEnable && (8356 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3220_0 <=( _mesh_19_4_io_out_last_0) ^ ((fiEnable && (8357 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3221_0 <=( _mesh_20_4_io_out_last_0) ^ ((fiEnable && (8358 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3222_0 <=( _mesh_21_4_io_out_last_0) ^ ((fiEnable && (8359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3223_0 <=( _mesh_22_4_io_out_last_0) ^ ((fiEnable && (8360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3224_0 <=( _mesh_23_4_io_out_last_0) ^ ((fiEnable && (8361 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3225_0 <=( _mesh_24_4_io_out_last_0) ^ ((fiEnable && (8362 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3226_0 <=( _mesh_25_4_io_out_last_0) ^ ((fiEnable && (8363 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3227_0 <=( _mesh_26_4_io_out_last_0) ^ ((fiEnable && (8364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3228_0 <=( _mesh_27_4_io_out_last_0) ^ ((fiEnable && (8365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3229_0 <=( _mesh_28_4_io_out_last_0) ^ ((fiEnable && (8366 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3230_0 <=( _mesh_29_4_io_out_last_0) ^ ((fiEnable && (8367 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3231_0 <=( _mesh_30_4_io_out_last_0) ^ ((fiEnable && (8368 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3232_0 <=( io_in_last_5_0) ^ ((fiEnable && (8369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3233_0 <=( _mesh_0_5_io_out_last_0) ^ ((fiEnable && (8370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3234_0 <=( _mesh_1_5_io_out_last_0) ^ ((fiEnable && (8371 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3235_0 <=( _mesh_2_5_io_out_last_0) ^ ((fiEnable && (8372 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3236_0 <=( _mesh_3_5_io_out_last_0) ^ ((fiEnable && (8373 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3237_0 <=( _mesh_4_5_io_out_last_0) ^ ((fiEnable && (8374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3238_0 <=( _mesh_5_5_io_out_last_0) ^ ((fiEnable && (8375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3239_0 <=( _mesh_6_5_io_out_last_0) ^ ((fiEnable && (8376 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3240_0 <=( _mesh_7_5_io_out_last_0) ^ ((fiEnable && (8377 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3241_0 <=( _mesh_8_5_io_out_last_0) ^ ((fiEnable && (8378 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3242_0 <=( _mesh_9_5_io_out_last_0) ^ ((fiEnable && (8379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3243_0 <=( _mesh_10_5_io_out_last_0) ^ ((fiEnable && (8380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3244_0 <=( _mesh_11_5_io_out_last_0) ^ ((fiEnable && (8381 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3245_0 <=( _mesh_12_5_io_out_last_0) ^ ((fiEnable && (8382 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3246_0 <=( _mesh_13_5_io_out_last_0) ^ ((fiEnable && (8383 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3247_0 <=( _mesh_14_5_io_out_last_0) ^ ((fiEnable && (8384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3248_0 <=( _mesh_15_5_io_out_last_0) ^ ((fiEnable && (8385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3249_0 <=( _mesh_16_5_io_out_last_0) ^ ((fiEnable && (8386 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3250_0 <=( _mesh_17_5_io_out_last_0) ^ ((fiEnable && (8387 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3251_0 <=( _mesh_18_5_io_out_last_0) ^ ((fiEnable && (8388 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3252_0 <=( _mesh_19_5_io_out_last_0) ^ ((fiEnable && (8389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3253_0 <=( _mesh_20_5_io_out_last_0) ^ ((fiEnable && (8390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3254_0 <=( _mesh_21_5_io_out_last_0) ^ ((fiEnable && (8391 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3255_0 <=( _mesh_22_5_io_out_last_0) ^ ((fiEnable && (8392 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3256_0 <=( _mesh_23_5_io_out_last_0) ^ ((fiEnable && (8393 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3257_0 <=( _mesh_24_5_io_out_last_0) ^ ((fiEnable && (8394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3258_0 <=( _mesh_25_5_io_out_last_0) ^ ((fiEnable && (8395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3259_0 <=( _mesh_26_5_io_out_last_0) ^ ((fiEnable && (8396 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3260_0 <=( _mesh_27_5_io_out_last_0) ^ ((fiEnable && (8397 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3261_0 <=( _mesh_28_5_io_out_last_0) ^ ((fiEnable && (8398 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3262_0 <=( _mesh_29_5_io_out_last_0) ^ ((fiEnable && (8399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3263_0 <=( _mesh_30_5_io_out_last_0) ^ ((fiEnable && (8400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3264_0 <=( io_in_last_6_0) ^ ((fiEnable && (8401 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3265_0 <=( _mesh_0_6_io_out_last_0) ^ ((fiEnable && (8402 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3266_0 <=( _mesh_1_6_io_out_last_0) ^ ((fiEnable && (8403 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3267_0 <=( _mesh_2_6_io_out_last_0) ^ ((fiEnable && (8404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3268_0 <=( _mesh_3_6_io_out_last_0) ^ ((fiEnable && (8405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3269_0 <=( _mesh_4_6_io_out_last_0) ^ ((fiEnable && (8406 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3270_0 <=( _mesh_5_6_io_out_last_0) ^ ((fiEnable && (8407 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3271_0 <=( _mesh_6_6_io_out_last_0) ^ ((fiEnable && (8408 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3272_0 <=( _mesh_7_6_io_out_last_0) ^ ((fiEnable && (8409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3273_0 <=( _mesh_8_6_io_out_last_0) ^ ((fiEnable && (8410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3274_0 <=( _mesh_9_6_io_out_last_0) ^ ((fiEnable && (8411 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3275_0 <=( _mesh_10_6_io_out_last_0) ^ ((fiEnable && (8412 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3276_0 <=( _mesh_11_6_io_out_last_0) ^ ((fiEnable && (8413 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3277_0 <=( _mesh_12_6_io_out_last_0) ^ ((fiEnable && (8414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3278_0 <=( _mesh_13_6_io_out_last_0) ^ ((fiEnable && (8415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3279_0 <=( _mesh_14_6_io_out_last_0) ^ ((fiEnable && (8416 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3280_0 <=( _mesh_15_6_io_out_last_0) ^ ((fiEnable && (8417 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3281_0 <=( _mesh_16_6_io_out_last_0) ^ ((fiEnable && (8418 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3282_0 <=( _mesh_17_6_io_out_last_0) ^ ((fiEnable && (8419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3283_0 <=( _mesh_18_6_io_out_last_0) ^ ((fiEnable && (8420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3284_0 <=( _mesh_19_6_io_out_last_0) ^ ((fiEnable && (8421 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3285_0 <=( _mesh_20_6_io_out_last_0) ^ ((fiEnable && (8422 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3286_0 <=( _mesh_21_6_io_out_last_0) ^ ((fiEnable && (8423 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3287_0 <=( _mesh_22_6_io_out_last_0) ^ ((fiEnable && (8424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3288_0 <=( _mesh_23_6_io_out_last_0) ^ ((fiEnable && (8425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3289_0 <=( _mesh_24_6_io_out_last_0) ^ ((fiEnable && (8426 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3290_0 <=( _mesh_25_6_io_out_last_0) ^ ((fiEnable && (8427 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3291_0 <=( _mesh_26_6_io_out_last_0) ^ ((fiEnable && (8428 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3292_0 <=( _mesh_27_6_io_out_last_0) ^ ((fiEnable && (8429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3293_0 <=( _mesh_28_6_io_out_last_0) ^ ((fiEnable && (8430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3294_0 <=( _mesh_29_6_io_out_last_0) ^ ((fiEnable && (8431 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3295_0 <=( _mesh_30_6_io_out_last_0) ^ ((fiEnable && (8432 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3296_0 <=( io_in_last_7_0) ^ ((fiEnable && (8433 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3297_0 <=( _mesh_0_7_io_out_last_0) ^ ((fiEnable && (8434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3298_0 <=( _mesh_1_7_io_out_last_0) ^ ((fiEnable && (8435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3299_0 <=( _mesh_2_7_io_out_last_0) ^ ((fiEnable && (8436 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3300_0 <=( _mesh_3_7_io_out_last_0) ^ ((fiEnable && (8437 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3301_0 <=( _mesh_4_7_io_out_last_0) ^ ((fiEnable && (8438 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3302_0 <=( _mesh_5_7_io_out_last_0) ^ ((fiEnable && (8439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3303_0 <=( _mesh_6_7_io_out_last_0) ^ ((fiEnable && (8440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3304_0 <=( _mesh_7_7_io_out_last_0) ^ ((fiEnable && (8441 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3305_0 <=( _mesh_8_7_io_out_last_0) ^ ((fiEnable && (8442 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3306_0 <=( _mesh_9_7_io_out_last_0) ^ ((fiEnable && (8443 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3307_0 <=( _mesh_10_7_io_out_last_0) ^ ((fiEnable && (8444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3308_0 <=( _mesh_11_7_io_out_last_0) ^ ((fiEnable && (8445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3309_0 <=( _mesh_12_7_io_out_last_0) ^ ((fiEnable && (8446 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3310_0 <=( _mesh_13_7_io_out_last_0) ^ ((fiEnable && (8447 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3311_0 <=( _mesh_14_7_io_out_last_0) ^ ((fiEnable && (8448 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3312_0 <=( _mesh_15_7_io_out_last_0) ^ ((fiEnable && (8449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3313_0 <=( _mesh_16_7_io_out_last_0) ^ ((fiEnable && (8450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3314_0 <=( _mesh_17_7_io_out_last_0) ^ ((fiEnable && (8451 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3315_0 <=( _mesh_18_7_io_out_last_0) ^ ((fiEnable && (8452 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3316_0 <=( _mesh_19_7_io_out_last_0) ^ ((fiEnable && (8453 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3317_0 <=( _mesh_20_7_io_out_last_0) ^ ((fiEnable && (8454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3318_0 <=( _mesh_21_7_io_out_last_0) ^ ((fiEnable && (8455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3319_0 <=( _mesh_22_7_io_out_last_0) ^ ((fiEnable && (8456 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3320_0 <=( _mesh_23_7_io_out_last_0) ^ ((fiEnable && (8457 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3321_0 <=( _mesh_24_7_io_out_last_0) ^ ((fiEnable && (8458 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3322_0 <=( _mesh_25_7_io_out_last_0) ^ ((fiEnable && (8459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3323_0 <=( _mesh_26_7_io_out_last_0) ^ ((fiEnable && (8460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3324_0 <=( _mesh_27_7_io_out_last_0) ^ ((fiEnable && (8461 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3325_0 <=( _mesh_28_7_io_out_last_0) ^ ((fiEnable && (8462 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3326_0 <=( _mesh_29_7_io_out_last_0) ^ ((fiEnable && (8463 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3327_0 <=( _mesh_30_7_io_out_last_0) ^ ((fiEnable && (8464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3328_0 <=( io_in_last_8_0) ^ ((fiEnable && (8465 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3329_0 <=( _mesh_0_8_io_out_last_0) ^ ((fiEnable && (8466 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3330_0 <=( _mesh_1_8_io_out_last_0) ^ ((fiEnable && (8467 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3331_0 <=( _mesh_2_8_io_out_last_0) ^ ((fiEnable && (8468 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3332_0 <=( _mesh_3_8_io_out_last_0) ^ ((fiEnable && (8469 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3333_0 <=( _mesh_4_8_io_out_last_0) ^ ((fiEnable && (8470 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3334_0 <=( _mesh_5_8_io_out_last_0) ^ ((fiEnable && (8471 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3335_0 <=( _mesh_6_8_io_out_last_0) ^ ((fiEnable && (8472 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3336_0 <=( _mesh_7_8_io_out_last_0) ^ ((fiEnable && (8473 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3337_0 <=( _mesh_8_8_io_out_last_0) ^ ((fiEnable && (8474 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3338_0 <=( _mesh_9_8_io_out_last_0) ^ ((fiEnable && (8475 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3339_0 <=( _mesh_10_8_io_out_last_0) ^ ((fiEnable && (8476 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3340_0 <=( _mesh_11_8_io_out_last_0) ^ ((fiEnable && (8477 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3341_0 <=( _mesh_12_8_io_out_last_0) ^ ((fiEnable && (8478 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3342_0 <=( _mesh_13_8_io_out_last_0) ^ ((fiEnable && (8479 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3343_0 <=( _mesh_14_8_io_out_last_0) ^ ((fiEnable && (8480 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3344_0 <=( _mesh_15_8_io_out_last_0) ^ ((fiEnable && (8481 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3345_0 <=( _mesh_16_8_io_out_last_0) ^ ((fiEnable && (8482 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3346_0 <=( _mesh_17_8_io_out_last_0) ^ ((fiEnable && (8483 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3347_0 <=( _mesh_18_8_io_out_last_0) ^ ((fiEnable && (8484 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3348_0 <=( _mesh_19_8_io_out_last_0) ^ ((fiEnable && (8485 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3349_0 <=( _mesh_20_8_io_out_last_0) ^ ((fiEnable && (8486 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3350_0 <=( _mesh_21_8_io_out_last_0) ^ ((fiEnable && (8487 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3351_0 <=( _mesh_22_8_io_out_last_0) ^ ((fiEnable && (8488 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3352_0 <=( _mesh_23_8_io_out_last_0) ^ ((fiEnable && (8489 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3353_0 <=( _mesh_24_8_io_out_last_0) ^ ((fiEnable && (8490 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3354_0 <=( _mesh_25_8_io_out_last_0) ^ ((fiEnable && (8491 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3355_0 <=( _mesh_26_8_io_out_last_0) ^ ((fiEnable && (8492 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3356_0 <=( _mesh_27_8_io_out_last_0) ^ ((fiEnable && (8493 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3357_0 <=( _mesh_28_8_io_out_last_0) ^ ((fiEnable && (8494 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3358_0 <=( _mesh_29_8_io_out_last_0) ^ ((fiEnable && (8495 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3359_0 <=( _mesh_30_8_io_out_last_0) ^ ((fiEnable && (8496 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3360_0 <=( io_in_last_9_0) ^ ((fiEnable && (8497 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3361_0 <=( _mesh_0_9_io_out_last_0) ^ ((fiEnable && (8498 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3362_0 <=( _mesh_1_9_io_out_last_0) ^ ((fiEnable && (8499 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3363_0 <=( _mesh_2_9_io_out_last_0) ^ ((fiEnable && (8500 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3364_0 <=( _mesh_3_9_io_out_last_0) ^ ((fiEnable && (8501 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3365_0 <=( _mesh_4_9_io_out_last_0) ^ ((fiEnable && (8502 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3366_0 <=( _mesh_5_9_io_out_last_0) ^ ((fiEnable && (8503 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3367_0 <=( _mesh_6_9_io_out_last_0) ^ ((fiEnable && (8504 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3368_0 <=( _mesh_7_9_io_out_last_0) ^ ((fiEnable && (8505 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3369_0 <=( _mesh_8_9_io_out_last_0) ^ ((fiEnable && (8506 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3370_0 <=( _mesh_9_9_io_out_last_0) ^ ((fiEnable && (8507 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3371_0 <=( _mesh_10_9_io_out_last_0) ^ ((fiEnable && (8508 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3372_0 <=( _mesh_11_9_io_out_last_0) ^ ((fiEnable && (8509 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3373_0 <=( _mesh_12_9_io_out_last_0) ^ ((fiEnable && (8510 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3374_0 <=( _mesh_13_9_io_out_last_0) ^ ((fiEnable && (8511 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3375_0 <=( _mesh_14_9_io_out_last_0) ^ ((fiEnable && (8512 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3376_0 <=( _mesh_15_9_io_out_last_0) ^ ((fiEnable && (8513 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3377_0 <=( _mesh_16_9_io_out_last_0) ^ ((fiEnable && (8514 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3378_0 <=( _mesh_17_9_io_out_last_0) ^ ((fiEnable && (8515 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3379_0 <=( _mesh_18_9_io_out_last_0) ^ ((fiEnable && (8516 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3380_0 <=( _mesh_19_9_io_out_last_0) ^ ((fiEnable && (8517 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3381_0 <=( _mesh_20_9_io_out_last_0) ^ ((fiEnable && (8518 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3382_0 <=( _mesh_21_9_io_out_last_0) ^ ((fiEnable && (8519 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3383_0 <=( _mesh_22_9_io_out_last_0) ^ ((fiEnable && (8520 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3384_0 <=( _mesh_23_9_io_out_last_0) ^ ((fiEnable && (8521 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3385_0 <=( _mesh_24_9_io_out_last_0) ^ ((fiEnable && (8522 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3386_0 <=( _mesh_25_9_io_out_last_0) ^ ((fiEnable && (8523 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3387_0 <=( _mesh_26_9_io_out_last_0) ^ ((fiEnable && (8524 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3388_0 <=( _mesh_27_9_io_out_last_0) ^ ((fiEnable && (8525 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3389_0 <=( _mesh_28_9_io_out_last_0) ^ ((fiEnable && (8526 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3390_0 <=( _mesh_29_9_io_out_last_0) ^ ((fiEnable && (8527 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3391_0 <=( _mesh_30_9_io_out_last_0) ^ ((fiEnable && (8528 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3392_0 <=( io_in_last_10_0) ^ ((fiEnable && (8529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3393_0 <=( _mesh_0_10_io_out_last_0) ^ ((fiEnable && (8530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3394_0 <=( _mesh_1_10_io_out_last_0) ^ ((fiEnable && (8531 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3395_0 <=( _mesh_2_10_io_out_last_0) ^ ((fiEnable && (8532 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3396_0 <=( _mesh_3_10_io_out_last_0) ^ ((fiEnable && (8533 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3397_0 <=( _mesh_4_10_io_out_last_0) ^ ((fiEnable && (8534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3398_0 <=( _mesh_5_10_io_out_last_0) ^ ((fiEnable && (8535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3399_0 <=( _mesh_6_10_io_out_last_0) ^ ((fiEnable && (8536 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3400_0 <=( _mesh_7_10_io_out_last_0) ^ ((fiEnable && (8537 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3401_0 <=( _mesh_8_10_io_out_last_0) ^ ((fiEnable && (8538 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3402_0 <=( _mesh_9_10_io_out_last_0) ^ ((fiEnable && (8539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3403_0 <=( _mesh_10_10_io_out_last_0) ^ ((fiEnable && (8540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3404_0 <=( _mesh_11_10_io_out_last_0) ^ ((fiEnable && (8541 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3405_0 <=( _mesh_12_10_io_out_last_0) ^ ((fiEnable && (8542 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3406_0 <=( _mesh_13_10_io_out_last_0) ^ ((fiEnable && (8543 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3407_0 <=( _mesh_14_10_io_out_last_0) ^ ((fiEnable && (8544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3408_0 <=( _mesh_15_10_io_out_last_0) ^ ((fiEnable && (8545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3409_0 <=( _mesh_16_10_io_out_last_0) ^ ((fiEnable && (8546 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3410_0 <=( _mesh_17_10_io_out_last_0) ^ ((fiEnable && (8547 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3411_0 <=( _mesh_18_10_io_out_last_0) ^ ((fiEnable && (8548 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3412_0 <=( _mesh_19_10_io_out_last_0) ^ ((fiEnable && (8549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3413_0 <=( _mesh_20_10_io_out_last_0) ^ ((fiEnable && (8550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3414_0 <=( _mesh_21_10_io_out_last_0) ^ ((fiEnable && (8551 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3415_0 <=( _mesh_22_10_io_out_last_0) ^ ((fiEnable && (8552 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3416_0 <=( _mesh_23_10_io_out_last_0) ^ ((fiEnable && (8553 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3417_0 <=( _mesh_24_10_io_out_last_0) ^ ((fiEnable && (8554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3418_0 <=( _mesh_25_10_io_out_last_0) ^ ((fiEnable && (8555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3419_0 <=( _mesh_26_10_io_out_last_0) ^ ((fiEnable && (8556 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3420_0 <=( _mesh_27_10_io_out_last_0) ^ ((fiEnable && (8557 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3421_0 <=( _mesh_28_10_io_out_last_0) ^ ((fiEnable && (8558 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3422_0 <=( _mesh_29_10_io_out_last_0) ^ ((fiEnable && (8559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3423_0 <=( _mesh_30_10_io_out_last_0) ^ ((fiEnable && (8560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3424_0 <=( io_in_last_11_0) ^ ((fiEnable && (8561 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3425_0 <=( _mesh_0_11_io_out_last_0) ^ ((fiEnable && (8562 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3426_0 <=( _mesh_1_11_io_out_last_0) ^ ((fiEnable && (8563 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3427_0 <=( _mesh_2_11_io_out_last_0) ^ ((fiEnable && (8564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3428_0 <=( _mesh_3_11_io_out_last_0) ^ ((fiEnable && (8565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3429_0 <=( _mesh_4_11_io_out_last_0) ^ ((fiEnable && (8566 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3430_0 <=( _mesh_5_11_io_out_last_0) ^ ((fiEnable && (8567 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3431_0 <=( _mesh_6_11_io_out_last_0) ^ ((fiEnable && (8568 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3432_0 <=( _mesh_7_11_io_out_last_0) ^ ((fiEnable && (8569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3433_0 <=( _mesh_8_11_io_out_last_0) ^ ((fiEnable && (8570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3434_0 <=( _mesh_9_11_io_out_last_0) ^ ((fiEnable && (8571 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3435_0 <=( _mesh_10_11_io_out_last_0) ^ ((fiEnable && (8572 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3436_0 <=( _mesh_11_11_io_out_last_0) ^ ((fiEnable && (8573 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3437_0 <=( _mesh_12_11_io_out_last_0) ^ ((fiEnable && (8574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3438_0 <=( _mesh_13_11_io_out_last_0) ^ ((fiEnable && (8575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3439_0 <=( _mesh_14_11_io_out_last_0) ^ ((fiEnable && (8576 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3440_0 <=( _mesh_15_11_io_out_last_0) ^ ((fiEnable && (8577 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3441_0 <=( _mesh_16_11_io_out_last_0) ^ ((fiEnable && (8578 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3442_0 <=( _mesh_17_11_io_out_last_0) ^ ((fiEnable && (8579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3443_0 <=( _mesh_18_11_io_out_last_0) ^ ((fiEnable && (8580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3444_0 <=( _mesh_19_11_io_out_last_0) ^ ((fiEnable && (8581 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3445_0 <=( _mesh_20_11_io_out_last_0) ^ ((fiEnable && (8582 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3446_0 <=( _mesh_21_11_io_out_last_0) ^ ((fiEnable && (8583 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3447_0 <=( _mesh_22_11_io_out_last_0) ^ ((fiEnable && (8584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3448_0 <=( _mesh_23_11_io_out_last_0) ^ ((fiEnable && (8585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3449_0 <=( _mesh_24_11_io_out_last_0) ^ ((fiEnable && (8586 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3450_0 <=( _mesh_25_11_io_out_last_0) ^ ((fiEnable && (8587 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3451_0 <=( _mesh_26_11_io_out_last_0) ^ ((fiEnable && (8588 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3452_0 <=( _mesh_27_11_io_out_last_0) ^ ((fiEnable && (8589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3453_0 <=( _mesh_28_11_io_out_last_0) ^ ((fiEnable && (8590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3454_0 <=( _mesh_29_11_io_out_last_0) ^ ((fiEnable && (8591 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3455_0 <=( _mesh_30_11_io_out_last_0) ^ ((fiEnable && (8592 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3456_0 <=( io_in_last_12_0) ^ ((fiEnable && (8593 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3457_0 <=( _mesh_0_12_io_out_last_0) ^ ((fiEnable && (8594 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3458_0 <=( _mesh_1_12_io_out_last_0) ^ ((fiEnable && (8595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3459_0 <=( _mesh_2_12_io_out_last_0) ^ ((fiEnable && (8596 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3460_0 <=( _mesh_3_12_io_out_last_0) ^ ((fiEnable && (8597 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3461_0 <=( _mesh_4_12_io_out_last_0) ^ ((fiEnable && (8598 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3462_0 <=( _mesh_5_12_io_out_last_0) ^ ((fiEnable && (8599 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3463_0 <=( _mesh_6_12_io_out_last_0) ^ ((fiEnable && (8600 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3464_0 <=( _mesh_7_12_io_out_last_0) ^ ((fiEnable && (8601 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3465_0 <=( _mesh_8_12_io_out_last_0) ^ ((fiEnable && (8602 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3466_0 <=( _mesh_9_12_io_out_last_0) ^ ((fiEnable && (8603 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3467_0 <=( _mesh_10_12_io_out_last_0) ^ ((fiEnable && (8604 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3468_0 <=( _mesh_11_12_io_out_last_0) ^ ((fiEnable && (8605 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3469_0 <=( _mesh_12_12_io_out_last_0) ^ ((fiEnable && (8606 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3470_0 <=( _mesh_13_12_io_out_last_0) ^ ((fiEnable && (8607 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3471_0 <=( _mesh_14_12_io_out_last_0) ^ ((fiEnable && (8608 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3472_0 <=( _mesh_15_12_io_out_last_0) ^ ((fiEnable && (8609 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3473_0 <=( _mesh_16_12_io_out_last_0) ^ ((fiEnable && (8610 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3474_0 <=( _mesh_17_12_io_out_last_0) ^ ((fiEnable && (8611 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3475_0 <=( _mesh_18_12_io_out_last_0) ^ ((fiEnable && (8612 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3476_0 <=( _mesh_19_12_io_out_last_0) ^ ((fiEnable && (8613 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3477_0 <=( _mesh_20_12_io_out_last_0) ^ ((fiEnable && (8614 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3478_0 <=( _mesh_21_12_io_out_last_0) ^ ((fiEnable && (8615 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3479_0 <=( _mesh_22_12_io_out_last_0) ^ ((fiEnable && (8616 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3480_0 <=( _mesh_23_12_io_out_last_0) ^ ((fiEnable && (8617 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3481_0 <=( _mesh_24_12_io_out_last_0) ^ ((fiEnable && (8618 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3482_0 <=( _mesh_25_12_io_out_last_0) ^ ((fiEnable && (8619 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3483_0 <=( _mesh_26_12_io_out_last_0) ^ ((fiEnable && (8620 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3484_0 <=( _mesh_27_12_io_out_last_0) ^ ((fiEnable && (8621 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3485_0 <=( _mesh_28_12_io_out_last_0) ^ ((fiEnable && (8622 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3486_0 <=( _mesh_29_12_io_out_last_0) ^ ((fiEnable && (8623 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3487_0 <=( _mesh_30_12_io_out_last_0) ^ ((fiEnable && (8624 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3488_0 <=( io_in_last_13_0) ^ ((fiEnable && (8625 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3489_0 <=( _mesh_0_13_io_out_last_0) ^ ((fiEnable && (8626 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3490_0 <=( _mesh_1_13_io_out_last_0) ^ ((fiEnable && (8627 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3491_0 <=( _mesh_2_13_io_out_last_0) ^ ((fiEnable && (8628 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3492_0 <=( _mesh_3_13_io_out_last_0) ^ ((fiEnable && (8629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3493_0 <=( _mesh_4_13_io_out_last_0) ^ ((fiEnable && (8630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3494_0 <=( _mesh_5_13_io_out_last_0) ^ ((fiEnable && (8631 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3495_0 <=( _mesh_6_13_io_out_last_0) ^ ((fiEnable && (8632 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3496_0 <=( _mesh_7_13_io_out_last_0) ^ ((fiEnable && (8633 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3497_0 <=( _mesh_8_13_io_out_last_0) ^ ((fiEnable && (8634 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3498_0 <=( _mesh_9_13_io_out_last_0) ^ ((fiEnable && (8635 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3499_0 <=( _mesh_10_13_io_out_last_0) ^ ((fiEnable && (8636 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3500_0 <=( _mesh_11_13_io_out_last_0) ^ ((fiEnable && (8637 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3501_0 <=( _mesh_12_13_io_out_last_0) ^ ((fiEnable && (8638 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3502_0 <=( _mesh_13_13_io_out_last_0) ^ ((fiEnable && (8639 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3503_0 <=( _mesh_14_13_io_out_last_0) ^ ((fiEnable && (8640 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3504_0 <=( _mesh_15_13_io_out_last_0) ^ ((fiEnable && (8641 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3505_0 <=( _mesh_16_13_io_out_last_0) ^ ((fiEnable && (8642 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3506_0 <=( _mesh_17_13_io_out_last_0) ^ ((fiEnable && (8643 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3507_0 <=( _mesh_18_13_io_out_last_0) ^ ((fiEnable && (8644 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3508_0 <=( _mesh_19_13_io_out_last_0) ^ ((fiEnable && (8645 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3509_0 <=( _mesh_20_13_io_out_last_0) ^ ((fiEnable && (8646 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3510_0 <=( _mesh_21_13_io_out_last_0) ^ ((fiEnable && (8647 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3511_0 <=( _mesh_22_13_io_out_last_0) ^ ((fiEnable && (8648 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3512_0 <=( _mesh_23_13_io_out_last_0) ^ ((fiEnable && (8649 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3513_0 <=( _mesh_24_13_io_out_last_0) ^ ((fiEnable && (8650 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3514_0 <=( _mesh_25_13_io_out_last_0) ^ ((fiEnable && (8651 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3515_0 <=( _mesh_26_13_io_out_last_0) ^ ((fiEnable && (8652 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3516_0 <=( _mesh_27_13_io_out_last_0) ^ ((fiEnable && (8653 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3517_0 <=( _mesh_28_13_io_out_last_0) ^ ((fiEnable && (8654 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3518_0 <=( _mesh_29_13_io_out_last_0) ^ ((fiEnable && (8655 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3519_0 <=( _mesh_30_13_io_out_last_0) ^ ((fiEnable && (8656 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3520_0 <=( io_in_last_14_0) ^ ((fiEnable && (8657 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3521_0 <=( _mesh_0_14_io_out_last_0) ^ ((fiEnable && (8658 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3522_0 <=( _mesh_1_14_io_out_last_0) ^ ((fiEnable && (8659 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3523_0 <=( _mesh_2_14_io_out_last_0) ^ ((fiEnable && (8660 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3524_0 <=( _mesh_3_14_io_out_last_0) ^ ((fiEnable && (8661 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3525_0 <=( _mesh_4_14_io_out_last_0) ^ ((fiEnable && (8662 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3526_0 <=( _mesh_5_14_io_out_last_0) ^ ((fiEnable && (8663 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3527_0 <=( _mesh_6_14_io_out_last_0) ^ ((fiEnable && (8664 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3528_0 <=( _mesh_7_14_io_out_last_0) ^ ((fiEnable && (8665 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3529_0 <=( _mesh_8_14_io_out_last_0) ^ ((fiEnable && (8666 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3530_0 <=( _mesh_9_14_io_out_last_0) ^ ((fiEnable && (8667 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3531_0 <=( _mesh_10_14_io_out_last_0) ^ ((fiEnable && (8668 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3532_0 <=( _mesh_11_14_io_out_last_0) ^ ((fiEnable && (8669 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3533_0 <=( _mesh_12_14_io_out_last_0) ^ ((fiEnable && (8670 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3534_0 <=( _mesh_13_14_io_out_last_0) ^ ((fiEnable && (8671 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3535_0 <=( _mesh_14_14_io_out_last_0) ^ ((fiEnable && (8672 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3536_0 <=( _mesh_15_14_io_out_last_0) ^ ((fiEnable && (8673 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3537_0 <=( _mesh_16_14_io_out_last_0) ^ ((fiEnable && (8674 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3538_0 <=( _mesh_17_14_io_out_last_0) ^ ((fiEnable && (8675 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3539_0 <=( _mesh_18_14_io_out_last_0) ^ ((fiEnable && (8676 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3540_0 <=( _mesh_19_14_io_out_last_0) ^ ((fiEnable && (8677 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3541_0 <=( _mesh_20_14_io_out_last_0) ^ ((fiEnable && (8678 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3542_0 <=( _mesh_21_14_io_out_last_0) ^ ((fiEnable && (8679 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3543_0 <=( _mesh_22_14_io_out_last_0) ^ ((fiEnable && (8680 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3544_0 <=( _mesh_23_14_io_out_last_0) ^ ((fiEnable && (8681 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3545_0 <=( _mesh_24_14_io_out_last_0) ^ ((fiEnable && (8682 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3546_0 <=( _mesh_25_14_io_out_last_0) ^ ((fiEnable && (8683 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3547_0 <=( _mesh_26_14_io_out_last_0) ^ ((fiEnable && (8684 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3548_0 <=( _mesh_27_14_io_out_last_0) ^ ((fiEnable && (8685 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3549_0 <=( _mesh_28_14_io_out_last_0) ^ ((fiEnable && (8686 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3550_0 <=( _mesh_29_14_io_out_last_0) ^ ((fiEnable && (8687 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3551_0 <=( _mesh_30_14_io_out_last_0) ^ ((fiEnable && (8688 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3552_0 <=( io_in_last_15_0) ^ ((fiEnable && (8689 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3553_0 <=( _mesh_0_15_io_out_last_0) ^ ((fiEnable && (8690 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3554_0 <=( _mesh_1_15_io_out_last_0) ^ ((fiEnable && (8691 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3555_0 <=( _mesh_2_15_io_out_last_0) ^ ((fiEnable && (8692 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3556_0 <=( _mesh_3_15_io_out_last_0) ^ ((fiEnable && (8693 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3557_0 <=( _mesh_4_15_io_out_last_0) ^ ((fiEnable && (8694 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3558_0 <=( _mesh_5_15_io_out_last_0) ^ ((fiEnable && (8695 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3559_0 <=( _mesh_6_15_io_out_last_0) ^ ((fiEnable && (8696 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3560_0 <=( _mesh_7_15_io_out_last_0) ^ ((fiEnable && (8697 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3561_0 <=( _mesh_8_15_io_out_last_0) ^ ((fiEnable && (8698 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3562_0 <=( _mesh_9_15_io_out_last_0) ^ ((fiEnable && (8699 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3563_0 <=( _mesh_10_15_io_out_last_0) ^ ((fiEnable && (8700 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3564_0 <=( _mesh_11_15_io_out_last_0) ^ ((fiEnable && (8701 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3565_0 <=( _mesh_12_15_io_out_last_0) ^ ((fiEnable && (8702 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3566_0 <=( _mesh_13_15_io_out_last_0) ^ ((fiEnable && (8703 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3567_0 <=( _mesh_14_15_io_out_last_0) ^ ((fiEnable && (8704 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3568_0 <=( _mesh_15_15_io_out_last_0) ^ ((fiEnable && (8705 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3569_0 <=( _mesh_16_15_io_out_last_0) ^ ((fiEnable && (8706 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3570_0 <=( _mesh_17_15_io_out_last_0) ^ ((fiEnable && (8707 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3571_0 <=( _mesh_18_15_io_out_last_0) ^ ((fiEnable && (8708 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3572_0 <=( _mesh_19_15_io_out_last_0) ^ ((fiEnable && (8709 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3573_0 <=( _mesh_20_15_io_out_last_0) ^ ((fiEnable && (8710 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3574_0 <=( _mesh_21_15_io_out_last_0) ^ ((fiEnable && (8711 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3575_0 <=( _mesh_22_15_io_out_last_0) ^ ((fiEnable && (8712 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3576_0 <=( _mesh_23_15_io_out_last_0) ^ ((fiEnable && (8713 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3577_0 <=( _mesh_24_15_io_out_last_0) ^ ((fiEnable && (8714 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3578_0 <=( _mesh_25_15_io_out_last_0) ^ ((fiEnable && (8715 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3579_0 <=( _mesh_26_15_io_out_last_0) ^ ((fiEnable && (8716 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3580_0 <=( _mesh_27_15_io_out_last_0) ^ ((fiEnable && (8717 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3581_0 <=( _mesh_28_15_io_out_last_0) ^ ((fiEnable && (8718 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3582_0 <=( _mesh_29_15_io_out_last_0) ^ ((fiEnable && (8719 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3583_0 <=( _mesh_30_15_io_out_last_0) ^ ((fiEnable && (8720 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3584_0 <=( io_in_last_16_0) ^ ((fiEnable && (8721 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3585_0 <=( _mesh_0_16_io_out_last_0) ^ ((fiEnable && (8722 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3586_0 <=( _mesh_1_16_io_out_last_0) ^ ((fiEnable && (8723 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3587_0 <=( _mesh_2_16_io_out_last_0) ^ ((fiEnable && (8724 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3588_0 <=( _mesh_3_16_io_out_last_0) ^ ((fiEnable && (8725 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3589_0 <=( _mesh_4_16_io_out_last_0) ^ ((fiEnable && (8726 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3590_0 <=( _mesh_5_16_io_out_last_0) ^ ((fiEnable && (8727 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3591_0 <=( _mesh_6_16_io_out_last_0) ^ ((fiEnable && (8728 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3592_0 <=( _mesh_7_16_io_out_last_0) ^ ((fiEnable && (8729 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3593_0 <=( _mesh_8_16_io_out_last_0) ^ ((fiEnable && (8730 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3594_0 <=( _mesh_9_16_io_out_last_0) ^ ((fiEnable && (8731 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3595_0 <=( _mesh_10_16_io_out_last_0) ^ ((fiEnable && (8732 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3596_0 <=( _mesh_11_16_io_out_last_0) ^ ((fiEnable && (8733 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3597_0 <=( _mesh_12_16_io_out_last_0) ^ ((fiEnable && (8734 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3598_0 <=( _mesh_13_16_io_out_last_0) ^ ((fiEnable && (8735 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3599_0 <=( _mesh_14_16_io_out_last_0) ^ ((fiEnable && (8736 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3600_0 <=( _mesh_15_16_io_out_last_0) ^ ((fiEnable && (8737 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3601_0 <=( _mesh_16_16_io_out_last_0) ^ ((fiEnable && (8738 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3602_0 <=( _mesh_17_16_io_out_last_0) ^ ((fiEnable && (8739 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3603_0 <=( _mesh_18_16_io_out_last_0) ^ ((fiEnable && (8740 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3604_0 <=( _mesh_19_16_io_out_last_0) ^ ((fiEnable && (8741 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3605_0 <=( _mesh_20_16_io_out_last_0) ^ ((fiEnable && (8742 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3606_0 <=( _mesh_21_16_io_out_last_0) ^ ((fiEnable && (8743 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3607_0 <=( _mesh_22_16_io_out_last_0) ^ ((fiEnable && (8744 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3608_0 <=( _mesh_23_16_io_out_last_0) ^ ((fiEnable && (8745 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3609_0 <=( _mesh_24_16_io_out_last_0) ^ ((fiEnable && (8746 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3610_0 <=( _mesh_25_16_io_out_last_0) ^ ((fiEnable && (8747 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3611_0 <=( _mesh_26_16_io_out_last_0) ^ ((fiEnable && (8748 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3612_0 <=( _mesh_27_16_io_out_last_0) ^ ((fiEnable && (8749 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3613_0 <=( _mesh_28_16_io_out_last_0) ^ ((fiEnable && (8750 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3614_0 <=( _mesh_29_16_io_out_last_0) ^ ((fiEnable && (8751 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3615_0 <=( _mesh_30_16_io_out_last_0) ^ ((fiEnable && (8752 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3616_0 <=( io_in_last_17_0) ^ ((fiEnable && (8753 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3617_0 <=( _mesh_0_17_io_out_last_0) ^ ((fiEnable && (8754 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3618_0 <=( _mesh_1_17_io_out_last_0) ^ ((fiEnable && (8755 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3619_0 <=( _mesh_2_17_io_out_last_0) ^ ((fiEnable && (8756 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3620_0 <=( _mesh_3_17_io_out_last_0) ^ ((fiEnable && (8757 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3621_0 <=( _mesh_4_17_io_out_last_0) ^ ((fiEnable && (8758 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3622_0 <=( _mesh_5_17_io_out_last_0) ^ ((fiEnable && (8759 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3623_0 <=( _mesh_6_17_io_out_last_0) ^ ((fiEnable && (8760 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3624_0 <=( _mesh_7_17_io_out_last_0) ^ ((fiEnable && (8761 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3625_0 <=( _mesh_8_17_io_out_last_0) ^ ((fiEnable && (8762 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3626_0 <=( _mesh_9_17_io_out_last_0) ^ ((fiEnable && (8763 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3627_0 <=( _mesh_10_17_io_out_last_0) ^ ((fiEnable && (8764 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3628_0 <=( _mesh_11_17_io_out_last_0) ^ ((fiEnable && (8765 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3629_0 <=( _mesh_12_17_io_out_last_0) ^ ((fiEnable && (8766 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3630_0 <=( _mesh_13_17_io_out_last_0) ^ ((fiEnable && (8767 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3631_0 <=( _mesh_14_17_io_out_last_0) ^ ((fiEnable && (8768 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3632_0 <=( _mesh_15_17_io_out_last_0) ^ ((fiEnable && (8769 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3633_0 <=( _mesh_16_17_io_out_last_0) ^ ((fiEnable && (8770 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3634_0 <=( _mesh_17_17_io_out_last_0) ^ ((fiEnable && (8771 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3635_0 <=( _mesh_18_17_io_out_last_0) ^ ((fiEnable && (8772 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3636_0 <=( _mesh_19_17_io_out_last_0) ^ ((fiEnable && (8773 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3637_0 <=( _mesh_20_17_io_out_last_0) ^ ((fiEnable && (8774 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3638_0 <=( _mesh_21_17_io_out_last_0) ^ ((fiEnable && (8775 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3639_0 <=( _mesh_22_17_io_out_last_0) ^ ((fiEnable && (8776 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3640_0 <=( _mesh_23_17_io_out_last_0) ^ ((fiEnable && (8777 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3641_0 <=( _mesh_24_17_io_out_last_0) ^ ((fiEnable && (8778 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3642_0 <=( _mesh_25_17_io_out_last_0) ^ ((fiEnable && (8779 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3643_0 <=( _mesh_26_17_io_out_last_0) ^ ((fiEnable && (8780 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3644_0 <=( _mesh_27_17_io_out_last_0) ^ ((fiEnable && (8781 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3645_0 <=( _mesh_28_17_io_out_last_0) ^ ((fiEnable && (8782 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3646_0 <=( _mesh_29_17_io_out_last_0) ^ ((fiEnable && (8783 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3647_0 <=( _mesh_30_17_io_out_last_0) ^ ((fiEnable && (8784 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3648_0 <=( io_in_last_18_0) ^ ((fiEnable && (8785 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3649_0 <=( _mesh_0_18_io_out_last_0) ^ ((fiEnable && (8786 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3650_0 <=( _mesh_1_18_io_out_last_0) ^ ((fiEnable && (8787 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3651_0 <=( _mesh_2_18_io_out_last_0) ^ ((fiEnable && (8788 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3652_0 <=( _mesh_3_18_io_out_last_0) ^ ((fiEnable && (8789 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3653_0 <=( _mesh_4_18_io_out_last_0) ^ ((fiEnable && (8790 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3654_0 <=( _mesh_5_18_io_out_last_0) ^ ((fiEnable && (8791 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3655_0 <=( _mesh_6_18_io_out_last_0) ^ ((fiEnable && (8792 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3656_0 <=( _mesh_7_18_io_out_last_0) ^ ((fiEnable && (8793 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3657_0 <=( _mesh_8_18_io_out_last_0) ^ ((fiEnable && (8794 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3658_0 <=( _mesh_9_18_io_out_last_0) ^ ((fiEnable && (8795 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3659_0 <=( _mesh_10_18_io_out_last_0) ^ ((fiEnable && (8796 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3660_0 <=( _mesh_11_18_io_out_last_0) ^ ((fiEnable && (8797 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3661_0 <=( _mesh_12_18_io_out_last_0) ^ ((fiEnable && (8798 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3662_0 <=( _mesh_13_18_io_out_last_0) ^ ((fiEnable && (8799 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3663_0 <=( _mesh_14_18_io_out_last_0) ^ ((fiEnable && (8800 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3664_0 <=( _mesh_15_18_io_out_last_0) ^ ((fiEnable && (8801 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3665_0 <=( _mesh_16_18_io_out_last_0) ^ ((fiEnable && (8802 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3666_0 <=( _mesh_17_18_io_out_last_0) ^ ((fiEnable && (8803 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3667_0 <=( _mesh_18_18_io_out_last_0) ^ ((fiEnable && (8804 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3668_0 <=( _mesh_19_18_io_out_last_0) ^ ((fiEnable && (8805 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3669_0 <=( _mesh_20_18_io_out_last_0) ^ ((fiEnable && (8806 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3670_0 <=( _mesh_21_18_io_out_last_0) ^ ((fiEnable && (8807 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3671_0 <=( _mesh_22_18_io_out_last_0) ^ ((fiEnable && (8808 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3672_0 <=( _mesh_23_18_io_out_last_0) ^ ((fiEnable && (8809 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3673_0 <=( _mesh_24_18_io_out_last_0) ^ ((fiEnable && (8810 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3674_0 <=( _mesh_25_18_io_out_last_0) ^ ((fiEnable && (8811 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3675_0 <=( _mesh_26_18_io_out_last_0) ^ ((fiEnable && (8812 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3676_0 <=( _mesh_27_18_io_out_last_0) ^ ((fiEnable && (8813 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3677_0 <=( _mesh_28_18_io_out_last_0) ^ ((fiEnable && (8814 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3678_0 <=( _mesh_29_18_io_out_last_0) ^ ((fiEnable && (8815 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3679_0 <=( _mesh_30_18_io_out_last_0) ^ ((fiEnable && (8816 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3680_0 <=( io_in_last_19_0) ^ ((fiEnable && (8817 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3681_0 <=( _mesh_0_19_io_out_last_0) ^ ((fiEnable && (8818 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3682_0 <=( _mesh_1_19_io_out_last_0) ^ ((fiEnable && (8819 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3683_0 <=( _mesh_2_19_io_out_last_0) ^ ((fiEnable && (8820 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3684_0 <=( _mesh_3_19_io_out_last_0) ^ ((fiEnable && (8821 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3685_0 <=( _mesh_4_19_io_out_last_0) ^ ((fiEnable && (8822 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3686_0 <=( _mesh_5_19_io_out_last_0) ^ ((fiEnable && (8823 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3687_0 <=( _mesh_6_19_io_out_last_0) ^ ((fiEnable && (8824 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3688_0 <=( _mesh_7_19_io_out_last_0) ^ ((fiEnable && (8825 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3689_0 <=( _mesh_8_19_io_out_last_0) ^ ((fiEnable && (8826 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3690_0 <=( _mesh_9_19_io_out_last_0) ^ ((fiEnable && (8827 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3691_0 <=( _mesh_10_19_io_out_last_0) ^ ((fiEnable && (8828 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3692_0 <=( _mesh_11_19_io_out_last_0) ^ ((fiEnable && (8829 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3693_0 <=( _mesh_12_19_io_out_last_0) ^ ((fiEnable && (8830 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3694_0 <=( _mesh_13_19_io_out_last_0) ^ ((fiEnable && (8831 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3695_0 <=( _mesh_14_19_io_out_last_0) ^ ((fiEnable && (8832 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3696_0 <=( _mesh_15_19_io_out_last_0) ^ ((fiEnable && (8833 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3697_0 <=( _mesh_16_19_io_out_last_0) ^ ((fiEnable && (8834 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3698_0 <=( _mesh_17_19_io_out_last_0) ^ ((fiEnable && (8835 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3699_0 <=( _mesh_18_19_io_out_last_0) ^ ((fiEnable && (8836 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3700_0 <=( _mesh_19_19_io_out_last_0) ^ ((fiEnable && (8837 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3701_0 <=( _mesh_20_19_io_out_last_0) ^ ((fiEnable && (8838 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3702_0 <=( _mesh_21_19_io_out_last_0) ^ ((fiEnable && (8839 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3703_0 <=( _mesh_22_19_io_out_last_0) ^ ((fiEnable && (8840 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3704_0 <=( _mesh_23_19_io_out_last_0) ^ ((fiEnable && (8841 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3705_0 <=( _mesh_24_19_io_out_last_0) ^ ((fiEnable && (8842 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3706_0 <=( _mesh_25_19_io_out_last_0) ^ ((fiEnable && (8843 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3707_0 <=( _mesh_26_19_io_out_last_0) ^ ((fiEnable && (8844 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3708_0 <=( _mesh_27_19_io_out_last_0) ^ ((fiEnable && (8845 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3709_0 <=( _mesh_28_19_io_out_last_0) ^ ((fiEnable && (8846 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3710_0 <=( _mesh_29_19_io_out_last_0) ^ ((fiEnable && (8847 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3711_0 <=( _mesh_30_19_io_out_last_0) ^ ((fiEnable && (8848 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3712_0 <=( io_in_last_20_0) ^ ((fiEnable && (8849 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3713_0 <=( _mesh_0_20_io_out_last_0) ^ ((fiEnable && (8850 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3714_0 <=( _mesh_1_20_io_out_last_0) ^ ((fiEnable && (8851 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3715_0 <=( _mesh_2_20_io_out_last_0) ^ ((fiEnable && (8852 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3716_0 <=( _mesh_3_20_io_out_last_0) ^ ((fiEnable && (8853 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3717_0 <=( _mesh_4_20_io_out_last_0) ^ ((fiEnable && (8854 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3718_0 <=( _mesh_5_20_io_out_last_0) ^ ((fiEnable && (8855 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3719_0 <=( _mesh_6_20_io_out_last_0) ^ ((fiEnable && (8856 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3720_0 <=( _mesh_7_20_io_out_last_0) ^ ((fiEnable && (8857 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3721_0 <=( _mesh_8_20_io_out_last_0) ^ ((fiEnable && (8858 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3722_0 <=( _mesh_9_20_io_out_last_0) ^ ((fiEnable && (8859 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3723_0 <=( _mesh_10_20_io_out_last_0) ^ ((fiEnable && (8860 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3724_0 <=( _mesh_11_20_io_out_last_0) ^ ((fiEnable && (8861 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3725_0 <=( _mesh_12_20_io_out_last_0) ^ ((fiEnable && (8862 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3726_0 <=( _mesh_13_20_io_out_last_0) ^ ((fiEnable && (8863 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3727_0 <=( _mesh_14_20_io_out_last_0) ^ ((fiEnable && (8864 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3728_0 <=( _mesh_15_20_io_out_last_0) ^ ((fiEnable && (8865 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3729_0 <=( _mesh_16_20_io_out_last_0) ^ ((fiEnable && (8866 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3730_0 <=( _mesh_17_20_io_out_last_0) ^ ((fiEnable && (8867 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3731_0 <=( _mesh_18_20_io_out_last_0) ^ ((fiEnable && (8868 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3732_0 <=( _mesh_19_20_io_out_last_0) ^ ((fiEnable && (8869 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3733_0 <=( _mesh_20_20_io_out_last_0) ^ ((fiEnable && (8870 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3734_0 <=( _mesh_21_20_io_out_last_0) ^ ((fiEnable && (8871 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3735_0 <=( _mesh_22_20_io_out_last_0) ^ ((fiEnable && (8872 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3736_0 <=( _mesh_23_20_io_out_last_0) ^ ((fiEnable && (8873 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3737_0 <=( _mesh_24_20_io_out_last_0) ^ ((fiEnable && (8874 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3738_0 <=( _mesh_25_20_io_out_last_0) ^ ((fiEnable && (8875 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3739_0 <=( _mesh_26_20_io_out_last_0) ^ ((fiEnable && (8876 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3740_0 <=( _mesh_27_20_io_out_last_0) ^ ((fiEnable && (8877 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3741_0 <=( _mesh_28_20_io_out_last_0) ^ ((fiEnable && (8878 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3742_0 <=( _mesh_29_20_io_out_last_0) ^ ((fiEnable && (8879 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3743_0 <=( _mesh_30_20_io_out_last_0) ^ ((fiEnable && (8880 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3744_0 <=( io_in_last_21_0) ^ ((fiEnable && (8881 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3745_0 <=( _mesh_0_21_io_out_last_0) ^ ((fiEnable && (8882 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3746_0 <=( _mesh_1_21_io_out_last_0) ^ ((fiEnable && (8883 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3747_0 <=( _mesh_2_21_io_out_last_0) ^ ((fiEnable && (8884 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3748_0 <=( _mesh_3_21_io_out_last_0) ^ ((fiEnable && (8885 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3749_0 <=( _mesh_4_21_io_out_last_0) ^ ((fiEnable && (8886 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3750_0 <=( _mesh_5_21_io_out_last_0) ^ ((fiEnable && (8887 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3751_0 <=( _mesh_6_21_io_out_last_0) ^ ((fiEnable && (8888 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3752_0 <=( _mesh_7_21_io_out_last_0) ^ ((fiEnable && (8889 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3753_0 <=( _mesh_8_21_io_out_last_0) ^ ((fiEnable && (8890 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3754_0 <=( _mesh_9_21_io_out_last_0) ^ ((fiEnable && (8891 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3755_0 <=( _mesh_10_21_io_out_last_0) ^ ((fiEnable && (8892 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3756_0 <=( _mesh_11_21_io_out_last_0) ^ ((fiEnable && (8893 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3757_0 <=( _mesh_12_21_io_out_last_0) ^ ((fiEnable && (8894 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3758_0 <=( _mesh_13_21_io_out_last_0) ^ ((fiEnable && (8895 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3759_0 <=( _mesh_14_21_io_out_last_0) ^ ((fiEnable && (8896 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3760_0 <=( _mesh_15_21_io_out_last_0) ^ ((fiEnable && (8897 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3761_0 <=( _mesh_16_21_io_out_last_0) ^ ((fiEnable && (8898 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3762_0 <=( _mesh_17_21_io_out_last_0) ^ ((fiEnable && (8899 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3763_0 <=( _mesh_18_21_io_out_last_0) ^ ((fiEnable && (8900 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3764_0 <=( _mesh_19_21_io_out_last_0) ^ ((fiEnable && (8901 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3765_0 <=( _mesh_20_21_io_out_last_0) ^ ((fiEnable && (8902 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3766_0 <=( _mesh_21_21_io_out_last_0) ^ ((fiEnable && (8903 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3767_0 <=( _mesh_22_21_io_out_last_0) ^ ((fiEnable && (8904 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3768_0 <=( _mesh_23_21_io_out_last_0) ^ ((fiEnable && (8905 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3769_0 <=( _mesh_24_21_io_out_last_0) ^ ((fiEnable && (8906 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3770_0 <=( _mesh_25_21_io_out_last_0) ^ ((fiEnable && (8907 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3771_0 <=( _mesh_26_21_io_out_last_0) ^ ((fiEnable && (8908 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3772_0 <=( _mesh_27_21_io_out_last_0) ^ ((fiEnable && (8909 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3773_0 <=( _mesh_28_21_io_out_last_0) ^ ((fiEnable && (8910 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3774_0 <=( _mesh_29_21_io_out_last_0) ^ ((fiEnable && (8911 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3775_0 <=( _mesh_30_21_io_out_last_0) ^ ((fiEnable && (8912 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3776_0 <=( io_in_last_22_0) ^ ((fiEnable && (8913 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3777_0 <=( _mesh_0_22_io_out_last_0) ^ ((fiEnable && (8914 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3778_0 <=( _mesh_1_22_io_out_last_0) ^ ((fiEnable && (8915 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3779_0 <=( _mesh_2_22_io_out_last_0) ^ ((fiEnable && (8916 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3780_0 <=( _mesh_3_22_io_out_last_0) ^ ((fiEnable && (8917 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3781_0 <=( _mesh_4_22_io_out_last_0) ^ ((fiEnable && (8918 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3782_0 <=( _mesh_5_22_io_out_last_0) ^ ((fiEnable && (8919 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3783_0 <=( _mesh_6_22_io_out_last_0) ^ ((fiEnable && (8920 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3784_0 <=( _mesh_7_22_io_out_last_0) ^ ((fiEnable && (8921 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3785_0 <=( _mesh_8_22_io_out_last_0) ^ ((fiEnable && (8922 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3786_0 <=( _mesh_9_22_io_out_last_0) ^ ((fiEnable && (8923 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3787_0 <=( _mesh_10_22_io_out_last_0) ^ ((fiEnable && (8924 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3788_0 <=( _mesh_11_22_io_out_last_0) ^ ((fiEnable && (8925 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3789_0 <=( _mesh_12_22_io_out_last_0) ^ ((fiEnable && (8926 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3790_0 <=( _mesh_13_22_io_out_last_0) ^ ((fiEnable && (8927 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3791_0 <=( _mesh_14_22_io_out_last_0) ^ ((fiEnable && (8928 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3792_0 <=( _mesh_15_22_io_out_last_0) ^ ((fiEnable && (8929 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3793_0 <=( _mesh_16_22_io_out_last_0) ^ ((fiEnable && (8930 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3794_0 <=( _mesh_17_22_io_out_last_0) ^ ((fiEnable && (8931 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3795_0 <=( _mesh_18_22_io_out_last_0) ^ ((fiEnable && (8932 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3796_0 <=( _mesh_19_22_io_out_last_0) ^ ((fiEnable && (8933 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3797_0 <=( _mesh_20_22_io_out_last_0) ^ ((fiEnable && (8934 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3798_0 <=( _mesh_21_22_io_out_last_0) ^ ((fiEnable && (8935 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3799_0 <=( _mesh_22_22_io_out_last_0) ^ ((fiEnable && (8936 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3800_0 <=( _mesh_23_22_io_out_last_0) ^ ((fiEnable && (8937 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3801_0 <=( _mesh_24_22_io_out_last_0) ^ ((fiEnable && (8938 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3802_0 <=( _mesh_25_22_io_out_last_0) ^ ((fiEnable && (8939 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3803_0 <=( _mesh_26_22_io_out_last_0) ^ ((fiEnable && (8940 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3804_0 <=( _mesh_27_22_io_out_last_0) ^ ((fiEnable && (8941 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3805_0 <=( _mesh_28_22_io_out_last_0) ^ ((fiEnable && (8942 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3806_0 <=( _mesh_29_22_io_out_last_0) ^ ((fiEnable && (8943 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3807_0 <=( _mesh_30_22_io_out_last_0) ^ ((fiEnable && (8944 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3808_0 <=( io_in_last_23_0) ^ ((fiEnable && (8945 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3809_0 <=( _mesh_0_23_io_out_last_0) ^ ((fiEnable && (8946 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3810_0 <=( _mesh_1_23_io_out_last_0) ^ ((fiEnable && (8947 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3811_0 <=( _mesh_2_23_io_out_last_0) ^ ((fiEnable && (8948 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3812_0 <=( _mesh_3_23_io_out_last_0) ^ ((fiEnable && (8949 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3813_0 <=( _mesh_4_23_io_out_last_0) ^ ((fiEnable && (8950 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3814_0 <=( _mesh_5_23_io_out_last_0) ^ ((fiEnable && (8951 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3815_0 <=( _mesh_6_23_io_out_last_0) ^ ((fiEnable && (8952 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3816_0 <=( _mesh_7_23_io_out_last_0) ^ ((fiEnable && (8953 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3817_0 <=( _mesh_8_23_io_out_last_0) ^ ((fiEnable && (8954 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3818_0 <=( _mesh_9_23_io_out_last_0) ^ ((fiEnable && (8955 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3819_0 <=( _mesh_10_23_io_out_last_0) ^ ((fiEnable && (8956 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3820_0 <=( _mesh_11_23_io_out_last_0) ^ ((fiEnable && (8957 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3821_0 <=( _mesh_12_23_io_out_last_0) ^ ((fiEnable && (8958 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3822_0 <=( _mesh_13_23_io_out_last_0) ^ ((fiEnable && (8959 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3823_0 <=( _mesh_14_23_io_out_last_0) ^ ((fiEnable && (8960 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3824_0 <=( _mesh_15_23_io_out_last_0) ^ ((fiEnable && (8961 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3825_0 <=( _mesh_16_23_io_out_last_0) ^ ((fiEnable && (8962 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3826_0 <=( _mesh_17_23_io_out_last_0) ^ ((fiEnable && (8963 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3827_0 <=( _mesh_18_23_io_out_last_0) ^ ((fiEnable && (8964 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3828_0 <=( _mesh_19_23_io_out_last_0) ^ ((fiEnable && (8965 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3829_0 <=( _mesh_20_23_io_out_last_0) ^ ((fiEnable && (8966 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3830_0 <=( _mesh_21_23_io_out_last_0) ^ ((fiEnable && (8967 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3831_0 <=( _mesh_22_23_io_out_last_0) ^ ((fiEnable && (8968 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3832_0 <=( _mesh_23_23_io_out_last_0) ^ ((fiEnable && (8969 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3833_0 <=( _mesh_24_23_io_out_last_0) ^ ((fiEnable && (8970 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3834_0 <=( _mesh_25_23_io_out_last_0) ^ ((fiEnable && (8971 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3835_0 <=( _mesh_26_23_io_out_last_0) ^ ((fiEnable && (8972 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3836_0 <=( _mesh_27_23_io_out_last_0) ^ ((fiEnable && (8973 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3837_0 <=( _mesh_28_23_io_out_last_0) ^ ((fiEnable && (8974 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3838_0 <=( _mesh_29_23_io_out_last_0) ^ ((fiEnable && (8975 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3839_0 <=( _mesh_30_23_io_out_last_0) ^ ((fiEnable && (8976 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3840_0 <=( io_in_last_24_0) ^ ((fiEnable && (8977 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3841_0 <=( _mesh_0_24_io_out_last_0) ^ ((fiEnable && (8978 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3842_0 <=( _mesh_1_24_io_out_last_0) ^ ((fiEnable && (8979 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3843_0 <=( _mesh_2_24_io_out_last_0) ^ ((fiEnable && (8980 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3844_0 <=( _mesh_3_24_io_out_last_0) ^ ((fiEnable && (8981 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3845_0 <=( _mesh_4_24_io_out_last_0) ^ ((fiEnable && (8982 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3846_0 <=( _mesh_5_24_io_out_last_0) ^ ((fiEnable && (8983 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3847_0 <=( _mesh_6_24_io_out_last_0) ^ ((fiEnable && (8984 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3848_0 <=( _mesh_7_24_io_out_last_0) ^ ((fiEnable && (8985 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3849_0 <=( _mesh_8_24_io_out_last_0) ^ ((fiEnable && (8986 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3850_0 <=( _mesh_9_24_io_out_last_0) ^ ((fiEnable && (8987 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3851_0 <=( _mesh_10_24_io_out_last_0) ^ ((fiEnable && (8988 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3852_0 <=( _mesh_11_24_io_out_last_0) ^ ((fiEnable && (8989 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3853_0 <=( _mesh_12_24_io_out_last_0) ^ ((fiEnable && (8990 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3854_0 <=( _mesh_13_24_io_out_last_0) ^ ((fiEnable && (8991 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3855_0 <=( _mesh_14_24_io_out_last_0) ^ ((fiEnable && (8992 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3856_0 <=( _mesh_15_24_io_out_last_0) ^ ((fiEnable && (8993 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3857_0 <=( _mesh_16_24_io_out_last_0) ^ ((fiEnable && (8994 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3858_0 <=( _mesh_17_24_io_out_last_0) ^ ((fiEnable && (8995 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3859_0 <=( _mesh_18_24_io_out_last_0) ^ ((fiEnable && (8996 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3860_0 <=( _mesh_19_24_io_out_last_0) ^ ((fiEnable && (8997 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3861_0 <=( _mesh_20_24_io_out_last_0) ^ ((fiEnable && (8998 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3862_0 <=( _mesh_21_24_io_out_last_0) ^ ((fiEnable && (8999 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3863_0 <=( _mesh_22_24_io_out_last_0) ^ ((fiEnable && (9000 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3864_0 <=( _mesh_23_24_io_out_last_0) ^ ((fiEnable && (9001 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3865_0 <=( _mesh_24_24_io_out_last_0) ^ ((fiEnable && (9002 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3866_0 <=( _mesh_25_24_io_out_last_0) ^ ((fiEnable && (9003 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3867_0 <=( _mesh_26_24_io_out_last_0) ^ ((fiEnable && (9004 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3868_0 <=( _mesh_27_24_io_out_last_0) ^ ((fiEnable && (9005 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3869_0 <=( _mesh_28_24_io_out_last_0) ^ ((fiEnable && (9006 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3870_0 <=( _mesh_29_24_io_out_last_0) ^ ((fiEnable && (9007 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3871_0 <=( _mesh_30_24_io_out_last_0) ^ ((fiEnable && (9008 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3872_0 <=( io_in_last_25_0) ^ ((fiEnable && (9009 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3873_0 <=( _mesh_0_25_io_out_last_0) ^ ((fiEnable && (9010 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3874_0 <=( _mesh_1_25_io_out_last_0) ^ ((fiEnable && (9011 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3875_0 <=( _mesh_2_25_io_out_last_0) ^ ((fiEnable && (9012 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3876_0 <=( _mesh_3_25_io_out_last_0) ^ ((fiEnable && (9013 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3877_0 <=( _mesh_4_25_io_out_last_0) ^ ((fiEnable && (9014 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3878_0 <=( _mesh_5_25_io_out_last_0) ^ ((fiEnable && (9015 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3879_0 <=( _mesh_6_25_io_out_last_0) ^ ((fiEnable && (9016 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3880_0 <=( _mesh_7_25_io_out_last_0) ^ ((fiEnable && (9017 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3881_0 <=( _mesh_8_25_io_out_last_0) ^ ((fiEnable && (9018 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3882_0 <=( _mesh_9_25_io_out_last_0) ^ ((fiEnable && (9019 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3883_0 <=( _mesh_10_25_io_out_last_0) ^ ((fiEnable && (9020 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3884_0 <=( _mesh_11_25_io_out_last_0) ^ ((fiEnable && (9021 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3885_0 <=( _mesh_12_25_io_out_last_0) ^ ((fiEnable && (9022 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3886_0 <=( _mesh_13_25_io_out_last_0) ^ ((fiEnable && (9023 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3887_0 <=( _mesh_14_25_io_out_last_0) ^ ((fiEnable && (9024 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3888_0 <=( _mesh_15_25_io_out_last_0) ^ ((fiEnable && (9025 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3889_0 <=( _mesh_16_25_io_out_last_0) ^ ((fiEnable && (9026 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3890_0 <=( _mesh_17_25_io_out_last_0) ^ ((fiEnable && (9027 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3891_0 <=( _mesh_18_25_io_out_last_0) ^ ((fiEnable && (9028 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3892_0 <=( _mesh_19_25_io_out_last_0) ^ ((fiEnable && (9029 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3893_0 <=( _mesh_20_25_io_out_last_0) ^ ((fiEnable && (9030 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3894_0 <=( _mesh_21_25_io_out_last_0) ^ ((fiEnable && (9031 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3895_0 <=( _mesh_22_25_io_out_last_0) ^ ((fiEnable && (9032 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3896_0 <=( _mesh_23_25_io_out_last_0) ^ ((fiEnable && (9033 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3897_0 <=( _mesh_24_25_io_out_last_0) ^ ((fiEnable && (9034 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3898_0 <=( _mesh_25_25_io_out_last_0) ^ ((fiEnable && (9035 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3899_0 <=( _mesh_26_25_io_out_last_0) ^ ((fiEnable && (9036 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3900_0 <=( _mesh_27_25_io_out_last_0) ^ ((fiEnable && (9037 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3901_0 <=( _mesh_28_25_io_out_last_0) ^ ((fiEnable && (9038 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3902_0 <=( _mesh_29_25_io_out_last_0) ^ ((fiEnable && (9039 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3903_0 <=( _mesh_30_25_io_out_last_0) ^ ((fiEnable && (9040 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3904_0 <=( io_in_last_26_0) ^ ((fiEnable && (9041 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3905_0 <=( _mesh_0_26_io_out_last_0) ^ ((fiEnable && (9042 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3906_0 <=( _mesh_1_26_io_out_last_0) ^ ((fiEnable && (9043 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3907_0 <=( _mesh_2_26_io_out_last_0) ^ ((fiEnable && (9044 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3908_0 <=( _mesh_3_26_io_out_last_0) ^ ((fiEnable && (9045 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3909_0 <=( _mesh_4_26_io_out_last_0) ^ ((fiEnable && (9046 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3910_0 <=( _mesh_5_26_io_out_last_0) ^ ((fiEnable && (9047 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3911_0 <=( _mesh_6_26_io_out_last_0) ^ ((fiEnable && (9048 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3912_0 <=( _mesh_7_26_io_out_last_0) ^ ((fiEnable && (9049 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3913_0 <=( _mesh_8_26_io_out_last_0) ^ ((fiEnable && (9050 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3914_0 <=( _mesh_9_26_io_out_last_0) ^ ((fiEnable && (9051 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3915_0 <=( _mesh_10_26_io_out_last_0) ^ ((fiEnable && (9052 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3916_0 <=( _mesh_11_26_io_out_last_0) ^ ((fiEnable && (9053 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3917_0 <=( _mesh_12_26_io_out_last_0) ^ ((fiEnable && (9054 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3918_0 <=( _mesh_13_26_io_out_last_0) ^ ((fiEnable && (9055 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3919_0 <=( _mesh_14_26_io_out_last_0) ^ ((fiEnable && (9056 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3920_0 <=( _mesh_15_26_io_out_last_0) ^ ((fiEnable && (9057 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3921_0 <=( _mesh_16_26_io_out_last_0) ^ ((fiEnable && (9058 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3922_0 <=( _mesh_17_26_io_out_last_0) ^ ((fiEnable && (9059 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3923_0 <=( _mesh_18_26_io_out_last_0) ^ ((fiEnable && (9060 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3924_0 <=( _mesh_19_26_io_out_last_0) ^ ((fiEnable && (9061 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3925_0 <=( _mesh_20_26_io_out_last_0) ^ ((fiEnable && (9062 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3926_0 <=( _mesh_21_26_io_out_last_0) ^ ((fiEnable && (9063 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3927_0 <=( _mesh_22_26_io_out_last_0) ^ ((fiEnable && (9064 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3928_0 <=( _mesh_23_26_io_out_last_0) ^ ((fiEnable && (9065 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3929_0 <=( _mesh_24_26_io_out_last_0) ^ ((fiEnable && (9066 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3930_0 <=( _mesh_25_26_io_out_last_0) ^ ((fiEnable && (9067 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3931_0 <=( _mesh_26_26_io_out_last_0) ^ ((fiEnable && (9068 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3932_0 <=( _mesh_27_26_io_out_last_0) ^ ((fiEnable && (9069 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3933_0 <=( _mesh_28_26_io_out_last_0) ^ ((fiEnable && (9070 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3934_0 <=( _mesh_29_26_io_out_last_0) ^ ((fiEnable && (9071 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3935_0 <=( _mesh_30_26_io_out_last_0) ^ ((fiEnable && (9072 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3936_0 <=( io_in_last_27_0) ^ ((fiEnable && (9073 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3937_0 <=( _mesh_0_27_io_out_last_0) ^ ((fiEnable && (9074 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3938_0 <=( _mesh_1_27_io_out_last_0) ^ ((fiEnable && (9075 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3939_0 <=( _mesh_2_27_io_out_last_0) ^ ((fiEnable && (9076 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3940_0 <=( _mesh_3_27_io_out_last_0) ^ ((fiEnable && (9077 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3941_0 <=( _mesh_4_27_io_out_last_0) ^ ((fiEnable && (9078 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3942_0 <=( _mesh_5_27_io_out_last_0) ^ ((fiEnable && (9079 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3943_0 <=( _mesh_6_27_io_out_last_0) ^ ((fiEnable && (9080 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3944_0 <=( _mesh_7_27_io_out_last_0) ^ ((fiEnable && (9081 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3945_0 <=( _mesh_8_27_io_out_last_0) ^ ((fiEnable && (9082 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3946_0 <=( _mesh_9_27_io_out_last_0) ^ ((fiEnable && (9083 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3947_0 <=( _mesh_10_27_io_out_last_0) ^ ((fiEnable && (9084 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3948_0 <=( _mesh_11_27_io_out_last_0) ^ ((fiEnable && (9085 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3949_0 <=( _mesh_12_27_io_out_last_0) ^ ((fiEnable && (9086 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3950_0 <=( _mesh_13_27_io_out_last_0) ^ ((fiEnable && (9087 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3951_0 <=( _mesh_14_27_io_out_last_0) ^ ((fiEnable && (9088 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3952_0 <=( _mesh_15_27_io_out_last_0) ^ ((fiEnable && (9089 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3953_0 <=( _mesh_16_27_io_out_last_0) ^ ((fiEnable && (9090 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3954_0 <=( _mesh_17_27_io_out_last_0) ^ ((fiEnable && (9091 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3955_0 <=( _mesh_18_27_io_out_last_0) ^ ((fiEnable && (9092 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3956_0 <=( _mesh_19_27_io_out_last_0) ^ ((fiEnable && (9093 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3957_0 <=( _mesh_20_27_io_out_last_0) ^ ((fiEnable && (9094 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3958_0 <=( _mesh_21_27_io_out_last_0) ^ ((fiEnable && (9095 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3959_0 <=( _mesh_22_27_io_out_last_0) ^ ((fiEnable && (9096 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3960_0 <=( _mesh_23_27_io_out_last_0) ^ ((fiEnable && (9097 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3961_0 <=( _mesh_24_27_io_out_last_0) ^ ((fiEnable && (9098 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3962_0 <=( _mesh_25_27_io_out_last_0) ^ ((fiEnable && (9099 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3963_0 <=( _mesh_26_27_io_out_last_0) ^ ((fiEnable && (9100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3964_0 <=( _mesh_27_27_io_out_last_0) ^ ((fiEnable && (9101 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3965_0 <=( _mesh_28_27_io_out_last_0) ^ ((fiEnable && (9102 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3966_0 <=( _mesh_29_27_io_out_last_0) ^ ((fiEnable && (9103 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3967_0 <=( _mesh_30_27_io_out_last_0) ^ ((fiEnable && (9104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3968_0 <=( io_in_last_28_0) ^ ((fiEnable && (9105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3969_0 <=( _mesh_0_28_io_out_last_0) ^ ((fiEnable && (9106 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3970_0 <=( _mesh_1_28_io_out_last_0) ^ ((fiEnable && (9107 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3971_0 <=( _mesh_2_28_io_out_last_0) ^ ((fiEnable && (9108 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3972_0 <=( _mesh_3_28_io_out_last_0) ^ ((fiEnable && (9109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3973_0 <=( _mesh_4_28_io_out_last_0) ^ ((fiEnable && (9110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3974_0 <=( _mesh_5_28_io_out_last_0) ^ ((fiEnable && (9111 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3975_0 <=( _mesh_6_28_io_out_last_0) ^ ((fiEnable && (9112 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3976_0 <=( _mesh_7_28_io_out_last_0) ^ ((fiEnable && (9113 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3977_0 <=( _mesh_8_28_io_out_last_0) ^ ((fiEnable && (9114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3978_0 <=( _mesh_9_28_io_out_last_0) ^ ((fiEnable && (9115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3979_0 <=( _mesh_10_28_io_out_last_0) ^ ((fiEnable && (9116 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3980_0 <=( _mesh_11_28_io_out_last_0) ^ ((fiEnable && (9117 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3981_0 <=( _mesh_12_28_io_out_last_0) ^ ((fiEnable && (9118 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3982_0 <=( _mesh_13_28_io_out_last_0) ^ ((fiEnable && (9119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3983_0 <=( _mesh_14_28_io_out_last_0) ^ ((fiEnable && (9120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3984_0 <=( _mesh_15_28_io_out_last_0) ^ ((fiEnable && (9121 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3985_0 <=( _mesh_16_28_io_out_last_0) ^ ((fiEnable && (9122 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3986_0 <=( _mesh_17_28_io_out_last_0) ^ ((fiEnable && (9123 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3987_0 <=( _mesh_18_28_io_out_last_0) ^ ((fiEnable && (9124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3988_0 <=( _mesh_19_28_io_out_last_0) ^ ((fiEnable && (9125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3989_0 <=( _mesh_20_28_io_out_last_0) ^ ((fiEnable && (9126 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3990_0 <=( _mesh_21_28_io_out_last_0) ^ ((fiEnable && (9127 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3991_0 <=( _mesh_22_28_io_out_last_0) ^ ((fiEnable && (9128 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3992_0 <=( _mesh_23_28_io_out_last_0) ^ ((fiEnable && (9129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3993_0 <=( _mesh_24_28_io_out_last_0) ^ ((fiEnable && (9130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3994_0 <=( _mesh_25_28_io_out_last_0) ^ ((fiEnable && (9131 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3995_0 <=( _mesh_26_28_io_out_last_0) ^ ((fiEnable && (9132 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3996_0 <=( _mesh_27_28_io_out_last_0) ^ ((fiEnable && (9133 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3997_0 <=( _mesh_28_28_io_out_last_0) ^ ((fiEnable && (9134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3998_0 <=( _mesh_29_28_io_out_last_0) ^ ((fiEnable && (9135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_3999_0 <=( _mesh_30_28_io_out_last_0) ^ ((fiEnable && (9136 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4000_0 <=( io_in_last_29_0) ^ ((fiEnable && (9137 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4001_0 <=( _mesh_0_29_io_out_last_0) ^ ((fiEnable && (9138 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4002_0 <=( _mesh_1_29_io_out_last_0) ^ ((fiEnable && (9139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4003_0 <=( _mesh_2_29_io_out_last_0) ^ ((fiEnable && (9140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4004_0 <=( _mesh_3_29_io_out_last_0) ^ ((fiEnable && (9141 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4005_0 <=( _mesh_4_29_io_out_last_0) ^ ((fiEnable && (9142 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4006_0 <=( _mesh_5_29_io_out_last_0) ^ ((fiEnable && (9143 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4007_0 <=( _mesh_6_29_io_out_last_0) ^ ((fiEnable && (9144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4008_0 <=( _mesh_7_29_io_out_last_0) ^ ((fiEnable && (9145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4009_0 <=( _mesh_8_29_io_out_last_0) ^ ((fiEnable && (9146 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4010_0 <=( _mesh_9_29_io_out_last_0) ^ ((fiEnable && (9147 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4011_0 <=( _mesh_10_29_io_out_last_0) ^ ((fiEnable && (9148 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4012_0 <=( _mesh_11_29_io_out_last_0) ^ ((fiEnable && (9149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4013_0 <=( _mesh_12_29_io_out_last_0) ^ ((fiEnable && (9150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4014_0 <=( _mesh_13_29_io_out_last_0) ^ ((fiEnable && (9151 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4015_0 <=( _mesh_14_29_io_out_last_0) ^ ((fiEnable && (9152 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4016_0 <=( _mesh_15_29_io_out_last_0) ^ ((fiEnable && (9153 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4017_0 <=( _mesh_16_29_io_out_last_0) ^ ((fiEnable && (9154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4018_0 <=( _mesh_17_29_io_out_last_0) ^ ((fiEnable && (9155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4019_0 <=( _mesh_18_29_io_out_last_0) ^ ((fiEnable && (9156 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4020_0 <=( _mesh_19_29_io_out_last_0) ^ ((fiEnable && (9157 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4021_0 <=( _mesh_20_29_io_out_last_0) ^ ((fiEnable && (9158 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4022_0 <=( _mesh_21_29_io_out_last_0) ^ ((fiEnable && (9159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4023_0 <=( _mesh_22_29_io_out_last_0) ^ ((fiEnable && (9160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4024_0 <=( _mesh_23_29_io_out_last_0) ^ ((fiEnable && (9161 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4025_0 <=( _mesh_24_29_io_out_last_0) ^ ((fiEnable && (9162 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4026_0 <=( _mesh_25_29_io_out_last_0) ^ ((fiEnable && (9163 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4027_0 <=( _mesh_26_29_io_out_last_0) ^ ((fiEnable && (9164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4028_0 <=( _mesh_27_29_io_out_last_0) ^ ((fiEnable && (9165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4029_0 <=( _mesh_28_29_io_out_last_0) ^ ((fiEnable && (9166 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4030_0 <=( _mesh_29_29_io_out_last_0) ^ ((fiEnable && (9167 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4031_0 <=( _mesh_30_29_io_out_last_0) ^ ((fiEnable && (9168 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4032_0 <=( io_in_last_30_0) ^ ((fiEnable && (9169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4033_0 <=( _mesh_0_30_io_out_last_0) ^ ((fiEnable && (9170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4034_0 <=( _mesh_1_30_io_out_last_0) ^ ((fiEnable && (9171 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4035_0 <=( _mesh_2_30_io_out_last_0) ^ ((fiEnable && (9172 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4036_0 <=( _mesh_3_30_io_out_last_0) ^ ((fiEnable && (9173 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4037_0 <=( _mesh_4_30_io_out_last_0) ^ ((fiEnable && (9174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4038_0 <=( _mesh_5_30_io_out_last_0) ^ ((fiEnable && (9175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4039_0 <=( _mesh_6_30_io_out_last_0) ^ ((fiEnable && (9176 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4040_0 <=( _mesh_7_30_io_out_last_0) ^ ((fiEnable && (9177 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4041_0 <=( _mesh_8_30_io_out_last_0) ^ ((fiEnable && (9178 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4042_0 <=( _mesh_9_30_io_out_last_0) ^ ((fiEnable && (9179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4043_0 <=( _mesh_10_30_io_out_last_0) ^ ((fiEnable && (9180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4044_0 <=( _mesh_11_30_io_out_last_0) ^ ((fiEnable && (9181 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4045_0 <=( _mesh_12_30_io_out_last_0) ^ ((fiEnable && (9182 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4046_0 <=( _mesh_13_30_io_out_last_0) ^ ((fiEnable && (9183 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4047_0 <=( _mesh_14_30_io_out_last_0) ^ ((fiEnable && (9184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4048_0 <=( _mesh_15_30_io_out_last_0) ^ ((fiEnable && (9185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4049_0 <=( _mesh_16_30_io_out_last_0) ^ ((fiEnable && (9186 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4050_0 <=( _mesh_17_30_io_out_last_0) ^ ((fiEnable && (9187 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4051_0 <=( _mesh_18_30_io_out_last_0) ^ ((fiEnable && (9188 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4052_0 <=( _mesh_19_30_io_out_last_0) ^ ((fiEnable && (9189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4053_0 <=( _mesh_20_30_io_out_last_0) ^ ((fiEnable && (9190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4054_0 <=( _mesh_21_30_io_out_last_0) ^ ((fiEnable && (9191 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4055_0 <=( _mesh_22_30_io_out_last_0) ^ ((fiEnable && (9192 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4056_0 <=( _mesh_23_30_io_out_last_0) ^ ((fiEnable && (9193 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4057_0 <=( _mesh_24_30_io_out_last_0) ^ ((fiEnable && (9194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4058_0 <=( _mesh_25_30_io_out_last_0) ^ ((fiEnable && (9195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4059_0 <=( _mesh_26_30_io_out_last_0) ^ ((fiEnable && (9196 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4060_0 <=( _mesh_27_30_io_out_last_0) ^ ((fiEnable && (9197 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4061_0 <=( _mesh_28_30_io_out_last_0) ^ ((fiEnable && (9198 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4062_0 <=( _mesh_29_30_io_out_last_0) ^ ((fiEnable && (9199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4063_0 <=( _mesh_30_30_io_out_last_0) ^ ((fiEnable && (9200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4064_0 <=( io_in_last_31_0) ^ ((fiEnable && (9201 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4065_0 <=( _mesh_0_31_io_out_last_0) ^ ((fiEnable && (9202 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4066_0 <=( _mesh_1_31_io_out_last_0) ^ ((fiEnable && (9203 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4067_0 <=( _mesh_2_31_io_out_last_0) ^ ((fiEnable && (9204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4068_0 <=( _mesh_3_31_io_out_last_0) ^ ((fiEnable && (9205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4069_0 <=( _mesh_4_31_io_out_last_0) ^ ((fiEnable && (9206 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4070_0 <=( _mesh_5_31_io_out_last_0) ^ ((fiEnable && (9207 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4071_0 <=( _mesh_6_31_io_out_last_0) ^ ((fiEnable && (9208 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4072_0 <=( _mesh_7_31_io_out_last_0) ^ ((fiEnable && (9209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4073_0 <=( _mesh_8_31_io_out_last_0) ^ ((fiEnable && (9210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4074_0 <=( _mesh_9_31_io_out_last_0) ^ ((fiEnable && (9211 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4075_0 <=( _mesh_10_31_io_out_last_0) ^ ((fiEnable && (9212 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4076_0 <=( _mesh_11_31_io_out_last_0) ^ ((fiEnable && (9213 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4077_0 <=( _mesh_12_31_io_out_last_0) ^ ((fiEnable && (9214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4078_0 <=( _mesh_13_31_io_out_last_0) ^ ((fiEnable && (9215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4079_0 <=( _mesh_14_31_io_out_last_0) ^ ((fiEnable && (9216 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4080_0 <=( _mesh_15_31_io_out_last_0) ^ ((fiEnable && (9217 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4081_0 <=( _mesh_16_31_io_out_last_0) ^ ((fiEnable && (9218 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4082_0 <=( _mesh_17_31_io_out_last_0) ^ ((fiEnable && (9219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4083_0 <=( _mesh_18_31_io_out_last_0) ^ ((fiEnable && (9220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4084_0 <=( _mesh_19_31_io_out_last_0) ^ ((fiEnable && (9221 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4085_0 <=( _mesh_20_31_io_out_last_0) ^ ((fiEnable && (9222 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4086_0 <=( _mesh_21_31_io_out_last_0) ^ ((fiEnable && (9223 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4087_0 <=( _mesh_22_31_io_out_last_0) ^ ((fiEnable && (9224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4088_0 <=( _mesh_23_31_io_out_last_0) ^ ((fiEnable && (9225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4089_0 <=( _mesh_24_31_io_out_last_0) ^ ((fiEnable && (9226 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4090_0 <=( _mesh_25_31_io_out_last_0) ^ ((fiEnable && (9227 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4091_0 <=( _mesh_26_31_io_out_last_0) ^ ((fiEnable && (9228 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4092_0 <=( _mesh_27_31_io_out_last_0) ^ ((fiEnable && (9229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4093_0 <=( _mesh_28_31_io_out_last_0) ^ ((fiEnable && (9230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4094_0 <=( _mesh_29_31_io_out_last_0) ^ ((fiEnable && (9231 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4095_0 <=( _mesh_30_31_io_out_last_0) ^ ((fiEnable && (9232 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4096_0 <=( _mesh_31_0_io_out_b_0) ^ ((fiEnable && (9233 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4097_0 <=( _mesh_31_0_io_out_c_0) ^ ((fiEnable && (9234 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4098_0 <=( _mesh_31_0_io_out_valid_0) ^ ((fiEnable && (9235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4099_0_dataflow <=( _mesh_31_0_io_out_control_0_dataflow) ^ ((fiEnable && (9236 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4100_0 <=( _mesh_31_0_io_out_id_0) ^ ((fiEnable && (9237 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_4101_0 <=( _mesh_31_0_io_out_last_0) ^ ((fiEnable && (9238 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_4102_0 <=( _mesh_31_1_io_out_b_0) ^ ((fiEnable && (9239 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4103_0 <=( _mesh_31_1_io_out_c_0) ^ ((fiEnable && (9240 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4108_0 <=( _mesh_31_2_io_out_b_0) ^ ((fiEnable && (9241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4109_0 <=( _mesh_31_2_io_out_c_0) ^ ((fiEnable && (9242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4114_0 <=( _mesh_31_3_io_out_b_0) ^ ((fiEnable && (9243 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4115_0 <=( _mesh_31_3_io_out_c_0) ^ ((fiEnable && (9244 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4120_0 <=( _mesh_31_4_io_out_b_0) ^ ((fiEnable && (9245 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4121_0 <=( _mesh_31_4_io_out_c_0) ^ ((fiEnable && (9246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4126_0 <=( _mesh_31_5_io_out_b_0) ^ ((fiEnable && (9247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4127_0 <=( _mesh_31_5_io_out_c_0) ^ ((fiEnable && (9248 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4132_0 <=( _mesh_31_6_io_out_b_0) ^ ((fiEnable && (9249 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4133_0 <=( _mesh_31_6_io_out_c_0) ^ ((fiEnable && (9250 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4138_0 <=( _mesh_31_7_io_out_b_0) ^ ((fiEnable && (9251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4139_0 <=( _mesh_31_7_io_out_c_0) ^ ((fiEnable && (9252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4144_0 <=( _mesh_31_8_io_out_b_0) ^ ((fiEnable && (9253 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4145_0 <=( _mesh_31_8_io_out_c_0) ^ ((fiEnable && (9254 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4150_0 <=( _mesh_31_9_io_out_b_0) ^ ((fiEnable && (9255 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4151_0 <=( _mesh_31_9_io_out_c_0) ^ ((fiEnable && (9256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4156_0 <=( _mesh_31_10_io_out_b_0) ^ ((fiEnable && (9257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4157_0 <=( _mesh_31_10_io_out_c_0) ^ ((fiEnable && (9258 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4162_0 <=( _mesh_31_11_io_out_b_0) ^ ((fiEnable && (9259 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4163_0 <=( _mesh_31_11_io_out_c_0) ^ ((fiEnable && (9260 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4168_0 <=( _mesh_31_12_io_out_b_0) ^ ((fiEnable && (9261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4169_0 <=( _mesh_31_12_io_out_c_0) ^ ((fiEnable && (9262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4174_0 <=( _mesh_31_13_io_out_b_0) ^ ((fiEnable && (9263 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4175_0 <=( _mesh_31_13_io_out_c_0) ^ ((fiEnable && (9264 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4180_0 <=( _mesh_31_14_io_out_b_0) ^ ((fiEnable && (9265 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4181_0 <=( _mesh_31_14_io_out_c_0) ^ ((fiEnable && (9266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4186_0 <=( _mesh_31_15_io_out_b_0) ^ ((fiEnable && (9267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4187_0 <=( _mesh_31_15_io_out_c_0) ^ ((fiEnable && (9268 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4192_0 <=( _mesh_31_16_io_out_b_0) ^ ((fiEnable && (9269 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4193_0 <=( _mesh_31_16_io_out_c_0) ^ ((fiEnable && (9270 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4198_0 <=( _mesh_31_17_io_out_b_0) ^ ((fiEnable && (9271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4199_0 <=( _mesh_31_17_io_out_c_0) ^ ((fiEnable && (9272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4204_0 <=( _mesh_31_18_io_out_b_0) ^ ((fiEnable && (9273 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4205_0 <=( _mesh_31_18_io_out_c_0) ^ ((fiEnable && (9274 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4210_0 <=( _mesh_31_19_io_out_b_0) ^ ((fiEnable && (9275 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4211_0 <=( _mesh_31_19_io_out_c_0) ^ ((fiEnable && (9276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4216_0 <=( _mesh_31_20_io_out_b_0) ^ ((fiEnable && (9277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4217_0 <=( _mesh_31_20_io_out_c_0) ^ ((fiEnable && (9278 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4222_0 <=( _mesh_31_21_io_out_b_0) ^ ((fiEnable && (9279 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4223_0 <=( _mesh_31_21_io_out_c_0) ^ ((fiEnable && (9280 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4228_0 <=( _mesh_31_22_io_out_b_0) ^ ((fiEnable && (9281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4229_0 <=( _mesh_31_22_io_out_c_0) ^ ((fiEnable && (9282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4234_0 <=( _mesh_31_23_io_out_b_0) ^ ((fiEnable && (9283 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4235_0 <=( _mesh_31_23_io_out_c_0) ^ ((fiEnable && (9284 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4240_0 <=( _mesh_31_24_io_out_b_0) ^ ((fiEnable && (9285 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4241_0 <=( _mesh_31_24_io_out_c_0) ^ ((fiEnable && (9286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4246_0 <=( _mesh_31_25_io_out_b_0) ^ ((fiEnable && (9287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4247_0 <=( _mesh_31_25_io_out_c_0) ^ ((fiEnable && (9288 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4252_0 <=( _mesh_31_26_io_out_b_0) ^ ((fiEnable && (9289 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4253_0 <=( _mesh_31_26_io_out_c_0) ^ ((fiEnable && (9290 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4258_0 <=( _mesh_31_27_io_out_b_0) ^ ((fiEnable && (9291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4259_0 <=( _mesh_31_27_io_out_c_0) ^ ((fiEnable && (9292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4264_0 <=( _mesh_31_28_io_out_b_0) ^ ((fiEnable && (9293 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4265_0 <=( _mesh_31_28_io_out_c_0) ^ ((fiEnable && (9294 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4270_0 <=( _mesh_31_29_io_out_b_0) ^ ((fiEnable && (9295 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4271_0 <=( _mesh_31_29_io_out_c_0) ^ ((fiEnable && (9296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4276_0 <=( _mesh_31_30_io_out_b_0) ^ ((fiEnable && (9297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4277_0 <=( _mesh_31_30_io_out_c_0) ^ ((fiEnable && (9298 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4282_0 <=( _mesh_31_31_io_out_b_0) ^ ((fiEnable && (9299 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4283_0 <=( _mesh_31_31_io_out_c_0) ^ ((fiEnable && (9300 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	logic [31:0] _RANDOM_3;
	logic [31:0] _RANDOM_4;
	logic [31:0] _RANDOM_5;
	logic [31:0] _RANDOM_6;
	logic [31:0] _RANDOM_7;
	logic [31:0] _RANDOM_8;
	logic [31:0] _RANDOM_9;
	logic [31:0] _RANDOM_10;
	logic [31:0] _RANDOM_11;
	logic [31:0] _RANDOM_12;
	logic [31:0] _RANDOM_13;
	logic [31:0] _RANDOM_14;
	logic [31:0] _RANDOM_15;
	logic [31:0] _RANDOM_16;
	logic [31:0] _RANDOM_17;
	logic [31:0] _RANDOM_18;
	logic [31:0] _RANDOM_19;
	logic [31:0] _RANDOM_20;
	logic [31:0] _RANDOM_21;
	logic [31:0] _RANDOM_22;
	logic [31:0] _RANDOM_23;
	logic [31:0] _RANDOM_24;
	logic [31:0] _RANDOM_25;
	logic [31:0] _RANDOM_26;
	logic [31:0] _RANDOM_27;
	logic [31:0] _RANDOM_28;
	logic [31:0] _RANDOM_29;
	logic [31:0] _RANDOM_30;
	logic [31:0] _RANDOM_31;
	logic [31:0] _RANDOM_32;
	logic [31:0] _RANDOM_33;
	logic [31:0] _RANDOM_34;
	logic [31:0] _RANDOM_35;
	logic [31:0] _RANDOM_36;
	logic [31:0] _RANDOM_37;
	logic [31:0] _RANDOM_38;
	logic [31:0] _RANDOM_39;
	logic [31:0] _RANDOM_40;
	logic [31:0] _RANDOM_41;
	logic [31:0] _RANDOM_42;
	logic [31:0] _RANDOM_43;
	logic [31:0] _RANDOM_44;
	logic [31:0] _RANDOM_45;
	logic [31:0] _RANDOM_46;
	logic [31:0] _RANDOM_47;
	logic [31:0] _RANDOM_48;
	logic [31:0] _RANDOM_49;
	logic [31:0] _RANDOM_50;
	logic [31:0] _RANDOM_51;
	logic [31:0] _RANDOM_52;
	logic [31:0] _RANDOM_53;
	logic [31:0] _RANDOM_54;
	logic [31:0] _RANDOM_55;
	logic [31:0] _RANDOM_56;
	logic [31:0] _RANDOM_57;
	logic [31:0] _RANDOM_58;
	logic [31:0] _RANDOM_59;
	logic [31:0] _RANDOM_60;
	logic [31:0] _RANDOM_61;
	logic [31:0] _RANDOM_62;
	logic [31:0] _RANDOM_63;
	logic [31:0] _RANDOM_64;
	logic [31:0] _RANDOM_65;
	logic [31:0] _RANDOM_66;
	logic [31:0] _RANDOM_67;
	logic [31:0] _RANDOM_68;
	logic [31:0] _RANDOM_69;
	logic [31:0] _RANDOM_70;
	logic [31:0] _RANDOM_71;
	logic [31:0] _RANDOM_72;
	logic [31:0] _RANDOM_73;
	logic [31:0] _RANDOM_74;
	logic [31:0] _RANDOM_75;
	logic [31:0] _RANDOM_76;
	logic [31:0] _RANDOM_77;
	logic [31:0] _RANDOM_78;
	logic [31:0] _RANDOM_79;
	logic [31:0] _RANDOM_80;
	logic [31:0] _RANDOM_81;
	logic [31:0] _RANDOM_82;
	logic [31:0] _RANDOM_83;
	logic [31:0] _RANDOM_84;
	logic [31:0] _RANDOM_85;
	logic [31:0] _RANDOM_86;
	logic [31:0] _RANDOM_87;
	logic [31:0] _RANDOM_88;
	logic [31:0] _RANDOM_89;
	logic [31:0] _RANDOM_90;
	logic [31:0] _RANDOM_91;
	logic [31:0] _RANDOM_92;
	logic [31:0] _RANDOM_93;
	logic [31:0] _RANDOM_94;
	logic [31:0] _RANDOM_95;
	logic [31:0] _RANDOM_96;
	logic [31:0] _RANDOM_97;
	logic [31:0] _RANDOM_98;
	logic [31:0] _RANDOM_99;
	logic [31:0] _RANDOM_100;
	logic [31:0] _RANDOM_101;
	logic [31:0] _RANDOM_102;
	logic [31:0] _RANDOM_103;
	logic [31:0] _RANDOM_104;
	logic [31:0] _RANDOM_105;
	logic [31:0] _RANDOM_106;
	logic [31:0] _RANDOM_107;
	logic [31:0] _RANDOM_108;
	logic [31:0] _RANDOM_109;
	logic [31:0] _RANDOM_110;
	logic [31:0] _RANDOM_111;
	logic [31:0] _RANDOM_112;
	logic [31:0] _RANDOM_113;
	logic [31:0] _RANDOM_114;
	logic [31:0] _RANDOM_115;
	logic [31:0] _RANDOM_116;
	logic [31:0] _RANDOM_117;
	logic [31:0] _RANDOM_118;
	logic [31:0] _RANDOM_119;
	logic [31:0] _RANDOM_120;
	logic [31:0] _RANDOM_121;
	logic [31:0] _RANDOM_122;
	logic [31:0] _RANDOM_123;
	logic [31:0] _RANDOM_124;
	logic [31:0] _RANDOM_125;
	logic [31:0] _RANDOM_126;
	logic [31:0] _RANDOM_127;
	logic [31:0] _RANDOM_128;
	logic [31:0] _RANDOM_129;
	logic [31:0] _RANDOM_130;
	logic [31:0] _RANDOM_131;
	logic [31:0] _RANDOM_132;
	logic [31:0] _RANDOM_133;
	logic [31:0] _RANDOM_134;
	logic [31:0] _RANDOM_135;
	logic [31:0] _RANDOM_136;
	logic [31:0] _RANDOM_137;
	logic [31:0] _RANDOM_138;
	logic [31:0] _RANDOM_139;
	logic [31:0] _RANDOM_140;
	logic [31:0] _RANDOM_141;
	logic [31:0] _RANDOM_142;
	logic [31:0] _RANDOM_143;
	logic [31:0] _RANDOM_144;
	logic [31:0] _RANDOM_145;
	logic [31:0] _RANDOM_146;
	logic [31:0] _RANDOM_147;
	logic [31:0] _RANDOM_148;
	logic [31:0] _RANDOM_149;
	logic [31:0] _RANDOM_150;
	logic [31:0] _RANDOM_151;
	logic [31:0] _RANDOM_152;
	logic [31:0] _RANDOM_153;
	logic [31:0] _RANDOM_154;
	logic [31:0] _RANDOM_155;
	logic [31:0] _RANDOM_156;
	logic [31:0] _RANDOM_157;
	logic [31:0] _RANDOM_158;
	logic [31:0] _RANDOM_159;
	logic [31:0] _RANDOM_160;
	logic [31:0] _RANDOM_161;
	logic [31:0] _RANDOM_162;
	logic [31:0] _RANDOM_163;
	logic [31:0] _RANDOM_164;
	logic [31:0] _RANDOM_165;
	logic [31:0] _RANDOM_166;
	logic [31:0] _RANDOM_167;
	logic [31:0] _RANDOM_168;
	logic [31:0] _RANDOM_169;
	logic [31:0] _RANDOM_170;
	logic [31:0] _RANDOM_171;
	logic [31:0] _RANDOM_172;
	logic [31:0] _RANDOM_173;
	logic [31:0] _RANDOM_174;
	logic [31:0] _RANDOM_175;
	logic [31:0] _RANDOM_176;
	logic [31:0] _RANDOM_177;
	logic [31:0] _RANDOM_178;
	logic [31:0] _RANDOM_179;
	logic [31:0] _RANDOM_180;
	logic [31:0] _RANDOM_181;
	logic [31:0] _RANDOM_182;
	logic [31:0] _RANDOM_183;
	logic [31:0] _RANDOM_184;
	logic [31:0] _RANDOM_185;
	logic [31:0] _RANDOM_186;
	logic [31:0] _RANDOM_187;
	logic [31:0] _RANDOM_188;
	logic [31:0] _RANDOM_189;
	logic [31:0] _RANDOM_190;
	logic [31:0] _RANDOM_191;
	logic [31:0] _RANDOM_192;
	logic [31:0] _RANDOM_193;
	logic [31:0] _RANDOM_194;
	logic [31:0] _RANDOM_195;
	logic [31:0] _RANDOM_196;
	logic [31:0] _RANDOM_197;
	logic [31:0] _RANDOM_198;
	logic [31:0] _RANDOM_199;
	logic [31:0] _RANDOM_200;
	logic [31:0] _RANDOM_201;
	logic [31:0] _RANDOM_202;
	logic [31:0] _RANDOM_203;
	logic [31:0] _RANDOM_204;
	logic [31:0] _RANDOM_205;
	logic [31:0] _RANDOM_206;
	logic [31:0] _RANDOM_207;
	logic [31:0] _RANDOM_208;
	logic [31:0] _RANDOM_209;
	logic [31:0] _RANDOM_210;
	logic [31:0] _RANDOM_211;
	logic [31:0] _RANDOM_212;
	logic [31:0] _RANDOM_213;
	logic [31:0] _RANDOM_214;
	logic [31:0] _RANDOM_215;
	logic [31:0] _RANDOM_216;
	logic [31:0] _RANDOM_217;
	logic [31:0] _RANDOM_218;
	logic [31:0] _RANDOM_219;
	logic [31:0] _RANDOM_220;
	logic [31:0] _RANDOM_221;
	logic [31:0] _RANDOM_222;
	logic [31:0] _RANDOM_223;
	logic [31:0] _RANDOM_224;
	logic [31:0] _RANDOM_225;
	logic [31:0] _RANDOM_226;
	logic [31:0] _RANDOM_227;
	logic [31:0] _RANDOM_228;
	logic [31:0] _RANDOM_229;
	logic [31:0] _RANDOM_230;
	logic [31:0] _RANDOM_231;
	logic [31:0] _RANDOM_232;
	logic [31:0] _RANDOM_233;
	logic [31:0] _RANDOM_234;
	logic [31:0] _RANDOM_235;
	logic [31:0] _RANDOM_236;
	logic [31:0] _RANDOM_237;
	logic [31:0] _RANDOM_238;
	logic [31:0] _RANDOM_239;
	logic [31:0] _RANDOM_240;
	logic [31:0] _RANDOM_241;
	logic [31:0] _RANDOM_242;
	logic [31:0] _RANDOM_243;
	logic [31:0] _RANDOM_244;
	logic [31:0] _RANDOM_245;
	logic [31:0] _RANDOM_246;
	logic [31:0] _RANDOM_247;
	logic [31:0] _RANDOM_248;
	logic [31:0] _RANDOM_249;
	logic [31:0] _RANDOM_250;
	logic [31:0] _RANDOM_251;
	logic [31:0] _RANDOM_252;
	logic [31:0] _RANDOM_253;
	logic [31:0] _RANDOM_254;
	logic [31:0] _RANDOM_255;
	logic [31:0] _RANDOM_256;
	logic [31:0] _RANDOM_257;
	logic [31:0] _RANDOM_258;
	logic [31:0] _RANDOM_259;
	logic [31:0] _RANDOM_260;
	logic [31:0] _RANDOM_261;
	logic [31:0] _RANDOM_262;
	logic [31:0] _RANDOM_263;
	logic [31:0] _RANDOM_264;
	logic [31:0] _RANDOM_265;
	logic [31:0] _RANDOM_266;
	logic [31:0] _RANDOM_267;
	logic [31:0] _RANDOM_268;
	logic [31:0] _RANDOM_269;
	logic [31:0] _RANDOM_270;
	logic [31:0] _RANDOM_271;
	logic [31:0] _RANDOM_272;
	logic [31:0] _RANDOM_273;
	logic [31:0] _RANDOM_274;
	logic [31:0] _RANDOM_275;
	logic [31:0] _RANDOM_276;
	logic [31:0] _RANDOM_277;
	logic [31:0] _RANDOM_278;
	logic [31:0] _RANDOM_279;
	logic [31:0] _RANDOM_280;
	logic [31:0] _RANDOM_281;
	logic [31:0] _RANDOM_282;
	logic [31:0] _RANDOM_283;
	logic [31:0] _RANDOM_284;
	logic [31:0] _RANDOM_285;
	logic [31:0] _RANDOM_286;
	logic [31:0] _RANDOM_287;
	logic [31:0] _RANDOM_288;
	logic [31:0] _RANDOM_289;
	logic [31:0] _RANDOM_290;
	logic [31:0] _RANDOM_291;
	logic [31:0] _RANDOM_292;
	logic [31:0] _RANDOM_293;
	logic [31:0] _RANDOM_294;
	logic [31:0] _RANDOM_295;
	logic [31:0] _RANDOM_296;
	logic [31:0] _RANDOM_297;
	logic [31:0] _RANDOM_298;
	logic [31:0] _RANDOM_299;
	logic [31:0] _RANDOM_300;
	logic [31:0] _RANDOM_301;
	logic [31:0] _RANDOM_302;
	logic [31:0] _RANDOM_303;
	logic [31:0] _RANDOM_304;
	logic [31:0] _RANDOM_305;
	logic [31:0] _RANDOM_306;
	logic [31:0] _RANDOM_307;
	logic [31:0] _RANDOM_308;
	logic [31:0] _RANDOM_309;
	logic [31:0] _RANDOM_310;
	logic [31:0] _RANDOM_311;
	logic [31:0] _RANDOM_312;
	logic [31:0] _RANDOM_313;
	logic [31:0] _RANDOM_314;
	logic [31:0] _RANDOM_315;
	logic [31:0] _RANDOM_316;
	logic [31:0] _RANDOM_317;
	logic [31:0] _RANDOM_318;
	logic [31:0] _RANDOM_319;
	logic [31:0] _RANDOM_320;
	logic [31:0] _RANDOM_321;
	logic [31:0] _RANDOM_322;
	logic [31:0] _RANDOM_323;
	logic [31:0] _RANDOM_324;
	logic [31:0] _RANDOM_325;
	logic [31:0] _RANDOM_326;
	logic [31:0] _RANDOM_327;
	logic [31:0] _RANDOM_328;
	logic [31:0] _RANDOM_329;
	logic [31:0] _RANDOM_330;
	logic [31:0] _RANDOM_331;
	logic [31:0] _RANDOM_332;
	logic [31:0] _RANDOM_333;
	logic [31:0] _RANDOM_334;
	logic [31:0] _RANDOM_335;
	logic [31:0] _RANDOM_336;
	logic [31:0] _RANDOM_337;
	logic [31:0] _RANDOM_338;
	logic [31:0] _RANDOM_339;
	logic [31:0] _RANDOM_340;
	logic [31:0] _RANDOM_341;
	logic [31:0] _RANDOM_342;
	logic [31:0] _RANDOM_343;
	logic [31:0] _RANDOM_344;
	logic [31:0] _RANDOM_345;
	logic [31:0] _RANDOM_346;
	logic [31:0] _RANDOM_347;
	logic [31:0] _RANDOM_348;
	logic [31:0] _RANDOM_349;
	logic [31:0] _RANDOM_350;
	logic [31:0] _RANDOM_351;
	logic [31:0] _RANDOM_352;
	logic [31:0] _RANDOM_353;
	logic [31:0] _RANDOM_354;
	logic [31:0] _RANDOM_355;
	logic [31:0] _RANDOM_356;
	logic [31:0] _RANDOM_357;
	logic [31:0] _RANDOM_358;
	logic [31:0] _RANDOM_359;
	logic [31:0] _RANDOM_360;
	logic [31:0] _RANDOM_361;
	logic [31:0] _RANDOM_362;
	logic [31:0] _RANDOM_363;
	logic [31:0] _RANDOM_364;
	logic [31:0] _RANDOM_365;
	logic [31:0] _RANDOM_366;
	logic [31:0] _RANDOM_367;
	logic [31:0] _RANDOM_368;
	logic [31:0] _RANDOM_369;
	logic [31:0] _RANDOM_370;
	logic [31:0] _RANDOM_371;
	logic [31:0] _RANDOM_372;
	logic [31:0] _RANDOM_373;
	logic [31:0] _RANDOM_374;
	logic [31:0] _RANDOM_375;
	logic [31:0] _RANDOM_376;
	logic [31:0] _RANDOM_377;
	logic [31:0] _RANDOM_378;
	logic [31:0] _RANDOM_379;
	logic [31:0] _RANDOM_380;
	logic [31:0] _RANDOM_381;
	logic [31:0] _RANDOM_382;
	logic [31:0] _RANDOM_383;
	logic [31:0] _RANDOM_384;
	logic [31:0] _RANDOM_385;
	logic [31:0] _RANDOM_386;
	logic [31:0] _RANDOM_387;
	logic [31:0] _RANDOM_388;
	logic [31:0] _RANDOM_389;
	logic [31:0] _RANDOM_390;
	logic [31:0] _RANDOM_391;
	logic [31:0] _RANDOM_392;
	logic [31:0] _RANDOM_393;
	logic [31:0] _RANDOM_394;
	logic [31:0] _RANDOM_395;
	logic [31:0] _RANDOM_396;
	logic [31:0] _RANDOM_397;
	logic [31:0] _RANDOM_398;
	logic [31:0] _RANDOM_399;
	logic [31:0] _RANDOM_400;
	logic [31:0] _RANDOM_401;
	logic [31:0] _RANDOM_402;
	logic [31:0] _RANDOM_403;
	logic [31:0] _RANDOM_404;
	logic [31:0] _RANDOM_405;
	logic [31:0] _RANDOM_406;
	logic [31:0] _RANDOM_407;
	logic [31:0] _RANDOM_408;
	logic [31:0] _RANDOM_409;
	logic [31:0] _RANDOM_410;
	logic [31:0] _RANDOM_411;
	logic [31:0] _RANDOM_412;
	logic [31:0] _RANDOM_413;
	logic [31:0] _RANDOM_414;
	logic [31:0] _RANDOM_415;
	logic [31:0] _RANDOM_416;
	logic [31:0] _RANDOM_417;
	logic [31:0] _RANDOM_418;
	logic [31:0] _RANDOM_419;
	logic [31:0] _RANDOM_420;
	logic [31:0] _RANDOM_421;
	logic [31:0] _RANDOM_422;
	logic [31:0] _RANDOM_423;
	logic [31:0] _RANDOM_424;
	logic [31:0] _RANDOM_425;
	logic [31:0] _RANDOM_426;
	logic [31:0] _RANDOM_427;
	logic [31:0] _RANDOM_428;
	logic [31:0] _RANDOM_429;
	logic [31:0] _RANDOM_430;
	logic [31:0] _RANDOM_431;
	logic [31:0] _RANDOM_432;
	logic [31:0] _RANDOM_433;
	logic [31:0] _RANDOM_434;
	logic [31:0] _RANDOM_435;
	logic [31:0] _RANDOM_436;
	logic [31:0] _RANDOM_437;
	logic [31:0] _RANDOM_438;
	logic [31:0] _RANDOM_439;
	logic [31:0] _RANDOM_440;
	logic [31:0] _RANDOM_441;
	logic [31:0] _RANDOM_442;
	logic [31:0] _RANDOM_443;
	logic [31:0] _RANDOM_444;
	logic [31:0] _RANDOM_445;
	logic [31:0] _RANDOM_446;
	logic [31:0] _RANDOM_447;
	logic [31:0] _RANDOM_448;
	logic [31:0] _RANDOM_449;
	logic [31:0] _RANDOM_450;
	logic [31:0] _RANDOM_451;
	logic [31:0] _RANDOM_452;
	logic [31:0] _RANDOM_453;
	logic [31:0] _RANDOM_454;
	logic [31:0] _RANDOM_455;
	logic [31:0] _RANDOM_456;
	logic [31:0] _RANDOM_457;
	logic [31:0] _RANDOM_458;
	logic [31:0] _RANDOM_459;
	logic [31:0] _RANDOM_460;
	logic [31:0] _RANDOM_461;
	logic [31:0] _RANDOM_462;
	logic [31:0] _RANDOM_463;
	logic [31:0] _RANDOM_464;
	logic [31:0] _RANDOM_465;
	logic [31:0] _RANDOM_466;
	logic [31:0] _RANDOM_467;
	logic [31:0] _RANDOM_468;
	logic [31:0] _RANDOM_469;
	logic [31:0] _RANDOM_470;
	logic [31:0] _RANDOM_471;
	logic [31:0] _RANDOM_472;
	logic [31:0] _RANDOM_473;
	logic [31:0] _RANDOM_474;
	logic [31:0] _RANDOM_475;
	logic [31:0] _RANDOM_476;
	logic [31:0] _RANDOM_477;
	logic [31:0] _RANDOM_478;
	logic [31:0] _RANDOM_479;
	logic [31:0] _RANDOM_480;
	logic [31:0] _RANDOM_481;
	logic [31:0] _RANDOM_482;
	logic [31:0] _RANDOM_483;
	logic [31:0] _RANDOM_484;
	logic [31:0] _RANDOM_485;
	logic [31:0] _RANDOM_486;
	logic [31:0] _RANDOM_487;
	logic [31:0] _RANDOM_488;
	logic [31:0] _RANDOM_489;
	logic [31:0] _RANDOM_490;
	logic [31:0] _RANDOM_491;
	logic [31:0] _RANDOM_492;
	logic [31:0] _RANDOM_493;
	logic [31:0] _RANDOM_494;
	logic [31:0] _RANDOM_495;
	logic [31:0] _RANDOM_496;
	logic [31:0] _RANDOM_497;
	logic [31:0] _RANDOM_498;
	logic [31:0] _RANDOM_499;
	logic [31:0] _RANDOM_500;
	logic [31:0] _RANDOM_501;
	logic [31:0] _RANDOM_502;
	logic [31:0] _RANDOM_503;
	logic [31:0] _RANDOM_504;
	logic [31:0] _RANDOM_505;
	logic [31:0] _RANDOM_506;
	logic [31:0] _RANDOM_507;
	logic [31:0] _RANDOM_508;
	logic [31:0] _RANDOM_509;
	logic [31:0] _RANDOM_510;
	logic [31:0] _RANDOM_511;
	logic [31:0] _RANDOM_512;
	logic [31:0] _RANDOM_513;
	logic [31:0] _RANDOM_514;
	logic [31:0] _RANDOM_515;
	logic [31:0] _RANDOM_516;
	logic [31:0] _RANDOM_517;
	logic [31:0] _RANDOM_518;
	logic [31:0] _RANDOM_519;
	logic [31:0] _RANDOM_520;
	logic [31:0] _RANDOM_521;
	logic [31:0] _RANDOM_522;
	logic [31:0] _RANDOM_523;
	logic [31:0] _RANDOM_524;
	logic [31:0] _RANDOM_525;
	logic [31:0] _RANDOM_526;
	logic [31:0] _RANDOM_527;
	logic [31:0] _RANDOM_528;
	logic [31:0] _RANDOM_529;
	logic [31:0] _RANDOM_530;
	logic [31:0] _RANDOM_531;
	logic [31:0] _RANDOM_532;
	logic [31:0] _RANDOM_533;
	logic [31:0] _RANDOM_534;
	logic [31:0] _RANDOM_535;
	logic [31:0] _RANDOM_536;
	logic [31:0] _RANDOM_537;
	logic [31:0] _RANDOM_538;
	logic [31:0] _RANDOM_539;
	logic [31:0] _RANDOM_540;
	logic [31:0] _RANDOM_541;
	logic [31:0] _RANDOM_542;
	logic [31:0] _RANDOM_543;
	logic [31:0] _RANDOM_544;
	logic [31:0] _RANDOM_545;
	logic [31:0] _RANDOM_546;
	logic [31:0] _RANDOM_547;
	logic [31:0] _RANDOM_548;
	logic [31:0] _RANDOM_549;
	logic [31:0] _RANDOM_550;
	logic [31:0] _RANDOM_551;
	logic [31:0] _RANDOM_552;
	logic [31:0] _RANDOM_553;
	logic [31:0] _RANDOM_554;
	logic [31:0] _RANDOM_555;
	logic [31:0] _RANDOM_556;
	logic [31:0] _RANDOM_557;
	logic [31:0] _RANDOM_558;
	logic [31:0] _RANDOM_559;
	logic [31:0] _RANDOM_560;
	logic [31:0] _RANDOM_561;
	logic [31:0] _RANDOM_562;
	logic [31:0] _RANDOM_563;
	logic [31:0] _RANDOM_564;
	logic [31:0] _RANDOM_565;
	logic [31:0] _RANDOM_566;
	logic [31:0] _RANDOM_567;
	logic [31:0] _RANDOM_568;
	logic [31:0] _RANDOM_569;
	logic [31:0] _RANDOM_570;
	logic [31:0] _RANDOM_571;
	logic [31:0] _RANDOM_572;
	logic [31:0] _RANDOM_573;
	logic [31:0] _RANDOM_574;
	logic [31:0] _RANDOM_575;
	logic [31:0] _RANDOM_576;
	logic [31:0] _RANDOM_577;
	logic [31:0] _RANDOM_578;
	logic [31:0] _RANDOM_579;
	logic [31:0] _RANDOM_580;
	logic [31:0] _RANDOM_581;
	logic [31:0] _RANDOM_582;
	logic [31:0] _RANDOM_583;
	logic [31:0] _RANDOM_584;
	logic [31:0] _RANDOM_585;
	logic [31:0] _RANDOM_586;
	logic [31:0] _RANDOM_587;
	logic [31:0] _RANDOM_588;
	logic [31:0] _RANDOM_589;
	logic [31:0] _RANDOM_590;
	logic [31:0] _RANDOM_591;
	logic [31:0] _RANDOM_592;
	logic [31:0] _RANDOM_593;
	logic [31:0] _RANDOM_594;
	logic [31:0] _RANDOM_595;
	logic [31:0] _RANDOM_596;
	logic [31:0] _RANDOM_597;
	logic [31:0] _RANDOM_598;
	logic [31:0] _RANDOM_599;
	logic [31:0] _RANDOM_600;
	logic [31:0] _RANDOM_601;
	logic [31:0] _RANDOM_602;
	logic [31:0] _RANDOM_603;
	logic [31:0] _RANDOM_604;
	logic [31:0] _RANDOM_605;
	logic [31:0] _RANDOM_606;
	logic [31:0] _RANDOM_607;
	logic [31:0] _RANDOM_608;
	logic [31:0] _RANDOM_609;
	logic [31:0] _RANDOM_610;
	logic [31:0] _RANDOM_611;
	logic [31:0] _RANDOM_612;
	logic [31:0] _RANDOM_613;
	logic [31:0] _RANDOM_614;
	logic [31:0] _RANDOM_615;
	logic [31:0] _RANDOM_616;
	logic [31:0] _RANDOM_617;
	logic [31:0] _RANDOM_618;
	logic [31:0] _RANDOM_619;
	logic [31:0] _RANDOM_620;
	logic [31:0] _RANDOM_621;
	logic [31:0] _RANDOM_622;
	logic [31:0] _RANDOM_623;
	logic [31:0] _RANDOM_624;
	logic [31:0] _RANDOM_625;
	logic [31:0] _RANDOM_626;
	logic [31:0] _RANDOM_627;
	logic [31:0] _RANDOM_628;
	logic [31:0] _RANDOM_629;
	logic [31:0] _RANDOM_630;
	logic [31:0] _RANDOM_631;
	logic [31:0] _RANDOM_632;
	logic [31:0] _RANDOM_633;
	logic [31:0] _RANDOM_634;
	logic [31:0] _RANDOM_635;
	logic [31:0] _RANDOM_636;
	logic [31:0] _RANDOM_637;
	logic [31:0] _RANDOM_638;
	logic [31:0] _RANDOM_639;
	logic [31:0] _RANDOM_640;
	logic [31:0] _RANDOM_641;
	logic [31:0] _RANDOM_642;
	logic [31:0] _RANDOM_643;
	logic [31:0] _RANDOM_644;
	logic [31:0] _RANDOM_645;
	logic [31:0] _RANDOM_646;
	logic [31:0] _RANDOM_647;
	logic [31:0] _RANDOM_648;
	logic [31:0] _RANDOM_649;
	logic [31:0] _RANDOM_650;
	logic [31:0] _RANDOM_651;
	logic [31:0] _RANDOM_652;
	logic [31:0] _RANDOM_653;
	logic [31:0] _RANDOM_654;
	logic [31:0] _RANDOM_655;
	logic [31:0] _RANDOM_656;
	logic [31:0] _RANDOM_657;
	logic [31:0] _RANDOM_658;
	logic [31:0] _RANDOM_659;
	logic [31:0] _RANDOM_660;
	logic [31:0] _RANDOM_661;
	logic [31:0] _RANDOM_662;
	logic [31:0] _RANDOM_663;
	logic [31:0] _RANDOM_664;
	logic [31:0] _RANDOM_665;
	logic [31:0] _RANDOM_666;
	logic [31:0] _RANDOM_667;
	logic [31:0] _RANDOM_668;
	logic [31:0] _RANDOM_669;
	logic [31:0] _RANDOM_670;
	logic [31:0] _RANDOM_671;
	logic [31:0] _RANDOM_672;
	logic [31:0] _RANDOM_673;
	logic [31:0] _RANDOM_674;
	logic [31:0] _RANDOM_675;
	logic [31:0] _RANDOM_676;
	logic [31:0] _RANDOM_677;
	logic [31:0] _RANDOM_678;
	logic [31:0] _RANDOM_679;
	logic [31:0] _RANDOM_680;
	logic [31:0] _RANDOM_681;
	logic [31:0] _RANDOM_682;
	logic [31:0] _RANDOM_683;
	logic [31:0] _RANDOM_684;
	logic [31:0] _RANDOM_685;
	logic [31:0] _RANDOM_686;
	logic [31:0] _RANDOM_687;
	logic [31:0] _RANDOM_688;
	logic [31:0] _RANDOM_689;
	logic [31:0] _RANDOM_690;
	logic [31:0] _RANDOM_691;
	logic [31:0] _RANDOM_692;
	logic [31:0] _RANDOM_693;
	logic [31:0] _RANDOM_694;
	logic [31:0] _RANDOM_695;
	logic [31:0] _RANDOM_696;
	logic [31:0] _RANDOM_697;
	logic [31:0] _RANDOM_698;
	logic [31:0] _RANDOM_699;
	logic [31:0] _RANDOM_700;
	logic [31:0] _RANDOM_701;
	logic [31:0] _RANDOM_702;
	logic [31:0] _RANDOM_703;
	logic [31:0] _RANDOM_704;
	logic [31:0] _RANDOM_705;
	logic [31:0] _RANDOM_706;
	logic [31:0] _RANDOM_707;
	logic [31:0] _RANDOM_708;
	logic [31:0] _RANDOM_709;
	logic [31:0] _RANDOM_710;
	logic [31:0] _RANDOM_711;
	logic [31:0] _RANDOM_712;
	logic [31:0] _RANDOM_713;
	logic [31:0] _RANDOM_714;
	logic [31:0] _RANDOM_715;
	logic [31:0] _RANDOM_716;
	logic [31:0] _RANDOM_717;
	logic [31:0] _RANDOM_718;
	logic [31:0] _RANDOM_719;
	logic [31:0] _RANDOM_720;
	logic [31:0] _RANDOM_721;
	logic [31:0] _RANDOM_722;
	logic [31:0] _RANDOM_723;
	logic [31:0] _RANDOM_724;
	logic [31:0] _RANDOM_725;
	logic [31:0] _RANDOM_726;
	logic [31:0] _RANDOM_727;
	logic [31:0] _RANDOM_728;
	logic [31:0] _RANDOM_729;
	logic [31:0] _RANDOM_730;
	logic [31:0] _RANDOM_731;
	logic [31:0] _RANDOM_732;
	logic [31:0] _RANDOM_733;
	logic [31:0] _RANDOM_734;
	logic [31:0] _RANDOM_735;
	logic [31:0] _RANDOM_736;
	logic [31:0] _RANDOM_737;
	logic [31:0] _RANDOM_738;
	logic [31:0] _RANDOM_739;
	logic [31:0] _RANDOM_740;
	logic [31:0] _RANDOM_741;
	logic [31:0] _RANDOM_742;
	logic [31:0] _RANDOM_743;
	logic [31:0] _RANDOM_744;
	logic [31:0] _RANDOM_745;
	logic [31:0] _RANDOM_746;
	logic [31:0] _RANDOM_747;
	logic [31:0] _RANDOM_748;
	logic [31:0] _RANDOM_749;
	logic [31:0] _RANDOM_750;
	logic [31:0] _RANDOM_751;
	logic [31:0] _RANDOM_752;
	logic [31:0] _RANDOM_753;
	logic [31:0] _RANDOM_754;
	logic [31:0] _RANDOM_755;
	logic [31:0] _RANDOM_756;
	logic [31:0] _RANDOM_757;
	logic [31:0] _RANDOM_758;
	logic [31:0] _RANDOM_759;
	logic [31:0] _RANDOM_760;
	logic [31:0] _RANDOM_761;
	logic [31:0] _RANDOM_762;
	logic [31:0] _RANDOM_763;
	logic [31:0] _RANDOM_764;
	logic [31:0] _RANDOM_765;
	logic [31:0] _RANDOM_766;
	logic [31:0] _RANDOM_767;
	logic [31:0] _RANDOM_768;
	logic [31:0] _RANDOM_769;
	logic [31:0] _RANDOM_770;
	logic [31:0] _RANDOM_771;
	logic [31:0] _RANDOM_772;
	logic [31:0] _RANDOM_773;
	logic [31:0] _RANDOM_774;
	logic [31:0] _RANDOM_775;
	logic [31:0] _RANDOM_776;
	logic [31:0] _RANDOM_777;
	logic [31:0] _RANDOM_778;
	logic [31:0] _RANDOM_779;
	logic [31:0] _RANDOM_780;
	logic [31:0] _RANDOM_781;
	logic [31:0] _RANDOM_782;
	logic [31:0] _RANDOM_783;
	logic [31:0] _RANDOM_784;
	logic [31:0] _RANDOM_785;
	logic [31:0] _RANDOM_786;
	logic [31:0] _RANDOM_787;
	logic [31:0] _RANDOM_788;
	logic [31:0] _RANDOM_789;
	logic [31:0] _RANDOM_790;
	logic [31:0] _RANDOM_791;
	logic [31:0] _RANDOM_792;
	logic [31:0] _RANDOM_793;
	logic [31:0] _RANDOM_794;
	logic [31:0] _RANDOM_795;
	logic [31:0] _RANDOM_796;
	logic [31:0] _RANDOM_797;
	logic [31:0] _RANDOM_798;
	logic [31:0] _RANDOM_799;
	logic [31:0] _RANDOM_800;
	logic [31:0] _RANDOM_801;
	logic [31:0] _RANDOM_802;
	logic [31:0] _RANDOM_803;
	logic [31:0] _RANDOM_804;
	logic [31:0] _RANDOM_805;
	logic [31:0] _RANDOM_806;
	logic [31:0] _RANDOM_807;
	logic [31:0] _RANDOM_808;
	logic [31:0] _RANDOM_809;
	logic [31:0] _RANDOM_810;
	logic [31:0] _RANDOM_811;
	logic [31:0] _RANDOM_812;
	logic [31:0] _RANDOM_813;
	logic [31:0] _RANDOM_814;
	logic [31:0] _RANDOM_815;
	logic [31:0] _RANDOM_816;
	logic [31:0] _RANDOM_817;
	logic [31:0] _RANDOM_818;
	logic [31:0] _RANDOM_819;
	logic [31:0] _RANDOM_820;
	logic [31:0] _RANDOM_821;
	logic [31:0] _RANDOM_822;
	logic [31:0] _RANDOM_823;
	logic [31:0] _RANDOM_824;
	logic [31:0] _RANDOM_825;
	logic [31:0] _RANDOM_826;
	logic [31:0] _RANDOM_827;
	logic [31:0] _RANDOM_828;
	logic [31:0] _RANDOM_829;
	logic [31:0] _RANDOM_830;
	logic [31:0] _RANDOM_831;
	logic [31:0] _RANDOM_832;
	logic [31:0] _RANDOM_833;
	logic [31:0] _RANDOM_834;
	logic [31:0] _RANDOM_835;
	logic [31:0] _RANDOM_836;
	logic [31:0] _RANDOM_837;
	logic [31:0] _RANDOM_838;
	logic [31:0] _RANDOM_839;
	logic [31:0] _RANDOM_840;
	logic [31:0] _RANDOM_841;
	logic [31:0] _RANDOM_842;
	logic [31:0] _RANDOM_843;
	logic [31:0] _RANDOM_844;
	logic [31:0] _RANDOM_845;
	logic [31:0] _RANDOM_846;
	logic [31:0] _RANDOM_847;
	logic [31:0] _RANDOM_848;
	logic [31:0] _RANDOM_849;
	logic [31:0] _RANDOM_850;
	logic [31:0] _RANDOM_851;
	logic [31:0] _RANDOM_852;
	logic [31:0] _RANDOM_853;
	logic [31:0] _RANDOM_854;
	logic [31:0] _RANDOM_855;
	logic [31:0] _RANDOM_856;
	logic [31:0] _RANDOM_857;
	logic [31:0] _RANDOM_858;
	logic [31:0] _RANDOM_859;
	logic [31:0] _RANDOM_860;
	logic [31:0] _RANDOM_861;
	logic [31:0] _RANDOM_862;
	logic [31:0] _RANDOM_863;
	logic [31:0] _RANDOM_864;
	logic [31:0] _RANDOM_865;
	logic [31:0] _RANDOM_866;
	logic [31:0] _RANDOM_867;
	logic [31:0] _RANDOM_868;
	logic [31:0] _RANDOM_869;
	logic [31:0] _RANDOM_870;
	logic [31:0] _RANDOM_871;
	logic [31:0] _RANDOM_872;
	logic [31:0] _RANDOM_873;
	logic [31:0] _RANDOM_874;
	logic [31:0] _RANDOM_875;
	logic [31:0] _RANDOM_876;
	logic [31:0] _RANDOM_877;
	logic [31:0] _RANDOM_878;
	logic [31:0] _RANDOM_879;
	logic [31:0] _RANDOM_880;
	logic [31:0] _RANDOM_881;
	logic [31:0] _RANDOM_882;
	logic [31:0] _RANDOM_883;
	logic [31:0] _RANDOM_884;
	logic [31:0] _RANDOM_885;
	logic [31:0] _RANDOM_886;
	logic [31:0] _RANDOM_887;
	logic [31:0] _RANDOM_888;
	logic [31:0] _RANDOM_889;
	logic [31:0] _RANDOM_890;
	logic [31:0] _RANDOM_891;
	logic [31:0] _RANDOM_892;
	logic [31:0] _RANDOM_893;
	logic [31:0] _RANDOM_894;
	logic [31:0] _RANDOM_895;
	logic [31:0] _RANDOM_896;
	logic [31:0] _RANDOM_897;
	logic [31:0] _RANDOM_898;
	logic [31:0] _RANDOM_899;
	logic [31:0] _RANDOM_900;
	logic [31:0] _RANDOM_901;
	logic [31:0] _RANDOM_902;
	logic [31:0] _RANDOM_903;
	logic [31:0] _RANDOM_904;
	logic [31:0] _RANDOM_905;
	logic [31:0] _RANDOM_906;
	logic [31:0] _RANDOM_907;
	logic [31:0] _RANDOM_908;
	logic [31:0] _RANDOM_909;
	logic [31:0] _RANDOM_910;
	logic [31:0] _RANDOM_911;
	logic [31:0] _RANDOM_912;
	logic [31:0] _RANDOM_913;
	logic [31:0] _RANDOM_914;
	logic [31:0] _RANDOM_915;
	logic [31:0] _RANDOM_916;
	logic [31:0] _RANDOM_917;
	logic [31:0] _RANDOM_918;
	logic [31:0] _RANDOM_919;
	logic [31:0] _RANDOM_920;
	logic [31:0] _RANDOM_921;
	logic [31:0] _RANDOM_922;
	logic [31:0] _RANDOM_923;
	logic [31:0] _RANDOM_924;
	logic [31:0] _RANDOM_925;
	logic [31:0] _RANDOM_926;
	logic [31:0] _RANDOM_927;
	logic [31:0] _RANDOM_928;
	logic [31:0] _RANDOM_929;
	logic [31:0] _RANDOM_930;
	logic [31:0] _RANDOM_931;
	logic [31:0] _RANDOM_932;
	logic [31:0] _RANDOM_933;
	logic [31:0] _RANDOM_934;
	logic [31:0] _RANDOM_935;
	logic [31:0] _RANDOM_936;
	logic [31:0] _RANDOM_937;
	logic [31:0] _RANDOM_938;
	logic [31:0] _RANDOM_939;
	logic [31:0] _RANDOM_940;
	logic [31:0] _RANDOM_941;
	logic [31:0] _RANDOM_942;
	logic [31:0] _RANDOM_943;
	logic [31:0] _RANDOM_944;
	logic [31:0] _RANDOM_945;
	logic [31:0] _RANDOM_946;
	logic [31:0] _RANDOM_947;
	logic [31:0] _RANDOM_948;
	logic [31:0] _RANDOM_949;
	logic [31:0] _RANDOM_950;
	logic [31:0] _RANDOM_951;
	logic [31:0] _RANDOM_952;
	logic [31:0] _RANDOM_953;
	logic [31:0] _RANDOM_954;
	logic [31:0] _RANDOM_955;
	logic [31:0] _RANDOM_956;
	logic [31:0] _RANDOM_957;
	logic [31:0] _RANDOM_958;
	logic [31:0] _RANDOM_959;
	logic [31:0] _RANDOM_960;
	logic [31:0] _RANDOM_961;
	logic [31:0] _RANDOM_962;
	logic [31:0] _RANDOM_963;
	logic [31:0] _RANDOM_964;
	logic [31:0] _RANDOM_965;
	logic [31:0] _RANDOM_966;
	logic [31:0] _RANDOM_967;
	logic [31:0] _RANDOM_968;
	logic [31:0] _RANDOM_969;
	logic [31:0] _RANDOM_970;
	logic [31:0] _RANDOM_971;
	logic [31:0] _RANDOM_972;
	logic [31:0] _RANDOM_973;
	logic [31:0] _RANDOM_974;
	logic [31:0] _RANDOM_975;
	logic [31:0] _RANDOM_976;
	logic [31:0] _RANDOM_977;
	logic [31:0] _RANDOM_978;
	logic [31:0] _RANDOM_979;
	logic [31:0] _RANDOM_980;
	logic [31:0] _RANDOM_981;
	logic [31:0] _RANDOM_982;
	logic [31:0] _RANDOM_983;
	logic [31:0] _RANDOM_984;
	logic [31:0] _RANDOM_985;
	logic [31:0] _RANDOM_986;
	logic [31:0] _RANDOM_987;
	logic [31:0] _RANDOM_988;
	logic [31:0] _RANDOM_989;
	logic [31:0] _RANDOM_990;
	logic [31:0] _RANDOM_991;
	logic [31:0] _RANDOM_992;
	logic [31:0] _RANDOM_993;
	logic [31:0] _RANDOM_994;
	logic [31:0] _RANDOM_995;
	logic [31:0] _RANDOM_996;
	logic [31:0] _RANDOM_997;
	logic [31:0] _RANDOM_998;
	logic [31:0] _RANDOM_999;
	logic [31:0] _RANDOM_1000;
	logic [31:0] _RANDOM_1001;
	logic [31:0] _RANDOM_1002;
	logic [31:0] _RANDOM_1003;
	logic [31:0] _RANDOM_1004;
	logic [31:0] _RANDOM_1005;
	logic [31:0] _RANDOM_1006;
	logic [31:0] _RANDOM_1007;
	logic [31:0] _RANDOM_1008;
	logic [31:0] _RANDOM_1009;
	logic [31:0] _RANDOM_1010;
	logic [31:0] _RANDOM_1011;
	logic [31:0] _RANDOM_1012;
	logic [31:0] _RANDOM_1013;
	logic [31:0] _RANDOM_1014;
	logic [31:0] _RANDOM_1015;
	logic [31:0] _RANDOM_1016;
	logic [31:0] _RANDOM_1017;
	logic [31:0] _RANDOM_1018;
	logic [31:0] _RANDOM_1019;
	logic [31:0] _RANDOM_1020;
	logic [31:0] _RANDOM_1021;
	logic [31:0] _RANDOM_1022;
	logic [31:0] _RANDOM_1023;
	logic [31:0] _RANDOM_1024;
	logic [31:0] _RANDOM_1025;
	logic [31:0] _RANDOM_1026;
	logic [31:0] _RANDOM_1027;
	logic [31:0] _RANDOM_1028;
	logic [31:0] _RANDOM_1029;
	logic [31:0] _RANDOM_1030;
	logic [31:0] _RANDOM_1031;
	logic [31:0] _RANDOM_1032;
	logic [31:0] _RANDOM_1033;
	logic [31:0] _RANDOM_1034;
	logic [31:0] _RANDOM_1035;
	logic [31:0] _RANDOM_1036;
	logic [31:0] _RANDOM_1037;
	logic [31:0] _RANDOM_1038;
	logic [31:0] _RANDOM_1039;
	logic [31:0] _RANDOM_1040;
	logic [31:0] _RANDOM_1041;
	logic [31:0] _RANDOM_1042;
	logic [31:0] _RANDOM_1043;
	logic [31:0] _RANDOM_1044;
	logic [31:0] _RANDOM_1045;
	logic [31:0] _RANDOM_1046;
	logic [31:0] _RANDOM_1047;
	logic [31:0] _RANDOM_1048;
	logic [31:0] _RANDOM_1049;
	logic [31:0] _RANDOM_1050;
	logic [31:0] _RANDOM_1051;
	logic [31:0] _RANDOM_1052;
	logic [31:0] _RANDOM_1053;
	logic [31:0] _RANDOM_1054;
	logic [31:0] _RANDOM_1055;
	logic [31:0] _RANDOM_1056;
	logic [31:0] _RANDOM_1057;
	logic [31:0] _RANDOM_1058;
	logic [31:0] _RANDOM_1059;
	logic [31:0] _RANDOM_1060;
	logic [31:0] _RANDOM_1061;
	logic [31:0] _RANDOM_1062;
	logic [31:0] _RANDOM_1063;
	logic [31:0] _RANDOM_1064;
	logic [31:0] _RANDOM_1065;
	logic [31:0] _RANDOM_1066;
	logic [31:0] _RANDOM_1067;
	logic [31:0] _RANDOM_1068;
	logic [31:0] _RANDOM_1069;
	logic [31:0] _RANDOM_1070;
	logic [31:0] _RANDOM_1071;
	logic [31:0] _RANDOM_1072;
	logic [31:0] _RANDOM_1073;
	logic [31:0] _RANDOM_1074;
	logic [31:0] _RANDOM_1075;
	logic [31:0] _RANDOM_1076;
	logic [31:0] _RANDOM_1077;
	logic [31:0] _RANDOM_1078;
	logic [31:0] _RANDOM_1079;
	logic [31:0] _RANDOM_1080;
	logic [31:0] _RANDOM_1081;
	logic [31:0] _RANDOM_1082;
	logic [31:0] _RANDOM_1083;
	logic [31:0] _RANDOM_1084;
	logic [31:0] _RANDOM_1085;
	logic [31:0] _RANDOM_1086;
	logic [31:0] _RANDOM_1087;
	logic [31:0] _RANDOM_1088;
	logic [31:0] _RANDOM_1089;
	logic [31:0] _RANDOM_1090;
	logic [31:0] _RANDOM_1091;
	logic [31:0] _RANDOM_1092;
	logic [31:0] _RANDOM_1093;
	logic [31:0] _RANDOM_1094;
	logic [31:0] _RANDOM_1095;
	logic [31:0] _RANDOM_1096;
	logic [31:0] _RANDOM_1097;
	logic [31:0] _RANDOM_1098;
	logic [31:0] _RANDOM_1099;
	logic [31:0] _RANDOM_1100;
	logic [31:0] _RANDOM_1101;
	logic [31:0] _RANDOM_1102;
	logic [31:0] _RANDOM_1103;
	logic [31:0] _RANDOM_1104;
	logic [31:0] _RANDOM_1105;
	logic [31:0] _RANDOM_1106;
	logic [31:0] _RANDOM_1107;
	logic [31:0] _RANDOM_1108;
	logic [31:0] _RANDOM_1109;
	logic [31:0] _RANDOM_1110;
	logic [31:0] _RANDOM_1111;
	logic [31:0] _RANDOM_1112;
	logic [31:0] _RANDOM_1113;
	logic [31:0] _RANDOM_1114;
	logic [31:0] _RANDOM_1115;
	logic [31:0] _RANDOM_1116;
	logic [31:0] _RANDOM_1117;
	logic [31:0] _RANDOM_1118;
	logic [31:0] _RANDOM_1119;
	logic [31:0] _RANDOM_1120;
	logic [31:0] _RANDOM_1121;
	logic [31:0] _RANDOM_1122;
	logic [31:0] _RANDOM_1123;
	logic [31:0] _RANDOM_1124;
	logic [31:0] _RANDOM_1125;
	logic [31:0] _RANDOM_1126;
	logic [31:0] _RANDOM_1127;
	logic [31:0] _RANDOM_1128;
	logic [31:0] _RANDOM_1129;
	logic [31:0] _RANDOM_1130;
	logic [31:0] _RANDOM_1131;
	logic [31:0] _RANDOM_1132;
	logic [31:0] _RANDOM_1133;
	logic [31:0] _RANDOM_1134;
	logic [31:0] _RANDOM_1135;
	logic [31:0] _RANDOM_1136;
	logic [31:0] _RANDOM_1137;
	logic [31:0] _RANDOM_1138;
	logic [31:0] _RANDOM_1139;
	logic [31:0] _RANDOM_1140;
	logic [31:0] _RANDOM_1141;
	logic [31:0] _RANDOM_1142;
	logic [31:0] _RANDOM_1143;
	logic [31:0] _RANDOM_1144;
	logic [31:0] _RANDOM_1145;
	logic [31:0] _RANDOM_1146;
	logic [31:0] _RANDOM_1147;
	logic [31:0] _RANDOM_1148;
	logic [31:0] _RANDOM_1149;
	logic [31:0] _RANDOM_1150;
	logic [31:0] _RANDOM_1151;
	logic [31:0] _RANDOM_1152;
	logic [31:0] _RANDOM_1153;
	logic [31:0] _RANDOM_1154;
	logic [31:0] _RANDOM_1155;
	logic [31:0] _RANDOM_1156;
	logic [31:0] _RANDOM_1157;
	logic [31:0] _RANDOM_1158;
	logic [31:0] _RANDOM_1159;
	logic [31:0] _RANDOM_1160;
	logic [31:0] _RANDOM_1161;
	logic [31:0] _RANDOM_1162;
	logic [31:0] _RANDOM_1163;
	logic [31:0] _RANDOM_1164;
	logic [31:0] _RANDOM_1165;
	logic [31:0] _RANDOM_1166;
	logic [31:0] _RANDOM_1167;
	logic [31:0] _RANDOM_1168;
	logic [31:0] _RANDOM_1169;
	logic [31:0] _RANDOM_1170;
	logic [31:0] _RANDOM_1171;
	logic [31:0] _RANDOM_1172;
	logic [31:0] _RANDOM_1173;
	logic [31:0] _RANDOM_1174;
	logic [31:0] _RANDOM_1175;
	logic [31:0] _RANDOM_1176;
	logic [31:0] _RANDOM_1177;
	logic [31:0] _RANDOM_1178;
	logic [31:0] _RANDOM_1179;
	logic [31:0] _RANDOM_1180;
	logic [31:0] _RANDOM_1181;
	logic [31:0] _RANDOM_1182;
	logic [31:0] _RANDOM_1183;
	logic [31:0] _RANDOM_1184;
	logic [31:0] _RANDOM_1185;
	logic [31:0] _RANDOM_1186;
	logic [31:0] _RANDOM_1187;
	logic [31:0] _RANDOM_1188;
	logic [31:0] _RANDOM_1189;
	logic [31:0] _RANDOM_1190;
	logic [31:0] _RANDOM_1191;
	logic [31:0] _RANDOM_1192;
	logic [31:0] _RANDOM_1193;
	logic [31:0] _RANDOM_1194;
	logic [31:0] _RANDOM_1195;
	logic [31:0] _RANDOM_1196;
	logic [31:0] _RANDOM_1197;
	logic [31:0] _RANDOM_1198;
	logic [31:0] _RANDOM_1199;
	logic [31:0] _RANDOM_1200;
	logic [31:0] _RANDOM_1201;
	logic [31:0] _RANDOM_1202;
	logic [31:0] _RANDOM_1203;
	logic [31:0] _RANDOM_1204;
	logic [31:0] _RANDOM_1205;
	logic [31:0] _RANDOM_1206;
	logic [31:0] _RANDOM_1207;
	logic [31:0] _RANDOM_1208;
	logic [31:0] _RANDOM_1209;
	logic [31:0] _RANDOM_1210;
	logic [31:0] _RANDOM_1211;
	logic [31:0] _RANDOM_1212;
	logic [31:0] _RANDOM_1213;
	logic [31:0] _RANDOM_1214;
	logic [31:0] _RANDOM_1215;
	logic [31:0] _RANDOM_1216;
	logic [31:0] _RANDOM_1217;
	logic [31:0] _RANDOM_1218;
	logic [31:0] _RANDOM_1219;
	logic [31:0] _RANDOM_1220;
	logic [31:0] _RANDOM_1221;
	logic [31:0] _RANDOM_1222;
	logic [31:0] _RANDOM_1223;
	logic [31:0] _RANDOM_1224;
	logic [31:0] _RANDOM_1225;
	logic [31:0] _RANDOM_1226;
	logic [31:0] _RANDOM_1227;
	logic [31:0] _RANDOM_1228;
	logic [31:0] _RANDOM_1229;
	logic [31:0] _RANDOM_1230;
	logic [31:0] _RANDOM_1231;
	logic [31:0] _RANDOM_1232;
	logic [31:0] _RANDOM_1233;
	logic [31:0] _RANDOM_1234;
	logic [31:0] _RANDOM_1235;
	logic [31:0] _RANDOM_1236;
	logic [31:0] _RANDOM_1237;
	logic [31:0] _RANDOM_1238;
	logic [31:0] _RANDOM_1239;
	logic [31:0] _RANDOM_1240;
	logic [31:0] _RANDOM_1241;
	logic [31:0] _RANDOM_1242;
	logic [31:0] _RANDOM_1243;
	logic [31:0] _RANDOM_1244;
	logic [31:0] _RANDOM_1245;
	logic [31:0] _RANDOM_1246;
	logic [31:0] _RANDOM_1247;
	logic [31:0] _RANDOM_1248;
	logic [31:0] _RANDOM_1249;
	logic [31:0] _RANDOM_1250;
	logic [31:0] _RANDOM_1251;
	logic [31:0] _RANDOM_1252;
	logic [31:0] _RANDOM_1253;
	logic [31:0] _RANDOM_1254;
	logic [31:0] _RANDOM_1255;
	logic [31:0] _RANDOM_1256;
	logic [31:0] _RANDOM_1257;
	logic [31:0] _RANDOM_1258;
	logic [31:0] _RANDOM_1259;
	logic [31:0] _RANDOM_1260;
	logic [31:0] _RANDOM_1261;
	logic [31:0] _RANDOM_1262;
	logic [31:0] _RANDOM_1263;
	logic [31:0] _RANDOM_1264;
	logic [31:0] _RANDOM_1265;
	logic [31:0] _RANDOM_1266;
	logic [31:0] _RANDOM_1267;
	logic [31:0] _RANDOM_1268;
	logic [31:0] _RANDOM_1269;
	logic [31:0] _RANDOM_1270;
	logic [31:0] _RANDOM_1271;
	logic [31:0] _RANDOM_1272;
	logic [31:0] _RANDOM_1273;
	logic [31:0] _RANDOM_1274;
	logic [31:0] _RANDOM_1275;
	logic [31:0] _RANDOM_1276;
	logic [31:0] _RANDOM_1277;
	logic [31:0] _RANDOM_1278;
	logic [31:0] _RANDOM_1279;
	logic [31:0] _RANDOM_1280;
	logic [31:0] _RANDOM_1281;
	logic [31:0] _RANDOM_1282;
	logic [31:0] _RANDOM_1283;
	logic [31:0] _RANDOM_1284;
	logic [31:0] _RANDOM_1285;
	logic [31:0] _RANDOM_1286;
	logic [31:0] _RANDOM_1287;
	logic [31:0] _RANDOM_1288;
	logic [31:0] _RANDOM_1289;
	logic [31:0] _RANDOM_1290;
	logic [31:0] _RANDOM_1291;
	logic [31:0] _RANDOM_1292;
	logic [31:0] _RANDOM_1293;
	logic [31:0] _RANDOM_1294;
	logic [31:0] _RANDOM_1295;
	logic [31:0] _RANDOM_1296;
	logic [31:0] _RANDOM_1297;
	logic [31:0] _RANDOM_1298;
	logic [31:0] _RANDOM_1299;
	logic [31:0] _RANDOM_1300;
	logic [31:0] _RANDOM_1301;
	logic [31:0] _RANDOM_1302;
	logic [31:0] _RANDOM_1303;
	logic [31:0] _RANDOM_1304;
	logic [31:0] _RANDOM_1305;
	logic [31:0] _RANDOM_1306;
	logic [31:0] _RANDOM_1307;
	logic [31:0] _RANDOM_1308;
	logic [31:0] _RANDOM_1309;
	logic [31:0] _RANDOM_1310;
	logic [31:0] _RANDOM_1311;
	logic [31:0] _RANDOM_1312;
	logic [31:0] _RANDOM_1313;
	logic [31:0] _RANDOM_1314;
	logic [31:0] _RANDOM_1315;
	logic [31:0] _RANDOM_1316;
	logic [31:0] _RANDOM_1317;
	logic [31:0] _RANDOM_1318;
	logic [31:0] _RANDOM_1319;
	logic [31:0] _RANDOM_1320;
	logic [31:0] _RANDOM_1321;
	logic [31:0] _RANDOM_1322;
	logic [31:0] _RANDOM_1323;
	logic [31:0] _RANDOM_1324;
	logic [31:0] _RANDOM_1325;
	logic [31:0] _RANDOM_1326;
	logic [31:0] _RANDOM_1327;
	logic [31:0] _RANDOM_1328;
	logic [31:0] _RANDOM_1329;
	logic [31:0] _RANDOM_1330;
	logic [31:0] _RANDOM_1331;
	logic [31:0] _RANDOM_1332;
	logic [31:0] _RANDOM_1333;
	logic [31:0] _RANDOM_1334;
	logic [31:0] _RANDOM_1335;
	logic [31:0] _RANDOM_1336;
	logic [31:0] _RANDOM_1337;
	logic [31:0] _RANDOM_1338;
	logic [31:0] _RANDOM_1339;
	logic [31:0] _RANDOM_1340;
	logic [31:0] _RANDOM_1341;
	logic [31:0] _RANDOM_1342;
	logic [31:0] _RANDOM_1343;
	logic [31:0] _RANDOM_1344;
	logic [31:0] _RANDOM_1345;
	logic [31:0] _RANDOM_1346;
	logic [31:0] _RANDOM_1347;
	logic [31:0] _RANDOM_1348;
	logic [31:0] _RANDOM_1349;
	logic [31:0] _RANDOM_1350;
	logic [31:0] _RANDOM_1351;
	logic [31:0] _RANDOM_1352;
	logic [31:0] _RANDOM_1353;
	logic [31:0] _RANDOM_1354;
	logic [31:0] _RANDOM_1355;
	logic [31:0] _RANDOM_1356;
	logic [31:0] _RANDOM_1357;
	logic [31:0] _RANDOM_1358;
	logic [31:0] _RANDOM_1359;
	logic [31:0] _RANDOM_1360;
	logic [31:0] _RANDOM_1361;
	logic [31:0] _RANDOM_1362;
	logic [31:0] _RANDOM_1363;
	logic [31:0] _RANDOM_1364;
	logic [31:0] _RANDOM_1365;
	logic [31:0] _RANDOM_1366;
	logic [31:0] _RANDOM_1367;
	logic [31:0] _RANDOM_1368;
	logic [31:0] _RANDOM_1369;
	logic [31:0] _RANDOM_1370;
	logic [31:0] _RANDOM_1371;
	logic [31:0] _RANDOM_1372;
	logic [31:0] _RANDOM_1373;
	logic [31:0] _RANDOM_1374;
	logic [31:0] _RANDOM_1375;
	logic [31:0] _RANDOM_1376;
	logic [31:0] _RANDOM_1377;
	logic [31:0] _RANDOM_1378;
	logic [31:0] _RANDOM_1379;
	logic [31:0] _RANDOM_1380;
	logic [31:0] _RANDOM_1381;
	logic [31:0] _RANDOM_1382;
	logic [31:0] _RANDOM_1383;
	logic [31:0] _RANDOM_1384;
	logic [31:0] _RANDOM_1385;
	logic [31:0] _RANDOM_1386;
	logic [31:0] _RANDOM_1387;
	logic [31:0] _RANDOM_1388;
	logic [31:0] _RANDOM_1389;
	logic [31:0] _RANDOM_1390;
	logic [31:0] _RANDOM_1391;
	logic [31:0] _RANDOM_1392;
	logic [31:0] _RANDOM_1393;
	logic [31:0] _RANDOM_1394;
	logic [31:0] _RANDOM_1395;
	logic [31:0] _RANDOM_1396;
	logic [31:0] _RANDOM_1397;
	logic [31:0] _RANDOM_1398;
	logic [31:0] _RANDOM_1399;
	logic [31:0] _RANDOM_1400;
	logic [31:0] _RANDOM_1401;
	logic [31:0] _RANDOM_1402;
	logic [31:0] _RANDOM_1403;
	logic [31:0] _RANDOM_1404;
	logic [31:0] _RANDOM_1405;
	logic [31:0] _RANDOM_1406;
	logic [31:0] _RANDOM_1407;
	logic [31:0] _RANDOM_1408;
	logic [31:0] _RANDOM_1409;
	logic [31:0] _RANDOM_1410;
	logic [31:0] _RANDOM_1411;
	logic [31:0] _RANDOM_1412;
	logic [31:0] _RANDOM_1413;
	logic [31:0] _RANDOM_1414;
	logic [31:0] _RANDOM_1415;
	logic [31:0] _RANDOM_1416;
	logic [31:0] _RANDOM_1417;
	logic [31:0] _RANDOM_1418;
	logic [31:0] _RANDOM_1419;
	logic [31:0] _RANDOM_1420;
	logic [31:0] _RANDOM_1421;
	logic [31:0] _RANDOM_1422;
	logic [31:0] _RANDOM_1423;
	logic [31:0] _RANDOM_1424;
	logic [31:0] _RANDOM_1425;
	logic [31:0] _RANDOM_1426;
	logic [31:0] _RANDOM_1427;
	logic [31:0] _RANDOM_1428;
	logic [31:0] _RANDOM_1429;
	logic [31:0] _RANDOM_1430;
	logic [31:0] _RANDOM_1431;
	logic [31:0] _RANDOM_1432;
	logic [31:0] _RANDOM_1433;
	logic [31:0] _RANDOM_1434;
	logic [31:0] _RANDOM_1435;
	logic [31:0] _RANDOM_1436;
	logic [31:0] _RANDOM_1437;
	logic [31:0] _RANDOM_1438;
	logic [31:0] _RANDOM_1439;
	logic [31:0] _RANDOM_1440;
	logic [31:0] _RANDOM_1441;
	logic [31:0] _RANDOM_1442;
	logic [31:0] _RANDOM_1443;
	logic [31:0] _RANDOM_1444;
	logic [31:0] _RANDOM_1445;
	logic [31:0] _RANDOM_1446;
	logic [31:0] _RANDOM_1447;
	logic [31:0] _RANDOM_1448;
	logic [31:0] _RANDOM_1449;
	logic [31:0] _RANDOM_1450;
	logic [31:0] _RANDOM_1451;
	logic [31:0] _RANDOM_1452;
	logic [31:0] _RANDOM_1453;
	logic [31:0] _RANDOM_1454;
	logic [31:0] _RANDOM_1455;
	logic [31:0] _RANDOM_1456;
	logic [31:0] _RANDOM_1457;
	logic [31:0] _RANDOM_1458;
	logic [31:0] _RANDOM_1459;
	logic [31:0] _RANDOM_1460;
	logic [31:0] _RANDOM_1461;
	logic [31:0] _RANDOM_1462;
	logic [31:0] _RANDOM_1463;
	logic [31:0] _RANDOM_1464;
	logic [31:0] _RANDOM_1465;
	logic [31:0] _RANDOM_1466;
	logic [31:0] _RANDOM_1467;
	logic [31:0] _RANDOM_1468;
	logic [31:0] _RANDOM_1469;
	logic [31:0] _RANDOM_1470;
	logic [31:0] _RANDOM_1471;
	logic [31:0] _RANDOM_1472;
	logic [31:0] _RANDOM_1473;
	logic [31:0] _RANDOM_1474;
	logic [31:0] _RANDOM_1475;
	logic [31:0] _RANDOM_1476;
	logic [31:0] _RANDOM_1477;
	logic [31:0] _RANDOM_1478;
	logic [31:0] _RANDOM_1479;
	logic [31:0] _RANDOM_1480;
	logic [31:0] _RANDOM_1481;
	logic [31:0] _RANDOM_1482;
	logic [31:0] _RANDOM_1483;
	logic [31:0] _RANDOM_1484;
	logic [31:0] _RANDOM_1485;
	logic [31:0] _RANDOM_1486;
	logic [31:0] _RANDOM_1487;
	logic [31:0] _RANDOM_1488;
	logic [31:0] _RANDOM_1489;
	logic [31:0] _RANDOM_1490;
	logic [31:0] _RANDOM_1491;
	logic [31:0] _RANDOM_1492;
	logic [31:0] _RANDOM_1493;
	logic [31:0] _RANDOM_1494;
	logic [31:0] _RANDOM_1495;
	logic [31:0] _RANDOM_1496;
	logic [31:0] _RANDOM_1497;
	logic [31:0] _RANDOM_1498;
	logic [31:0] _RANDOM_1499;
	logic [31:0] _RANDOM_1500;
	logic [31:0] _RANDOM_1501;
	logic [31:0] _RANDOM_1502;
	logic [31:0] _RANDOM_1503;
	logic [31:0] _RANDOM_1504;
	logic [31:0] _RANDOM_1505;
	logic [31:0] _RANDOM_1506;
	logic [31:0] _RANDOM_1507;
	logic [31:0] _RANDOM_1508;
	logic [31:0] _RANDOM_1509;
	logic [31:0] _RANDOM_1510;
	logic [31:0] _RANDOM_1511;
	logic [31:0] _RANDOM_1512;
	logic [31:0] _RANDOM_1513;
	logic [31:0] _RANDOM_1514;
	logic [31:0] _RANDOM_1515;
	logic [31:0] _RANDOM_1516;
	logic [31:0] _RANDOM_1517;
	logic [31:0] _RANDOM_1518;
	logic [31:0] _RANDOM_1519;
	logic [31:0] _RANDOM_1520;
	logic [31:0] _RANDOM_1521;
	logic [31:0] _RANDOM_1522;
	logic [31:0] _RANDOM_1523;
	logic [31:0] _RANDOM_1524;
	logic [31:0] _RANDOM_1525;
	logic [31:0] _RANDOM_1526;
	logic [31:0] _RANDOM_1527;
	logic [31:0] _RANDOM_1528;
	logic [31:0] _RANDOM_1529;
	logic [31:0] _RANDOM_1530;
	logic [31:0] _RANDOM_1531;
	logic [31:0] _RANDOM_1532;
	logic [31:0] _RANDOM_1533;
	logic [31:0] _RANDOM_1534;
	logic [31:0] _RANDOM_1535;
	logic [31:0] _RANDOM_1536;
	logic [31:0] _RANDOM_1537;
	logic [31:0] _RANDOM_1538;
	logic [31:0] _RANDOM_1539;
	logic [31:0] _RANDOM_1540;
	logic [31:0] _RANDOM_1541;
	logic [31:0] _RANDOM_1542;
	logic [31:0] _RANDOM_1543;
	logic [31:0] _RANDOM_1544;
	logic [31:0] _RANDOM_1545;
	logic [31:0] _RANDOM_1546;
	logic [31:0] _RANDOM_1547;
	logic [31:0] _RANDOM_1548;
	logic [31:0] _RANDOM_1549;
	logic [31:0] _RANDOM_1550;
	logic [31:0] _RANDOM_1551;
	logic [31:0] _RANDOM_1552;
	logic [31:0] _RANDOM_1553;
	logic [31:0] _RANDOM_1554;
	logic [31:0] _RANDOM_1555;
	logic [31:0] _RANDOM_1556;
	logic [31:0] _RANDOM_1557;
	logic [31:0] _RANDOM_1558;
	logic [31:0] _RANDOM_1559;
	logic [31:0] _RANDOM_1560;
	logic [31:0] _RANDOM_1561;
	logic [31:0] _RANDOM_1562;
	logic [31:0] _RANDOM_1563;
	logic [31:0] _RANDOM_1564;
	logic [31:0] _RANDOM_1565;
	logic [31:0] _RANDOM_1566;
	logic [31:0] _RANDOM_1567;
	logic [31:0] _RANDOM_1568;
	logic [31:0] _RANDOM_1569;
	logic [31:0] _RANDOM_1570;
	logic [31:0] _RANDOM_1571;
	logic [31:0] _RANDOM_1572;
	logic [31:0] _RANDOM_1573;
	logic [31:0] _RANDOM_1574;
	logic [31:0] _RANDOM_1575;
	logic [31:0] _RANDOM_1576;
	logic [31:0] _RANDOM_1577;
	logic [31:0] _RANDOM_1578;
	logic [31:0] _RANDOM_1579;
	logic [31:0] _RANDOM_1580;
	logic [31:0] _RANDOM_1581;
	logic [31:0] _RANDOM_1582;
	logic [31:0] _RANDOM_1583;
	logic [31:0] _RANDOM_1584;
	logic [31:0] _RANDOM_1585;
	logic [31:0] _RANDOM_1586;
	logic [31:0] _RANDOM_1587;
	logic [31:0] _RANDOM_1588;
	logic [31:0] _RANDOM_1589;
	logic [31:0] _RANDOM_1590;
	logic [31:0] _RANDOM_1591;
	logic [31:0] _RANDOM_1592;
	logic [31:0] _RANDOM_1593;
	logic [31:0] _RANDOM_1594;
	logic [31:0] _RANDOM_1595;
	logic [31:0] _RANDOM_1596;
	logic [31:0] _RANDOM_1597;
	logic [31:0] _RANDOM_1598;
	logic [31:0] _RANDOM_1599;
	logic [31:0] _RANDOM_1600;
	logic [31:0] _RANDOM_1601;
	logic [31:0] _RANDOM_1602;
	logic [31:0] _RANDOM_1603;
	logic [31:0] _RANDOM_1604;
	logic [31:0] _RANDOM_1605;
	logic [31:0] _RANDOM_1606;
	logic [31:0] _RANDOM_1607;
	logic [31:0] _RANDOM_1608;
	logic [31:0] _RANDOM_1609;
	logic [31:0] _RANDOM_1610;
	logic [31:0] _RANDOM_1611;
	logic [31:0] _RANDOM_1612;
	logic [31:0] _RANDOM_1613;
	logic [31:0] _RANDOM_1614;
	logic [31:0] _RANDOM_1615;
	logic [31:0] _RANDOM_1616;
	logic [31:0] _RANDOM_1617;
	logic [31:0] _RANDOM_1618;
	logic [31:0] _RANDOM_1619;
	logic [31:0] _RANDOM_1620;
	logic [31:0] _RANDOM_1621;
	logic [31:0] _RANDOM_1622;
	logic [31:0] _RANDOM_1623;
	logic [31:0] _RANDOM_1624;
	logic [31:0] _RANDOM_1625;
	logic [31:0] _RANDOM_1626;
	logic [31:0] _RANDOM_1627;
	logic [31:0] _RANDOM_1628;
	logic [31:0] _RANDOM_1629;
	logic [31:0] _RANDOM_1630;
	logic [31:0] _RANDOM_1631;
	logic [31:0] _RANDOM_1632;
	logic [31:0] _RANDOM_1633;
	logic [31:0] _RANDOM_1634;
	logic [31:0] _RANDOM_1635;
	logic [31:0] _RANDOM_1636;
	logic [31:0] _RANDOM_1637;
	logic [31:0] _RANDOM_1638;
	logic [31:0] _RANDOM_1639;
	logic [31:0] _RANDOM_1640;
	logic [31:0] _RANDOM_1641;
	logic [31:0] _RANDOM_1642;
	logic [31:0] _RANDOM_1643;
	logic [31:0] _RANDOM_1644;
	logic [31:0] _RANDOM_1645;
	logic [31:0] _RANDOM_1646;
	logic [31:0] _RANDOM_1647;
	logic [31:0] _RANDOM_1648;
	logic [31:0] _RANDOM_1649;
	logic [31:0] _RANDOM_1650;
	logic [31:0] _RANDOM_1651;
	logic [31:0] _RANDOM_1652;
	logic [31:0] _RANDOM_1653;
	logic [31:0] _RANDOM_1654;
	logic [31:0] _RANDOM_1655;
	logic [31:0] _RANDOM_1656;
	logic [31:0] _RANDOM_1657;
	logic [31:0] _RANDOM_1658;
	logic [31:0] _RANDOM_1659;
	logic [31:0] _RANDOM_1660;
	logic [31:0] _RANDOM_1661;
	logic [31:0] _RANDOM_1662;
	logic [31:0] _RANDOM_1663;
	logic [31:0] _RANDOM_1664;
	logic [31:0] _RANDOM_1665;
	logic [31:0] _RANDOM_1666;
	logic [31:0] _RANDOM_1667;
	logic [31:0] _RANDOM_1668;
	logic [31:0] _RANDOM_1669;
	logic [31:0] _RANDOM_1670;
	logic [31:0] _RANDOM_1671;
	logic [31:0] _RANDOM_1672;
	logic [31:0] _RANDOM_1673;
	logic [31:0] _RANDOM_1674;
	logic [31:0] _RANDOM_1675;
	logic [31:0] _RANDOM_1676;
	logic [31:0] _RANDOM_1677;
	logic [31:0] _RANDOM_1678;
	logic [31:0] _RANDOM_1679;
	logic [31:0] _RANDOM_1680;
	logic [31:0] _RANDOM_1681;
	logic [31:0] _RANDOM_1682;
	logic [31:0] _RANDOM_1683;
	logic [31:0] _RANDOM_1684;
	logic [31:0] _RANDOM_1685;
	logic [31:0] _RANDOM_1686;
	logic [31:0] _RANDOM_1687;
	logic [31:0] _RANDOM_1688;
	logic [31:0] _RANDOM_1689;
	logic [31:0] _RANDOM_1690;
	logic [31:0] _RANDOM_1691;
	logic [31:0] _RANDOM_1692;
	logic [31:0] _RANDOM_1693;
	logic [31:0] _RANDOM_1694;
	logic [31:0] _RANDOM_1695;
	logic [31:0] _RANDOM_1696;
	logic [31:0] _RANDOM_1697;
	logic [31:0] _RANDOM_1698;
	logic [31:0] _RANDOM_1699;
	logic [31:0] _RANDOM_1700;
	logic [31:0] _RANDOM_1701;
	logic [31:0] _RANDOM_1702;
	logic [31:0] _RANDOM_1703;
	logic [31:0] _RANDOM_1704;
	logic [31:0] _RANDOM_1705;
	logic [31:0] _RANDOM_1706;
	logic [31:0] _RANDOM_1707;
	logic [31:0] _RANDOM_1708;
	logic [31:0] _RANDOM_1709;
	logic [31:0] _RANDOM_1710;
	logic [31:0] _RANDOM_1711;
	logic [31:0] _RANDOM_1712;
	logic [31:0] _RANDOM_1713;
	logic [31:0] _RANDOM_1714;
	logic [31:0] _RANDOM_1715;
	logic [31:0] _RANDOM_1716;
	logic [31:0] _RANDOM_1717;
	logic [31:0] _RANDOM_1718;
	logic [31:0] _RANDOM_1719;
	logic [31:0] _RANDOM_1720;
	logic [31:0] _RANDOM_1721;
	logic [31:0] _RANDOM_1722;
	logic [31:0] _RANDOM_1723;
	logic [31:0] _RANDOM_1724;
	logic [31:0] _RANDOM_1725;
	logic [31:0] _RANDOM_1726;
	logic [31:0] _RANDOM_1727;
	logic [31:0] _RANDOM_1728;
	logic [31:0] _RANDOM_1729;
	logic [31:0] _RANDOM_1730;
	logic [31:0] _RANDOM_1731;
	logic [31:0] _RANDOM_1732;
	logic [31:0] _RANDOM_1733;
	logic [31:0] _RANDOM_1734;
	logic [31:0] _RANDOM_1735;
	logic [31:0] _RANDOM_1736;
	logic [31:0] _RANDOM_1737;
	logic [31:0] _RANDOM_1738;
	logic [31:0] _RANDOM_1739;
	logic [31:0] _RANDOM_1740;
	logic [31:0] _RANDOM_1741;
	logic [31:0] _RANDOM_1742;
	logic [31:0] _RANDOM_1743;
	logic [31:0] _RANDOM_1744;
	logic [31:0] _RANDOM_1745;
	logic [31:0] _RANDOM_1746;
	logic [31:0] _RANDOM_1747;
	logic [31:0] _RANDOM_1748;
	logic [31:0] _RANDOM_1749;
	logic [31:0] _RANDOM_1750;
	logic [31:0] _RANDOM_1751;
	logic [31:0] _RANDOM_1752;
	logic [31:0] _RANDOM_1753;
	logic [31:0] _RANDOM_1754;
	logic [31:0] _RANDOM_1755;
	logic [31:0] _RANDOM_1756;
	logic [31:0] _RANDOM_1757;
	logic [31:0] _RANDOM_1758;
	logic [31:0] _RANDOM_1759;
	logic [31:0] _RANDOM_1760;
	logic [31:0] _RANDOM_1761;
	logic [31:0] _RANDOM_1762;
	logic [31:0] _RANDOM_1763;
	logic [31:0] _RANDOM_1764;
	logic [31:0] _RANDOM_1765;
	logic [31:0] _RANDOM_1766;
	logic [31:0] _RANDOM_1767;
	logic [31:0] _RANDOM_1768;
	logic [31:0] _RANDOM_1769;
	logic [31:0] _RANDOM_1770;
	logic [31:0] _RANDOM_1771;
	logic [31:0] _RANDOM_1772;
	logic [31:0] _RANDOM_1773;
	logic [31:0] _RANDOM_1774;
	logic [31:0] _RANDOM_1775;
	logic [31:0] _RANDOM_1776;
	logic [31:0] _RANDOM_1777;
	logic [31:0] _RANDOM_1778;
	logic [31:0] _RANDOM_1779;
	logic [31:0] _RANDOM_1780;
	logic [31:0] _RANDOM_1781;
	logic [31:0] _RANDOM_1782;
	logic [31:0] _RANDOM_1783;
	logic [31:0] _RANDOM_1784;
	logic [31:0] _RANDOM_1785;
	logic [31:0] _RANDOM_1786;
	logic [31:0] _RANDOM_1787;
	logic [31:0] _RANDOM_1788;
	logic [31:0] _RANDOM_1789;
	logic [31:0] _RANDOM_1790;
	logic [31:0] _RANDOM_1791;
	logic [31:0] _RANDOM_1792;
	logic [31:0] _RANDOM_1793;
	logic [31:0] _RANDOM_1794;
	logic [31:0] _RANDOM_1795;
	logic [31:0] _RANDOM_1796;
	logic [31:0] _RANDOM_1797;
	logic [31:0] _RANDOM_1798;
	logic [31:0] _RANDOM_1799;
	logic [31:0] _RANDOM_1800;
	logic [31:0] _RANDOM_1801;
	logic [31:0] _RANDOM_1802;
	logic [31:0] _RANDOM_1803;
	logic [31:0] _RANDOM_1804;
	logic [31:0] _RANDOM_1805;
	logic [31:0] _RANDOM_1806;
	logic [31:0] _RANDOM_1807;
	logic [31:0] _RANDOM_1808;
	logic [31:0] _RANDOM_1809;
	logic [31:0] _RANDOM_1810;
	logic [31:0] _RANDOM_1811;
	logic [31:0] _RANDOM_1812;
	logic [31:0] _RANDOM_1813;
	logic [31:0] _RANDOM_1814;
	logic [31:0] _RANDOM_1815;
	logic [31:0] _RANDOM_1816;
	logic [31:0] _RANDOM_1817;
	logic [31:0] _RANDOM_1818;
	logic [31:0] _RANDOM_1819;
	logic [31:0] _RANDOM_1820;
	logic [31:0] _RANDOM_1821;
	logic [31:0] _RANDOM_1822;
	logic [31:0] _RANDOM_1823;
	logic [31:0] _RANDOM_1824;
	logic [31:0] _RANDOM_1825;
	logic [31:0] _RANDOM_1826;
	logic [31:0] _RANDOM_1827;
	logic [31:0] _RANDOM_1828;
	logic [31:0] _RANDOM_1829;
	logic [31:0] _RANDOM_1830;
	logic [31:0] _RANDOM_1831;
	logic [31:0] _RANDOM_1832;
	logic [31:0] _RANDOM_1833;
	logic [31:0] _RANDOM_1834;
	logic [31:0] _RANDOM_1835;
	logic [31:0] _RANDOM_1836;
	logic [31:0] _RANDOM_1837;
	logic [31:0] _RANDOM_1838;
	logic [31:0] _RANDOM_1839;
	logic [31:0] _RANDOM_1840;
	logic [31:0] _RANDOM_1841;
	logic [31:0] _RANDOM_1842;
	logic [31:0] _RANDOM_1843;
	logic [31:0] _RANDOM_1844;
	logic [31:0] _RANDOM_1845;
	logic [31:0] _RANDOM_1846;
	logic [31:0] _RANDOM_1847;
	logic [31:0] _RANDOM_1848;
	logic [31:0] _RANDOM_1849;
	logic [31:0] _RANDOM_1850;
	logic [31:0] _RANDOM_1851;
	logic [31:0] _RANDOM_1852;
	logic [31:0] _RANDOM_1853;
	logic [31:0] _RANDOM_1854;
	logic [31:0] _RANDOM_1855;
	logic [31:0] _RANDOM_1856;
	logic [31:0] _RANDOM_1857;
	logic [31:0] _RANDOM_1858;
	logic [31:0] _RANDOM_1859;
	logic [31:0] _RANDOM_1860;
	logic [31:0] _RANDOM_1861;
	logic [31:0] _RANDOM_1862;
	logic [31:0] _RANDOM_1863;
	logic [31:0] _RANDOM_1864;
	logic [31:0] _RANDOM_1865;
	logic [31:0] _RANDOM_1866;
	logic [31:0] _RANDOM_1867;
	logic [31:0] _RANDOM_1868;
	logic [31:0] _RANDOM_1869;
	logic [31:0] _RANDOM_1870;
	logic [31:0] _RANDOM_1871;
	logic [31:0] _RANDOM_1872;
	logic [31:0] _RANDOM_1873;
	logic [31:0] _RANDOM_1874;
	logic [31:0] _RANDOM_1875;
	logic [31:0] _RANDOM_1876;
	logic [31:0] _RANDOM_1877;
	logic [31:0] _RANDOM_1878;
	logic [31:0] _RANDOM_1879;
	logic [31:0] _RANDOM_1880;
	logic [31:0] _RANDOM_1881;
	logic [31:0] _RANDOM_1882;
	logic [31:0] _RANDOM_1883;
	logic [31:0] _RANDOM_1884;
	logic [31:0] _RANDOM_1885;
	logic [31:0] _RANDOM_1886;
	logic [31:0] _RANDOM_1887;
	logic [31:0] _RANDOM_1888;
	logic [31:0] _RANDOM_1889;
	logic [31:0] _RANDOM_1890;
	logic [31:0] _RANDOM_1891;
	logic [31:0] _RANDOM_1892;
	logic [31:0] _RANDOM_1893;
	logic [31:0] _RANDOM_1894;
	logic [31:0] _RANDOM_1895;
	logic [31:0] _RANDOM_1896;
	logic [31:0] _RANDOM_1897;
	logic [31:0] _RANDOM_1898;
	logic [31:0] _RANDOM_1899;
	logic [31:0] _RANDOM_1900;
	logic [31:0] _RANDOM_1901;
	logic [31:0] _RANDOM_1902;
	logic [31:0] _RANDOM_1903;
	logic [31:0] _RANDOM_1904;
	logic [31:0] _RANDOM_1905;
	logic [31:0] _RANDOM_1906;
	logic [31:0] _RANDOM_1907;
	logic [31:0] _RANDOM_1908;
	logic [31:0] _RANDOM_1909;
	logic [31:0] _RANDOM_1910;
	logic [31:0] _RANDOM_1911;
	logic [31:0] _RANDOM_1912;
	logic [31:0] _RANDOM_1913;
	logic [31:0] _RANDOM_1914;
	logic [31:0] _RANDOM_1915;
	logic [31:0] _RANDOM_1916;
	logic [31:0] _RANDOM_1917;
	logic [31:0] _RANDOM_1918;
	logic [31:0] _RANDOM_1919;
	logic [31:0] _RANDOM_1920;
	logic [31:0] _RANDOM_1921;
	logic [31:0] _RANDOM_1922;
	logic [31:0] _RANDOM_1923;
	logic [31:0] _RANDOM_1924;
	logic [31:0] _RANDOM_1925;
	logic [31:0] _RANDOM_1926;
	logic [31:0] _RANDOM_1927;
	logic [31:0] _RANDOM_1928;
	logic [31:0] _RANDOM_1929;
	logic [31:0] _RANDOM_1930;
	logic [31:0] _RANDOM_1931;
	logic [31:0] _RANDOM_1932;
	logic [31:0] _RANDOM_1933;
	logic [31:0] _RANDOM_1934;
	logic [31:0] _RANDOM_1935;
	logic [31:0] _RANDOM_1936;
	logic [31:0] _RANDOM_1937;
	logic [31:0] _RANDOM_1938;
	logic [31:0] _RANDOM_1939;
	logic [31:0] _RANDOM_1940;
	logic [31:0] _RANDOM_1941;
	logic [31:0] _RANDOM_1942;
	logic [31:0] _RANDOM_1943;
	logic [31:0] _RANDOM_1944;
	logic [31:0] _RANDOM_1945;
	logic [31:0] _RANDOM_1946;
	logic [31:0] _RANDOM_1947;
	logic [31:0] _RANDOM_1948;
	logic [31:0] _RANDOM_1949;
	logic [31:0] _RANDOM_1950;
	logic [31:0] _RANDOM_1951;
	logic [31:0] _RANDOM_1952;
	logic [31:0] _RANDOM_1953;
	logic [31:0] _RANDOM_1954;
	logic [31:0] _RANDOM_1955;
	logic [31:0] _RANDOM_1956;
	logic [31:0] _RANDOM_1957;
	logic [31:0] _RANDOM_1958;
	logic [31:0] _RANDOM_1959;
	logic [31:0] _RANDOM_1960;
	logic [31:0] _RANDOM_1961;
	logic [31:0] _RANDOM_1962;
	logic [31:0] _RANDOM_1963;
	logic [31:0] _RANDOM_1964;
	logic [31:0] _RANDOM_1965;
	logic [31:0] _RANDOM_1966;
	logic [31:0] _RANDOM_1967;
	logic [31:0] _RANDOM_1968;
	logic [31:0] _RANDOM_1969;
	logic [31:0] _RANDOM_1970;
	logic [31:0] _RANDOM_1971;
	logic [31:0] _RANDOM_1972;
	logic [31:0] _RANDOM_1973;
	logic [31:0] _RANDOM_1974;
	logic [31:0] _RANDOM_1975;
	logic [31:0] _RANDOM_1976;
	logic [31:0] _RANDOM_1977;
	logic [31:0] _RANDOM_1978;
	logic [31:0] _RANDOM_1979;
	logic [31:0] _RANDOM_1980;
	logic [31:0] _RANDOM_1981;
	logic [31:0] _RANDOM_1982;
	logic [31:0] _RANDOM_1983;
	logic [31:0] _RANDOM_1984;
	logic [31:0] _RANDOM_1985;
	logic [31:0] _RANDOM_1986;
	logic [31:0] _RANDOM_1987;
	logic [31:0] _RANDOM_1988;
	logic [31:0] _RANDOM_1989;
	logic [31:0] _RANDOM_1990;
	logic [31:0] _RANDOM_1991;
	logic [31:0] _RANDOM_1992;
	logic [31:0] _RANDOM_1993;
	logic [31:0] _RANDOM_1994;
	logic [31:0] _RANDOM_1995;
	logic [31:0] _RANDOM_1996;
	logic [31:0] _RANDOM_1997;
	logic [31:0] _RANDOM_1998;
	logic [31:0] _RANDOM_1999;
	logic [31:0] _RANDOM_2000;
	logic [31:0] _RANDOM_2001;
	logic [31:0] _RANDOM_2002;
	logic [31:0] _RANDOM_2003;
	logic [31:0] _RANDOM_2004;
	logic [31:0] _RANDOM_2005;
	logic [31:0] _RANDOM_2006;
	logic [31:0] _RANDOM_2007;
	logic [31:0] _RANDOM_2008;
	logic [31:0] _RANDOM_2009;
	logic [31:0] _RANDOM_2010;
	logic [31:0] _RANDOM_2011;
	logic [31:0] _RANDOM_2012;
	logic [31:0] _RANDOM_2013;
	logic [31:0] _RANDOM_2014;
	logic [31:0] _RANDOM_2015;
	logic [31:0] _RANDOM_2016;
	logic [31:0] _RANDOM_2017;
	logic [31:0] _RANDOM_2018;
	logic [31:0] _RANDOM_2019;
	logic [31:0] _RANDOM_2020;
	logic [31:0] _RANDOM_2021;
	logic [31:0] _RANDOM_2022;
	logic [31:0] _RANDOM_2023;
	logic [31:0] _RANDOM_2024;
	logic [31:0] _RANDOM_2025;
	logic [31:0] _RANDOM_2026;
	logic [31:0] _RANDOM_2027;
	logic [31:0] _RANDOM_2028;
	logic [31:0] _RANDOM_2029;
	logic [31:0] _RANDOM_2030;
	logic [31:0] _RANDOM_2031;
	logic [31:0] _RANDOM_2032;
	logic [31:0] _RANDOM_2033;
	logic [31:0] _RANDOM_2034;
	logic [31:0] _RANDOM_2035;
	logic [31:0] _RANDOM_2036;
	logic [31:0] _RANDOM_2037;
	logic [31:0] _RANDOM_2038;
	logic [31:0] _RANDOM_2039;
	logic [31:0] _RANDOM_2040;
	logic [31:0] _RANDOM_2041;
	logic [31:0] _RANDOM_2042;
	logic [31:0] _RANDOM_2043;
	logic [31:0] _RANDOM_2044;
	logic [31:0] _RANDOM_2045;
	logic [31:0] _RANDOM_2046;
	logic [31:0] _RANDOM_2047;
	logic [31:0] _RANDOM_2048;
	logic [31:0] _RANDOM_2049;
	logic [31:0] _RANDOM_2050;
	logic [31:0] _RANDOM_2051;
	logic [31:0] _RANDOM_2052;
	logic [31:0] _RANDOM_2053;
	logic [31:0] _RANDOM_2054;
	logic [31:0] _RANDOM_2055;
	logic [31:0] _RANDOM_2056;
	logic [31:0] _RANDOM_2057;
	logic [31:0] _RANDOM_2058;
	logic [31:0] _RANDOM_2059;
	logic [31:0] _RANDOM_2060;
	logic [31:0] _RANDOM_2061;
	logic [31:0] _RANDOM_2062;
	logic [31:0] _RANDOM_2063;
	logic [31:0] _RANDOM_2064;
	logic [31:0] _RANDOM_2065;
	logic [31:0] _RANDOM_2066;
	logic [31:0] _RANDOM_2067;
	logic [31:0] _RANDOM_2068;
	logic [31:0] _RANDOM_2069;
	logic [31:0] _RANDOM_2070;
	logic [31:0] _RANDOM_2071;
	logic [31:0] _RANDOM_2072;
	logic [31:0] _RANDOM_2073;
	logic [31:0] _RANDOM_2074;
	logic [31:0] _RANDOM_2075;
	logic [31:0] _RANDOM_2076;
	logic [31:0] _RANDOM_2077;
	logic [31:0] _RANDOM_2078;
	logic [31:0] _RANDOM_2079;
	logic [31:0] _RANDOM_2080;
	logic [31:0] _RANDOM_2081;
	logic [31:0] _RANDOM_2082;
	logic [31:0] _RANDOM_2083;
	logic [31:0] _RANDOM_2084;
	logic [31:0] _RANDOM_2085;
	logic [31:0] _RANDOM_2086;
	logic [31:0] _RANDOM_2087;
	logic [31:0] _RANDOM_2088;
	logic [31:0] _RANDOM_2089;
	logic [31:0] _RANDOM_2090;
	logic [31:0] _RANDOM_2091;
	logic [31:0] _RANDOM_2092;
	logic [31:0] _RANDOM_2093;
	logic [31:0] _RANDOM_2094;
	logic [31:0] _RANDOM_2095;
	logic [31:0] _RANDOM_2096;
	logic [31:0] _RANDOM_2097;
	logic [31:0] _RANDOM_2098;
	logic [31:0] _RANDOM_2099;
	logic [31:0] _RANDOM_2100;
	logic [31:0] _RANDOM_2101;
	logic [31:0] _RANDOM_2102;
	logic [31:0] _RANDOM_2103;
	logic [31:0] _RANDOM_2104;
	logic [31:0] _RANDOM_2105;
	logic [31:0] _RANDOM_2106;
	logic [31:0] _RANDOM_2107;
	logic [31:0] _RANDOM_2108;
	logic [31:0] _RANDOM_2109;
	logic [31:0] _RANDOM_2110;
	logic [31:0] _RANDOM_2111;
	logic [31:0] _RANDOM_2112;
	logic [31:0] _RANDOM_2113;
	logic [31:0] _RANDOM_2114;
	logic [31:0] _RANDOM_2115;
	logic [31:0] _RANDOM_2116;
	logic [31:0] _RANDOM_2117;
	logic [31:0] _RANDOM_2118;
	logic [31:0] _RANDOM_2119;
	logic [31:0] _RANDOM_2120;
	logic [31:0] _RANDOM_2121;
	logic [31:0] _RANDOM_2122;
	logic [31:0] _RANDOM_2123;
	logic [31:0] _RANDOM_2124;
	logic [31:0] _RANDOM_2125;
	logic [31:0] _RANDOM_2126;
	logic [31:0] _RANDOM_2127;
	logic [31:0] _RANDOM_2128;
	logic [31:0] _RANDOM_2129;
	logic [31:0] _RANDOM_2130;
	logic [31:0] _RANDOM_2131;
	logic [31:0] _RANDOM_2132;
	logic [31:0] _RANDOM_2133;
	logic [31:0] _RANDOM_2134;
	logic [31:0] _RANDOM_2135;
	logic [31:0] _RANDOM_2136;
	logic [31:0] _RANDOM_2137;
	logic [31:0] _RANDOM_2138;
	logic [31:0] _RANDOM_2139;
	logic [31:0] _RANDOM_2140;
	logic [31:0] _RANDOM_2141;
	logic [31:0] _RANDOM_2142;
	logic [31:0] _RANDOM_2143;
	logic [31:0] _RANDOM_2144;
	logic [31:0] _RANDOM_2145;
	logic [31:0] _RANDOM_2146;
	logic [31:0] _RANDOM_2147;
	logic [31:0] _RANDOM_2148;
	logic [31:0] _RANDOM_2149;
	logic [31:0] _RANDOM_2150;
	logic [31:0] _RANDOM_2151;
	logic [31:0] _RANDOM_2152;
	logic [31:0] _RANDOM_2153;
	logic [31:0] _RANDOM_2154;
	logic [31:0] _RANDOM_2155;
	logic [31:0] _RANDOM_2156;
	logic [31:0] _RANDOM_2157;
	logic [31:0] _RANDOM_2158;
	logic [31:0] _RANDOM_2159;
	logic [31:0] _RANDOM_2160;
	logic [31:0] _RANDOM_2161;
	logic [31:0] _RANDOM_2162;
	logic [31:0] _RANDOM_2163;
	logic [31:0] _RANDOM_2164;
	logic [31:0] _RANDOM_2165;
	logic [31:0] _RANDOM_2166;
	logic [31:0] _RANDOM_2167;
	logic [31:0] _RANDOM_2168;
	logic [31:0] _RANDOM_2169;
	logic [31:0] _RANDOM_2170;
	logic [31:0] _RANDOM_2171;
	logic [31:0] _RANDOM_2172;
	logic [31:0] _RANDOM_2173;
	logic [31:0] _RANDOM_2174;
	logic [31:0] _RANDOM_2175;
	logic [31:0] _RANDOM_2176;
	logic [31:0] _RANDOM_2177;
	logic [31:0] _RANDOM_2178;
	logic [31:0] _RANDOM_2179;
	logic [31:0] _RANDOM_2180;
	logic [31:0] _RANDOM_2181;
	logic [31:0] _RANDOM_2182;
	logic [31:0] _RANDOM_2183;
	logic [31:0] _RANDOM_2184;
	logic [31:0] _RANDOM_2185;
	logic [31:0] _RANDOM_2186;
	logic [31:0] _RANDOM_2187;
	logic [31:0] _RANDOM_2188;
	logic [31:0] _RANDOM_2189;
	logic [31:0] _RANDOM_2190;
	logic [31:0] _RANDOM_2191;
	logic [31:0] _RANDOM_2192;
	logic [31:0] _RANDOM_2193;
	logic [31:0] _RANDOM_2194;
	logic [31:0] _RANDOM_2195;
	logic [31:0] _RANDOM_2196;
	logic [31:0] _RANDOM_2197;
	logic [31:0] _RANDOM_2198;
	logic [31:0] _RANDOM_2199;
	logic [31:0] _RANDOM_2200;
	logic [31:0] _RANDOM_2201;
	logic [31:0] _RANDOM_2202;
	logic [31:0] _RANDOM_2203;
	logic [31:0] _RANDOM_2204;
	logic [31:0] _RANDOM_2205;
	logic [31:0] _RANDOM_2206;
	logic [31:0] _RANDOM_2207;
	logic [31:0] _RANDOM_2208;
	logic [31:0] _RANDOM_2209;
	logic [31:0] _RANDOM_2210;
	logic [31:0] _RANDOM_2211;
	logic [31:0] _RANDOM_2212;
	logic [31:0] _RANDOM_2213;
	logic [31:0] _RANDOM_2214;
	logic [31:0] _RANDOM_2215;
	logic [31:0] _RANDOM_2216;
	logic [31:0] _RANDOM_2217;
	logic [31:0] _RANDOM_2218;
	logic [31:0] _RANDOM_2219;
	logic [31:0] _RANDOM_2220;
	logic [31:0] _RANDOM_2221;
	logic [31:0] _RANDOM_2222;
	logic [31:0] _RANDOM_2223;
	logic [31:0] _RANDOM_2224;
	logic [31:0] _RANDOM_2225;
	logic [31:0] _RANDOM_2226;
	logic [31:0] _RANDOM_2227;
	logic [31:0] _RANDOM_2228;
	logic [31:0] _RANDOM_2229;
	logic [31:0] _RANDOM_2230;
	logic [31:0] _RANDOM_2231;
	logic [31:0] _RANDOM_2232;
	logic [31:0] _RANDOM_2233;
	logic [31:0] _RANDOM_2234;
	logic [31:0] _RANDOM_2235;
	logic [31:0] _RANDOM_2236;
	logic [31:0] _RANDOM_2237;
	logic [31:0] _RANDOM_2238;
	logic [31:0] _RANDOM_2239;
	logic [31:0] _RANDOM_2240;
	logic [31:0] _RANDOM_2241;
	logic [31:0] _RANDOM_2242;
	logic [31:0] _RANDOM_2243;
	logic [31:0] _RANDOM_2244;
	logic [31:0] _RANDOM_2245;
	logic [31:0] _RANDOM_2246;
	logic [31:0] _RANDOM_2247;
	logic [31:0] _RANDOM_2248;
	logic [31:0] _RANDOM_2249;
	logic [31:0] _RANDOM_2250;
	logic [31:0] _RANDOM_2251;
	logic [31:0] _RANDOM_2252;
	logic [31:0] _RANDOM_2253;
	logic [31:0] _RANDOM_2254;
	logic [31:0] _RANDOM_2255;
	logic [31:0] _RANDOM_2256;
	logic [31:0] _RANDOM_2257;
	logic [31:0] _RANDOM_2258;
	logic [31:0] _RANDOM_2259;
	logic [31:0] _RANDOM_2260;
	logic [31:0] _RANDOM_2261;
	logic [31:0] _RANDOM_2262;
	logic [31:0] _RANDOM_2263;
	logic [31:0] _RANDOM_2264;
	logic [31:0] _RANDOM_2265;
	logic [31:0] _RANDOM_2266;
	logic [31:0] _RANDOM_2267;
	logic [31:0] _RANDOM_2268;
	logic [31:0] _RANDOM_2269;
	logic [31:0] _RANDOM_2270;
	logic [31:0] _RANDOM_2271;
	logic [31:0] _RANDOM_2272;
	logic [31:0] _RANDOM_2273;
	logic [31:0] _RANDOM_2274;
	logic [31:0] _RANDOM_2275;
	logic [31:0] _RANDOM_2276;
	logic [31:0] _RANDOM_2277;
	logic [31:0] _RANDOM_2278;
	logic [31:0] _RANDOM_2279;
	logic [31:0] _RANDOM_2280;
	logic [31:0] _RANDOM_2281;
	logic [31:0] _RANDOM_2282;
	logic [31:0] _RANDOM_2283;
	logic [31:0] _RANDOM_2284;
	logic [31:0] _RANDOM_2285;
	logic [31:0] _RANDOM_2286;
	logic [31:0] _RANDOM_2287;
	logic [31:0] _RANDOM_2288;
	logic [31:0] _RANDOM_2289;
	logic [31:0] _RANDOM_2290;
	logic [31:0] _RANDOM_2291;
	logic [31:0] _RANDOM_2292;
	logic [31:0] _RANDOM_2293;
	logic [31:0] _RANDOM_2294;
	logic [31:0] _RANDOM_2295;
	logic [31:0] _RANDOM_2296;
	logic [31:0] _RANDOM_2297;
	logic [31:0] _RANDOM_2298;
	logic [31:0] _RANDOM_2299;
	logic [31:0] _RANDOM_2300;
	logic [31:0] _RANDOM_2301;
	logic [31:0] _RANDOM_2302;
	logic [31:0] _RANDOM_2303;
	logic [31:0] _RANDOM_2304;
	logic [31:0] _RANDOM_2305;
	logic [31:0] _RANDOM_2306;
	logic [31:0] _RANDOM_2307;
	logic [31:0] _RANDOM_2308;
	logic [31:0] _RANDOM_2309;
	logic [31:0] _RANDOM_2310;
	logic [31:0] _RANDOM_2311;
	logic [31:0] _RANDOM_2312;
	logic [31:0] _RANDOM_2313;
	logic [31:0] _RANDOM_2314;
	logic [31:0] _RANDOM_2315;
	logic [31:0] _RANDOM_2316;
	logic [31:0] _RANDOM_2317;
	logic [31:0] _RANDOM_2318;
	logic [31:0] _RANDOM_2319;
	logic [31:0] _RANDOM_2320;
	logic [31:0] _RANDOM_2321;
	logic [31:0] _RANDOM_2322;
	logic [31:0] _RANDOM_2323;
	logic [31:0] _RANDOM_2324;
	logic [31:0] _RANDOM_2325;
	logic [31:0] _RANDOM_2326;
	logic [31:0] _RANDOM_2327;
	logic [31:0] _RANDOM_2328;
	logic [31:0] _RANDOM_2329;
	logic [31:0] _RANDOM_2330;
	logic [31:0] _RANDOM_2331;
	logic [31:0] _RANDOM_2332;
	logic [31:0] _RANDOM_2333;
	logic [31:0] _RANDOM_2334;
	logic [31:0] _RANDOM_2335;
	logic [31:0] _RANDOM_2336;
	logic [31:0] _RANDOM_2337;
	logic [31:0] _RANDOM_2338;
	logic [31:0] _RANDOM_2339;
	logic [31:0] _RANDOM_2340;
	logic [31:0] _RANDOM_2341;
	logic [31:0] _RANDOM_2342;
	logic [31:0] _RANDOM_2343;
	logic [31:0] _RANDOM_2344;
	logic [31:0] _RANDOM_2345;
	logic [31:0] _RANDOM_2346;
	logic [31:0] _RANDOM_2347;
	logic [31:0] _RANDOM_2348;
	logic [31:0] _RANDOM_2349;
	logic [31:0] _RANDOM_2350;
	logic [31:0] _RANDOM_2351;
	logic [31:0] _RANDOM_2352;
	logic [31:0] _RANDOM_2353;
	logic [31:0] _RANDOM_2354;
	logic [31:0] _RANDOM_2355;
	logic [31:0] _RANDOM_2356;
	logic [31:0] _RANDOM_2357;
	logic [31:0] _RANDOM_2358;
	logic [31:0] _RANDOM_2359;
	logic [31:0] _RANDOM_2360;
	logic [31:0] _RANDOM_2361;
	logic [31:0] _RANDOM_2362;
	logic [31:0] _RANDOM_2363;
	logic [31:0] _RANDOM_2364;
	logic [31:0] _RANDOM_2365;
	logic [31:0] _RANDOM_2366;
	logic [31:0] _RANDOM_2367;
	logic [31:0] _RANDOM_2368;
	logic [31:0] _RANDOM_2369;
	logic [31:0] _RANDOM_2370;
	logic [31:0] _RANDOM_2371;
	logic [31:0] _RANDOM_2372;
	logic [31:0] _RANDOM_2373;
	logic [31:0] _RANDOM_2374;
	logic [31:0] _RANDOM_2375;
	logic [31:0] _RANDOM_2376;
	logic [31:0] _RANDOM_2377;
	logic [31:0] _RANDOM_2378;
	logic [31:0] _RANDOM_2379;
	logic [31:0] _RANDOM_2380;
	logic [31:0] _RANDOM_2381;
	logic [31:0] _RANDOM_2382;
	logic [31:0] _RANDOM_2383;
	logic [31:0] _RANDOM_2384;
	logic [31:0] _RANDOM_2385;
	logic [31:0] _RANDOM_2386;
	logic [31:0] _RANDOM_2387;
	logic [31:0] _RANDOM_2388;
	logic [31:0] _RANDOM_2389;
	logic [31:0] _RANDOM_2390;
	logic [31:0] _RANDOM_2391;
	logic [31:0] _RANDOM_2392;
	logic [31:0] _RANDOM_2393;
	logic [31:0] _RANDOM_2394;
	logic [31:0] _RANDOM_2395;
	logic [31:0] _RANDOM_2396;
	logic [31:0] _RANDOM_2397;
	logic [31:0] _RANDOM_2398;
	logic [31:0] _RANDOM_2399;
	logic [31:0] _RANDOM_2400;
	logic [31:0] _RANDOM_2401;
	logic [31:0] _RANDOM_2402;
	logic [31:0] _RANDOM_2403;
	logic [31:0] _RANDOM_2404;
	logic [31:0] _RANDOM_2405;
	logic [31:0] _RANDOM_2406;
	logic [31:0] _RANDOM_2407;
	logic [31:0] _RANDOM_2408;
	logic [31:0] _RANDOM_2409;
	logic [31:0] _RANDOM_2410;
	logic [31:0] _RANDOM_2411;
	logic [31:0] _RANDOM_2412;
	logic [31:0] _RANDOM_2413;
	logic [31:0] _RANDOM_2414;
	logic [31:0] _RANDOM_2415;
	logic [31:0] _RANDOM_2416;
	logic [31:0] _RANDOM_2417;
	logic [31:0] _RANDOM_2418;
	logic [31:0] _RANDOM_2419;
	logic [31:0] _RANDOM_2420;
	logic [31:0] _RANDOM_2421;
	logic [31:0] _RANDOM_2422;
	logic [31:0] _RANDOM_2423;
	logic [31:0] _RANDOM_2424;
	logic [31:0] _RANDOM_2425;
	logic [31:0] _RANDOM_2426;
	logic [31:0] _RANDOM_2427;
	logic [31:0] _RANDOM_2428;
	logic [31:0] _RANDOM_2429;
	logic [31:0] _RANDOM_2430;
	logic [31:0] _RANDOM_2431;
	logic [31:0] _RANDOM_2432;
	logic [31:0] _RANDOM_2433;
	logic [31:0] _RANDOM_2434;
	logic [31:0] _RANDOM_2435;
	logic [31:0] _RANDOM_2436;
	logic [31:0] _RANDOM_2437;
	logic [31:0] _RANDOM_2438;
	logic [31:0] _RANDOM_2439;
	logic [31:0] _RANDOM_2440;
	logic [31:0] _RANDOM_2441;
	logic [31:0] _RANDOM_2442;
	logic [31:0] _RANDOM_2443;
	logic [31:0] _RANDOM_2444;
	logic [31:0] _RANDOM_2445;
	logic [31:0] _RANDOM_2446;
	logic [31:0] _RANDOM_2447;
	logic [31:0] _RANDOM_2448;
	logic [31:0] _RANDOM_2449;
	logic [31:0] _RANDOM_2450;
	logic [31:0] _RANDOM_2451;
	logic [31:0] _RANDOM_2452;
	logic [31:0] _RANDOM_2453;
	logic [31:0] _RANDOM_2454;
	logic [31:0] _RANDOM_2455;
	logic [31:0] _RANDOM_2456;
	logic [31:0] _RANDOM_2457;
	logic [31:0] _RANDOM_2458;
	logic [31:0] _RANDOM_2459;
	logic [31:0] _RANDOM_2460;
	logic [31:0] _RANDOM_2461;
	logic [31:0] _RANDOM_2462;
	logic [31:0] _RANDOM_2463;
	logic [31:0] _RANDOM_2464;
	logic [31:0] _RANDOM_2465;
	logic [31:0] _RANDOM_2466;
	logic [31:0] _RANDOM_2467;
	logic [31:0] _RANDOM_2468;
	logic [31:0] _RANDOM_2469;
	logic [31:0] _RANDOM_2470;
	logic [31:0] _RANDOM_2471;
	logic [31:0] _RANDOM_2472;
	logic [31:0] _RANDOM_2473;
	logic [31:0] _RANDOM_2474;
	logic [31:0] _RANDOM_2475;
	logic [31:0] _RANDOM_2476;
	logic [31:0] _RANDOM_2477;
	logic [31:0] _RANDOM_2478;
	logic [31:0] _RANDOM_2479;
	logic [31:0] _RANDOM_2480;
	logic [31:0] _RANDOM_2481;
	logic [31:0] _RANDOM_2482;
	logic [31:0] _RANDOM_2483;
	logic [31:0] _RANDOM_2484;
	logic [31:0] _RANDOM_2485;
	logic [31:0] _RANDOM_2486;
	logic [31:0] _RANDOM_2487;
	logic [31:0] _RANDOM_2488;
	logic [31:0] _RANDOM_2489;
	logic [31:0] _RANDOM_2490;
	logic [31:0] _RANDOM_2491;
	logic [31:0] _RANDOM_2492;
	logic [31:0] _RANDOM_2493;
	logic [31:0] _RANDOM_2494;
	logic [31:0] _RANDOM_2495;
	logic [31:0] _RANDOM_2496;
	logic [31:0] _RANDOM_2497;
	logic [31:0] _RANDOM_2498;
	logic [31:0] _RANDOM_2499;
	logic [31:0] _RANDOM_2500;
	logic [31:0] _RANDOM_2501;
	logic [31:0] _RANDOM_2502;
	logic [31:0] _RANDOM_2503;
	logic [31:0] _RANDOM_2504;
	logic [31:0] _RANDOM_2505;
	logic [31:0] _RANDOM_2506;
	logic [31:0] _RANDOM_2507;
	logic [31:0] _RANDOM_2508;
	logic [31:0] _RANDOM_2509;
	logic [31:0] _RANDOM_2510;
	logic [31:0] _RANDOM_2511;
	logic [31:0] _RANDOM_2512;
	logic [31:0] _RANDOM_2513;
	logic [31:0] _RANDOM_2514;
	logic [31:0] _RANDOM_2515;
	logic [31:0] _RANDOM_2516;
	logic [31:0] _RANDOM_2517;
	logic [31:0] _RANDOM_2518;
	logic [31:0] _RANDOM_2519;
	logic [31:0] _RANDOM_2520;
	logic [31:0] _RANDOM_2521;
	logic [31:0] _RANDOM_2522;
	logic [31:0] _RANDOM_2523;
	logic [31:0] _RANDOM_2524;
	logic [31:0] _RANDOM_2525;
	logic [31:0] _RANDOM_2526;
	logic [31:0] _RANDOM_2527;
	logic [31:0] _RANDOM_2528;
	logic [31:0] _RANDOM_2529;
	logic [31:0] _RANDOM_2530;
	logic [31:0] _RANDOM_2531;
	logic [31:0] _RANDOM_2532;
	logic [31:0] _RANDOM_2533;
	logic [31:0] _RANDOM_2534;
	logic [31:0] _RANDOM_2535;
	logic [31:0] _RANDOM_2536;
	logic [31:0] _RANDOM_2537;
	logic [31:0] _RANDOM_2538;
	logic [31:0] _RANDOM_2539;
	logic [31:0] _RANDOM_2540;
	logic [31:0] _RANDOM_2541;
	logic [31:0] _RANDOM_2542;
	logic [31:0] _RANDOM_2543;
	logic [31:0] _RANDOM_2544;
	logic [31:0] _RANDOM_2545;
	logic [31:0] _RANDOM_2546;
	logic [31:0] _RANDOM_2547;
	logic [31:0] _RANDOM_2548;
	logic [31:0] _RANDOM_2549;
	logic [31:0] _RANDOM_2550;
	logic [31:0] _RANDOM_2551;
	logic [31:0] _RANDOM_2552;
	logic [31:0] _RANDOM_2553;
	logic [31:0] _RANDOM_2554;
	logic [31:0] _RANDOM_2555;
	logic [31:0] _RANDOM_2556;
	logic [31:0] _RANDOM_2557;
	logic [31:0] _RANDOM_2558;
	logic [31:0] _RANDOM_2559;
	logic [31:0] _RANDOM_2560;
	logic [31:0] _RANDOM_2561;
	logic [31:0] _RANDOM_2562;
	logic [31:0] _RANDOM_2563;
	logic [31:0] _RANDOM_2564;
	logic [31:0] _RANDOM_2565;
	logic [31:0] _RANDOM_2566;
	logic [31:0] _RANDOM_2567;
	logic [31:0] _RANDOM_2568;
	logic [31:0] _RANDOM_2569;
	logic [31:0] _RANDOM_2570;
	logic [31:0] _RANDOM_2571;
	logic [31:0] _RANDOM_2572;
	logic [31:0] _RANDOM_2573;
	logic [31:0] _RANDOM_2574;
	logic [31:0] _RANDOM_2575;
	logic [31:0] _RANDOM_2576;
	logic [31:0] _RANDOM_2577;
	logic [31:0] _RANDOM_2578;
	logic [31:0] _RANDOM_2579;
	logic [31:0] _RANDOM_2580;
	logic [31:0] _RANDOM_2581;
	logic [31:0] _RANDOM_2582;
	logic [31:0] _RANDOM_2583;
	logic [31:0] _RANDOM_2584;
	logic [31:0] _RANDOM_2585;
	logic [31:0] _RANDOM_2586;
	logic [31:0] _RANDOM_2587;
	logic [31:0] _RANDOM_2588;
	logic [31:0] _RANDOM_2589;
	logic [31:0] _RANDOM_2590;
	logic [31:0] _RANDOM_2591;
	logic [31:0] _RANDOM_2592;
	logic [31:0] _RANDOM_2593;
	logic [31:0] _RANDOM_2594;
	logic [31:0] _RANDOM_2595;
	logic [31:0] _RANDOM_2596;
	logic [31:0] _RANDOM_2597;
	logic [31:0] _RANDOM_2598;
	logic [31:0] _RANDOM_2599;
	logic [31:0] _RANDOM_2600;
	logic [31:0] _RANDOM_2601;
	logic [31:0] _RANDOM_2602;
	logic [31:0] _RANDOM_2603;
	logic [31:0] _RANDOM_2604;
	logic [31:0] _RANDOM_2605;
	logic [31:0] _RANDOM_2606;
	logic [31:0] _RANDOM_2607;
	logic [31:0] _RANDOM_2608;
	logic [31:0] _RANDOM_2609;
	logic [31:0] _RANDOM_2610;
	logic [31:0] _RANDOM_2611;
	logic [31:0] _RANDOM_2612;
	logic [31:0] _RANDOM_2613;
	logic [31:0] _RANDOM_2614;
	logic [31:0] _RANDOM_2615;
	logic [31:0] _RANDOM_2616;
	logic [31:0] _RANDOM_2617;
	logic [31:0] _RANDOM_2618;
	logic [31:0] _RANDOM_2619;
	logic [31:0] _RANDOM_2620;
	logic [31:0] _RANDOM_2621;
	logic [31:0] _RANDOM_2622;
	logic [31:0] _RANDOM_2623;
	logic [31:0] _RANDOM_2624;
	logic [31:0] _RANDOM_2625;
	logic [31:0] _RANDOM_2626;
	logic [31:0] _RANDOM_2627;
	logic [31:0] _RANDOM_2628;
	logic [31:0] _RANDOM_2629;
	logic [31:0] _RANDOM_2630;
	logic [31:0] _RANDOM_2631;
	logic [31:0] _RANDOM_2632;
	logic [31:0] _RANDOM_2633;
	logic [31:0] _RANDOM_2634;
	logic [31:0] _RANDOM_2635;
	logic [31:0] _RANDOM_2636;
	logic [31:0] _RANDOM_2637;
	logic [31:0] _RANDOM_2638;
	logic [31:0] _RANDOM_2639;
	logic [31:0] _RANDOM_2640;
	logic [31:0] _RANDOM_2641;
	logic [31:0] _RANDOM_2642;
	logic [31:0] _RANDOM_2643;
	logic [31:0] _RANDOM_2644;
	logic [31:0] _RANDOM_2645;
	logic [31:0] _RANDOM_2646;
	logic [31:0] _RANDOM_2647;
	logic [31:0] _RANDOM_2648;
	logic [31:0] _RANDOM_2649;
	logic [31:0] _RANDOM_2650;
	logic [31:0] _RANDOM_2651;
	logic [31:0] _RANDOM_2652;
	logic [31:0] _RANDOM_2653;
	logic [31:0] _RANDOM_2654;
	logic [31:0] _RANDOM_2655;
	logic [31:0] _RANDOM_2656;
	logic [31:0] _RANDOM_2657;
	logic [31:0] _RANDOM_2658;
	logic [31:0] _RANDOM_2659;
	logic [31:0] _RANDOM_2660;
	logic [31:0] _RANDOM_2661;
	logic [31:0] _RANDOM_2662;
	logic [31:0] _RANDOM_2663;
	logic [31:0] _RANDOM_2664;
	logic [31:0] _RANDOM_2665;
	logic [31:0] _RANDOM_2666;
	logic [31:0] _RANDOM_2667;
	logic [31:0] _RANDOM_2668;
	logic [31:0] _RANDOM_2669;
	logic [31:0] _RANDOM_2670;
	logic [31:0] _RANDOM_2671;
	logic [31:0] _RANDOM_2672;
	logic [31:0] _RANDOM_2673;
	logic [31:0] _RANDOM_2674;
	logic [31:0] _RANDOM_2675;
	logic [31:0] _RANDOM_2676;
	logic [31:0] _RANDOM_2677;
	logic [31:0] _RANDOM_2678;
	logic [31:0] _RANDOM_2679;
	logic [31:0] _RANDOM_2680;
	logic [31:0] _RANDOM_2681;
	logic [31:0] _RANDOM_2682;
	logic [31:0] _RANDOM_2683;
	logic [31:0] _RANDOM_2684;
	logic [31:0] _RANDOM_2685;
	logic [31:0] _RANDOM_2686;
	logic [31:0] _RANDOM_2687;
	logic [31:0] _RANDOM_2688;
	logic [31:0] _RANDOM_2689;
	logic [31:0] _RANDOM_2690;
	logic [31:0] _RANDOM_2691;
	logic [31:0] _RANDOM_2692;
	logic [31:0] _RANDOM_2693;
	logic [31:0] _RANDOM_2694;
	logic [31:0] _RANDOM_2695;
	logic [31:0] _RANDOM_2696;
	logic [31:0] _RANDOM_2697;
	logic [31:0] _RANDOM_2698;
	logic [31:0] _RANDOM_2699;
	logic [31:0] _RANDOM_2700;
	logic [31:0] _RANDOM_2701;
	logic [31:0] _RANDOM_2702;
	logic [31:0] _RANDOM_2703;
	logic [31:0] _RANDOM_2704;
	logic [31:0] _RANDOM_2705;
	logic [31:0] _RANDOM_2706;
	logic [31:0] _RANDOM_2707;
	logic [31:0] _RANDOM_2708;
	logic [31:0] _RANDOM_2709;
	logic [31:0] _RANDOM_2710;
	logic [31:0] _RANDOM_2711;
	logic [31:0] _RANDOM_2712;
	logic [31:0] _RANDOM_2713;
	logic [31:0] _RANDOM_2714;
	logic [31:0] _RANDOM_2715;
	logic [31:0] _RANDOM_2716;
	logic [31:0] _RANDOM_2717;
	logic [31:0] _RANDOM_2718;
	logic [31:0] _RANDOM_2719;
	logic [31:0] _RANDOM_2720;
	logic [31:0] _RANDOM_2721;
	logic [31:0] _RANDOM_2722;
	logic [31:0] _RANDOM_2723;
	logic [31:0] _RANDOM_2724;
	logic [31:0] _RANDOM_2725;
	logic [31:0] _RANDOM_2726;
	logic [31:0] _RANDOM_2727;
	logic [31:0] _RANDOM_2728;
	logic [31:0] _RANDOM_2729;
	logic [31:0] _RANDOM_2730;
	logic [31:0] _RANDOM_2731;
	logic [31:0] _RANDOM_2732;
	logic [31:0] _RANDOM_2733;
	logic [31:0] _RANDOM_2734;
	logic [31:0] _RANDOM_2735;
	logic [31:0] _RANDOM_2736;
	logic [31:0] _RANDOM_2737;
	logic [31:0] _RANDOM_2738;
	logic [31:0] _RANDOM_2739;
	logic [31:0] _RANDOM_2740;
	logic [31:0] _RANDOM_2741;
	logic [31:0] _RANDOM_2742;
	logic [31:0] _RANDOM_2743;
	logic [31:0] _RANDOM_2744;
	logic [31:0] _RANDOM_2745;
	logic [31:0] _RANDOM_2746;
	logic [31:0] _RANDOM_2747;
	logic [31:0] _RANDOM_2748;
	logic [31:0] _RANDOM_2749;
	logic [31:0] _RANDOM_2750;
	logic [31:0] _RANDOM_2751;
	logic [31:0] _RANDOM_2752;
	logic [31:0] _RANDOM_2753;
	logic [31:0] _RANDOM_2754;
	logic [31:0] _RANDOM_2755;
	logic [31:0] _RANDOM_2756;
	logic [31:0] _RANDOM_2757;
	logic [31:0] _RANDOM_2758;
	logic [31:0] _RANDOM_2759;
	logic [31:0] _RANDOM_2760;
	logic [31:0] _RANDOM_2761;
	logic [31:0] _RANDOM_2762;
	logic [31:0] _RANDOM_2763;
	logic [31:0] _RANDOM_2764;
	logic [31:0] _RANDOM_2765;
	logic [31:0] _RANDOM_2766;
	logic [31:0] _RANDOM_2767;
	logic [31:0] _RANDOM_2768;
	logic [31:0] _RANDOM_2769;
	logic [31:0] _RANDOM_2770;
	logic [31:0] _RANDOM_2771;
	logic [31:0] _RANDOM_2772;
	logic [31:0] _RANDOM_2773;
	logic [31:0] _RANDOM_2774;
	logic [31:0] _RANDOM_2775;
	logic [31:0] _RANDOM_2776;
	logic [31:0] _RANDOM_2777;
	logic [31:0] _RANDOM_2778;
	logic [31:0] _RANDOM_2779;
	logic [31:0] _RANDOM_2780;
	logic [31:0] _RANDOM_2781;
	logic [31:0] _RANDOM_2782;
	logic [31:0] _RANDOM_2783;
	logic [31:0] _RANDOM_2784;
	logic [31:0] _RANDOM_2785;
	logic [31:0] _RANDOM_2786;
	logic [31:0] _RANDOM_2787;
	logic [31:0] _RANDOM_2788;
	logic [31:0] _RANDOM_2789;
	logic [31:0] _RANDOM_2790;
	logic [31:0] _RANDOM_2791;
	logic [31:0] _RANDOM_2792;
	logic [31:0] _RANDOM_2793;
	logic [31:0] _RANDOM_2794;
	logic [31:0] _RANDOM_2795;
	logic [31:0] _RANDOM_2796;
	logic [31:0] _RANDOM_2797;
	logic [31:0] _RANDOM_2798;
	logic [31:0] _RANDOM_2799;
	logic [31:0] _RANDOM_2800;
	logic [31:0] _RANDOM_2801;
	logic [31:0] _RANDOM_2802;
	logic [31:0] _RANDOM_2803;
	logic [31:0] _RANDOM_2804;
	logic [31:0] _RANDOM_2805;
	logic [31:0] _RANDOM_2806;
	logic [31:0] _RANDOM_2807;
	logic [31:0] _RANDOM_2808;
	logic [31:0] _RANDOM_2809;
	logic [31:0] _RANDOM_2810;
	logic [31:0] _RANDOM_2811;
	logic [31:0] _RANDOM_2812;
	logic [31:0] _RANDOM_2813;
	logic [31:0] _RANDOM_2814;
	logic [31:0] _RANDOM_2815;
	logic [31:0] _RANDOM_2816;
	logic [31:0] _RANDOM_2817;
	logic [31:0] _RANDOM_2818;
	logic [31:0] _RANDOM_2819;
	logic [31:0] _RANDOM_2820;
	logic [31:0] _RANDOM_2821;
	logic [31:0] _RANDOM_2822;
	logic [31:0] _RANDOM_2823;
	logic [31:0] _RANDOM_2824;
	logic [31:0] _RANDOM_2825;
	logic [31:0] _RANDOM_2826;
	logic [31:0] _RANDOM_2827;
	logic [31:0] _RANDOM_2828;
	logic [31:0] _RANDOM_2829;
	logic [31:0] _RANDOM_2830;
	logic [31:0] _RANDOM_2831;
	logic [31:0] _RANDOM_2832;
	logic [31:0] _RANDOM_2833;
	logic [31:0] _RANDOM_2834;
	logic [31:0] _RANDOM_2835;
	logic [31:0] _RANDOM_2836;
	logic [31:0] _RANDOM_2837;
	logic [31:0] _RANDOM_2838;
	logic [31:0] _RANDOM_2839;
	logic [31:0] _RANDOM_2840;
	logic [31:0] _RANDOM_2841;
	logic [31:0] _RANDOM_2842;
	logic [31:0] _RANDOM_2843;
	logic [31:0] _RANDOM_2844;
	logic [31:0] _RANDOM_2845;
	logic [31:0] _RANDOM_2846;
	logic [31:0] _RANDOM_2847;
	logic [31:0] _RANDOM_2848;
	logic [31:0] _RANDOM_2849;
	logic [31:0] _RANDOM_2850;
	logic [31:0] _RANDOM_2851;
	logic [31:0] _RANDOM_2852;
	logic [31:0] _RANDOM_2853;
	logic [31:0] _RANDOM_2854;
	logic [31:0] _RANDOM_2855;
	logic [31:0] _RANDOM_2856;
	logic [31:0] _RANDOM_2857;
	logic [31:0] _RANDOM_2858;
	logic [31:0] _RANDOM_2859;
	logic [31:0] _RANDOM_2860;
	logic [31:0] _RANDOM_2861;
	logic [31:0] _RANDOM_2862;
	logic [31:0] _RANDOM_2863;
	logic [31:0] _RANDOM_2864;
	logic [31:0] _RANDOM_2865;
	logic [31:0] _RANDOM_2866;
	logic [31:0] _RANDOM_2867;
	logic [31:0] _RANDOM_2868;
	logic [31:0] _RANDOM_2869;
	logic [31:0] _RANDOM_2870;
	logic [31:0] _RANDOM_2871;
	logic [31:0] _RANDOM_2872;
	logic [31:0] _RANDOM_2873;
	logic [31:0] _RANDOM_2874;
	logic [31:0] _RANDOM_2875;
	logic [31:0] _RANDOM_2876;
	logic [31:0] _RANDOM_2877;
	logic [31:0] _RANDOM_2878;
	logic [31:0] _RANDOM_2879;
	logic [31:0] _RANDOM_2880;
	logic [31:0] _RANDOM_2881;
	logic [31:0] _RANDOM_2882;
	logic [31:0] _RANDOM_2883;
	logic [31:0] _RANDOM_2884;
	logic [31:0] _RANDOM_2885;
	logic [31:0] _RANDOM_2886;
	logic [31:0] _RANDOM_2887;
	logic [31:0] _RANDOM_2888;
	logic [31:0] _RANDOM_2889;
	logic [31:0] _RANDOM_2890;
	logic [31:0] _RANDOM_2891;
	logic [31:0] _RANDOM_2892;
	logic [31:0] _RANDOM_2893;
	logic [31:0] _RANDOM_2894;
	logic [31:0] _RANDOM_2895;
	logic [31:0] _RANDOM_2896;
	logic [31:0] _RANDOM_2897;
	logic [31:0] _RANDOM_2898;
	logic [31:0] _RANDOM_2899;
	logic [31:0] _RANDOM_2900;
	logic [31:0] _RANDOM_2901;
	logic [31:0] _RANDOM_2902;
	logic [31:0] _RANDOM_2903;
	logic [31:0] _RANDOM_2904;
	logic [31:0] _RANDOM_2905;
	logic [31:0] _RANDOM_2906;
	logic [31:0] _RANDOM_2907;
	logic [31:0] _RANDOM_2908;
	logic [31:0] _RANDOM_2909;
	logic [31:0] _RANDOM_2910;
	logic [31:0] _RANDOM_2911;
	logic [31:0] _RANDOM_2912;
	logic [31:0] _RANDOM_2913;
	logic [31:0] _RANDOM_2914;
	logic [31:0] _RANDOM_2915;
	logic [31:0] _RANDOM_2916;
	logic [31:0] _RANDOM_2917;
	logic [31:0] _RANDOM_2918;
	logic [31:0] _RANDOM_2919;
	logic [31:0] _RANDOM_2920;
	logic [31:0] _RANDOM_2921;
	logic [31:0] _RANDOM_2922;
	logic [31:0] _RANDOM_2923;
	logic [31:0] _RANDOM_2924;
	logic [31:0] _RANDOM_2925;
	logic [31:0] _RANDOM_2926;
	logic [31:0] _RANDOM_2927;
	logic [31:0] _RANDOM_2928;
	logic [31:0] _RANDOM_2929;
	logic [31:0] _RANDOM_2930;
	logic [31:0] _RANDOM_2931;
	logic [31:0] _RANDOM_2932;
	logic [31:0] _RANDOM_2933;
	logic [31:0] _RANDOM_2934;
	logic [31:0] _RANDOM_2935;
	logic [31:0] _RANDOM_2936;
	logic [31:0] _RANDOM_2937;
	logic [31:0] _RANDOM_2938;
	logic [31:0] _RANDOM_2939;
	logic [31:0] _RANDOM_2940;
	logic [31:0] _RANDOM_2941;
	logic [31:0] _RANDOM_2942;
	logic [31:0] _RANDOM_2943;
	logic [31:0] _RANDOM_2944;
	logic [31:0] _RANDOM_2945;
	logic [31:0] _RANDOM_2946;
	logic [31:0] _RANDOM_2947;
	logic [31:0] _RANDOM_2948;
	logic [31:0] _RANDOM_2949;
	logic [31:0] _RANDOM_2950;
	logic [31:0] _RANDOM_2951;
	logic [31:0] _RANDOM_2952;
	logic [31:0] _RANDOM_2953;
	logic [31:0] _RANDOM_2954;
	logic [31:0] _RANDOM_2955;
	logic [31:0] _RANDOM_2956;
	logic [31:0] _RANDOM_2957;
	logic [31:0] _RANDOM_2958;
	logic [31:0] _RANDOM_2959;
	logic [31:0] _RANDOM_2960;
	logic [31:0] _RANDOM_2961;
	logic [31:0] _RANDOM_2962;
	logic [31:0] _RANDOM_2963;
	logic [31:0] _RANDOM_2964;
	logic [31:0] _RANDOM_2965;
	logic [31:0] _RANDOM_2966;
	logic [31:0] _RANDOM_2967;
	logic [31:0] _RANDOM_2968;
	logic [31:0] _RANDOM_2969;
	logic [31:0] _RANDOM_2970;
	logic [31:0] _RANDOM_2971;
	logic [31:0] _RANDOM_2972;
	logic [31:0] _RANDOM_2973;
	logic [31:0] _RANDOM_2974;
	logic [31:0] _RANDOM_2975;
	logic [31:0] _RANDOM_2976;
	logic [31:0] _RANDOM_2977;
	logic [31:0] _RANDOM_2978;
	logic [31:0] _RANDOM_2979;
	logic [31:0] _RANDOM_2980;
	logic [31:0] _RANDOM_2981;
	logic [31:0] _RANDOM_2982;
	logic [31:0] _RANDOM_2983;
	logic [31:0] _RANDOM_2984;
	logic [31:0] _RANDOM_2985;
	logic [31:0] _RANDOM_2986;
	logic [31:0] _RANDOM_2987;
	logic [31:0] _RANDOM_2988;
	logic [31:0] _RANDOM_2989;
	logic [31:0] _RANDOM_2990;
	logic [31:0] _RANDOM_2991;
	logic [31:0] _RANDOM_2992;
	logic [31:0] _RANDOM_2993;
	logic [31:0] _RANDOM_2994;
	logic [31:0] _RANDOM_2995;
	logic [31:0] _RANDOM_2996;
	logic [31:0] _RANDOM_2997;
	logic [31:0] _RANDOM_2998;
	logic [31:0] _RANDOM_2999;
	logic [31:0] _RANDOM_3000;
	logic [31:0] _RANDOM_3001;
	logic [31:0] _RANDOM_3002;
	logic [31:0] _RANDOM_3003;
	logic [31:0] _RANDOM_3004;
	logic [31:0] _RANDOM_3005;
	logic [31:0] _RANDOM_3006;
	logic [31:0] _RANDOM_3007;
	logic [31:0] _RANDOM_3008;
	logic [31:0] _RANDOM_3009;
	logic [31:0] _RANDOM_3010;
	logic [31:0] _RANDOM_3011;
	logic [31:0] _RANDOM_3012;
	logic [31:0] _RANDOM_3013;
	logic [31:0] _RANDOM_3014;
	logic [31:0] _RANDOM_3015;
	logic [31:0] _RANDOM_3016;
	logic [31:0] _RANDOM_3017;
	logic [31:0] _RANDOM_3018;
	logic [31:0] _RANDOM_3019;
	logic [31:0] _RANDOM_3020;
	logic [31:0] _RANDOM_3021;
	logic [31:0] _RANDOM_3022;
	logic [31:0] _RANDOM_3023;
	logic [31:0] _RANDOM_3024;
	logic [31:0] _RANDOM_3025;
	logic [31:0] _RANDOM_3026;
	logic [31:0] _RANDOM_3027;
	logic [31:0] _RANDOM_3028;
	logic [31:0] _RANDOM_3029;
	logic [31:0] _RANDOM_3030;
	logic [31:0] _RANDOM_3031;
	logic [31:0] _RANDOM_3032;
	logic [31:0] _RANDOM_3033;
	logic [31:0] _RANDOM_3034;
	logic [31:0] _RANDOM_3035;
	logic [31:0] _RANDOM_3036;
	logic [31:0] _RANDOM_3037;
	logic [31:0] _RANDOM_3038;
	logic [31:0] _RANDOM_3039;
	logic [31:0] _RANDOM_3040;
	logic [31:0] _RANDOM_3041;
	logic [31:0] _RANDOM_3042;
	logic [31:0] _RANDOM_3043;
	logic [31:0] _RANDOM_3044;
	logic [31:0] _RANDOM_3045;
	logic [31:0] _RANDOM_3046;
	logic [31:0] _RANDOM_3047;
	logic [31:0] _RANDOM_3048;
	logic [31:0] _RANDOM_3049;
	logic [31:0] _RANDOM_3050;
	logic [31:0] _RANDOM_3051;
	logic [31:0] _RANDOM_3052;
	logic [31:0] _RANDOM_3053;
	logic [31:0] _RANDOM_3054;
	logic [31:0] _RANDOM_3055;
	logic [31:0] _RANDOM_3056;
	logic [31:0] _RANDOM_3057;
	logic [31:0] _RANDOM_3058;
	logic [31:0] _RANDOM_3059;
	logic [31:0] _RANDOM_3060;
	logic [31:0] _RANDOM_3061;
	logic [31:0] _RANDOM_3062;
	logic [31:0] _RANDOM_3063;
	logic [31:0] _RANDOM_3064;
	logic [31:0] _RANDOM_3065;
	logic [31:0] _RANDOM_3066;
	logic [31:0] _RANDOM_3067;
	logic [31:0] _RANDOM_3068;
	logic [31:0] _RANDOM_3069;
	logic [31:0] _RANDOM_3070;
	logic [31:0] _RANDOM_3071;
	logic [31:0] _RANDOM_3072;
	logic [31:0] _RANDOM_3073;
	logic [31:0] _RANDOM_3074;
	logic [31:0] _RANDOM_3075;
	logic [31:0] _RANDOM_3076;
	logic [31:0] _RANDOM_3077;
	logic [31:0] _RANDOM_3078;
	logic [31:0] _RANDOM_3079;
	logic [31:0] _RANDOM_3080;
	logic [31:0] _RANDOM_3081;
	logic [31:0] _RANDOM_3082;
	logic [31:0] _RANDOM_3083;
	logic [31:0] _RANDOM_3084;
	logic [31:0] _RANDOM_3085;
	logic [31:0] _RANDOM_3086;
	logic [31:0] _RANDOM_3087;
	logic [31:0] _RANDOM_3088;
	logic [31:0] _RANDOM_3089;
	logic [31:0] _RANDOM_3090;
	logic [31:0] _RANDOM_3091;
	logic [31:0] _RANDOM_3092;
	logic [31:0] _RANDOM_3093;
	logic [31:0] _RANDOM_3094;
	logic [31:0] _RANDOM_3095;
	logic [31:0] _RANDOM_3096;
	logic [31:0] _RANDOM_3097;
	logic [31:0] _RANDOM_3098;
	logic [31:0] _RANDOM_3099;
	logic [31:0] _RANDOM_3100;
	logic [31:0] _RANDOM_3101;
	logic [31:0] _RANDOM_3102;
	logic [31:0] _RANDOM_3103;
	logic [31:0] _RANDOM_3104;
	logic [31:0] _RANDOM_3105;
	logic [31:0] _RANDOM_3106;
	logic [31:0] _RANDOM_3107;
	logic [31:0] _RANDOM_3108;
	logic [31:0] _RANDOM_3109;
	logic [31:0] _RANDOM_3110;
	logic [31:0] _RANDOM_3111;
	logic [31:0] _RANDOM_3112;
	logic [31:0] _RANDOM_3113;
	logic [31:0] _RANDOM_3114;
	logic [31:0] _RANDOM_3115;
	logic [31:0] _RANDOM_3116;
	logic [31:0] _RANDOM_3117;
	logic [31:0] _RANDOM_3118;
	logic [31:0] _RANDOM_3119;
	logic [31:0] _RANDOM_3120;
	logic [31:0] _RANDOM_3121;
	logic [31:0] _RANDOM_3122;
	logic [31:0] _RANDOM_3123;
	logic [31:0] _RANDOM_3124;
	logic [31:0] _RANDOM_3125;
	logic [31:0] _RANDOM_3126;
	logic [31:0] _RANDOM_3127;
	logic [31:0] _RANDOM_3128;
	logic [31:0] _RANDOM_3129;
	logic [31:0] _RANDOM_3130;
	logic [31:0] _RANDOM_3131;
	logic [31:0] _RANDOM_3132;
	logic [31:0] _RANDOM_3133;
	logic [31:0] _RANDOM_3134;
	logic [31:0] _RANDOM_3135;
	logic [31:0] _RANDOM_3136;
	logic [31:0] _RANDOM_3137;
	logic [31:0] _RANDOM_3138;
	logic [31:0] _RANDOM_3139;
	logic [31:0] _RANDOM_3140;
	logic [31:0] _RANDOM_3141;
	logic [31:0] _RANDOM_3142;
	logic [31:0] _RANDOM_3143;
	logic [31:0] _RANDOM_3144;
	logic [31:0] _RANDOM_3145;
	logic [31:0] _RANDOM_3146;
	logic [31:0] _RANDOM_3147;
	logic [31:0] _RANDOM_3148;
	logic [31:0] _RANDOM_3149;
	logic [31:0] _RANDOM_3150;
	logic [31:0] _RANDOM_3151;
	logic [31:0] _RANDOM_3152;
	logic [31:0] _RANDOM_3153;
	logic [31:0] _RANDOM_3154;
	logic [31:0] _RANDOM_3155;
	logic [31:0] _RANDOM_3156;
	logic [31:0] _RANDOM_3157;
	logic [31:0] _RANDOM_3158;
	logic [31:0] _RANDOM_3159;
	logic [31:0] _RANDOM_3160;
	logic [31:0] _RANDOM_3161;
	logic [31:0] _RANDOM_3162;
	logic [31:0] _RANDOM_3163;
	logic [31:0] _RANDOM_3164;
	logic [31:0] _RANDOM_3165;
	logic [31:0] _RANDOM_3166;
	logic [31:0] _RANDOM_3167;
	logic [31:0] _RANDOM_3168;
	logic [31:0] _RANDOM_3169;
	logic [31:0] _RANDOM_3170;
	logic [31:0] _RANDOM_3171;
	logic [31:0] _RANDOM_3172;
	logic [31:0] _RANDOM_3173;
	logic [31:0] _RANDOM_3174;
	logic [31:0] _RANDOM_3175;
	logic [31:0] _RANDOM_3176;
	logic [31:0] _RANDOM_3177;
	logic [31:0] _RANDOM_3178;
	logic [31:0] _RANDOM_3179;
	logic [31:0] _RANDOM_3180;
	logic [31:0] _RANDOM_3181;
	logic [31:0] _RANDOM_3182;
	logic [31:0] _RANDOM_3183;
	logic [31:0] _RANDOM_3184;
	logic [31:0] _RANDOM_3185;
	logic [31:0] _RANDOM_3186;
	logic [31:0] _RANDOM_3187;
	logic [31:0] _RANDOM_3188;
	logic [31:0] _RANDOM_3189;
	logic [31:0] _RANDOM_3190;
	logic [31:0] _RANDOM_3191;
	logic [31:0] _RANDOM_3192;
	logic [31:0] _RANDOM_3193;
	logic [31:0] _RANDOM_3194;
	logic [31:0] _RANDOM_3195;
	logic [31:0] _RANDOM_3196;
	logic [31:0] _RANDOM_3197;
	logic [31:0] _RANDOM_3198;
	logic [31:0] _RANDOM_3199;
	logic [31:0] _RANDOM_3200;
	logic [31:0] _RANDOM_3201;
	logic [31:0] _RANDOM_3202;
	logic [31:0] _RANDOM_3203;
	logic [31:0] _RANDOM_3204;
	logic [31:0] _RANDOM_3205;
	logic [31:0] _RANDOM_3206;
	logic [31:0] _RANDOM_3207;
	logic [31:0] _RANDOM_3208;
	logic [31:0] _RANDOM_3209;
	logic [31:0] _RANDOM_3210;
	logic [31:0] _RANDOM_3211;
	logic [31:0] _RANDOM_3212;
	logic [31:0] _RANDOM_3213;
	logic [31:0] _RANDOM_3214;
	logic [31:0] _RANDOM_3215;
	logic [31:0] _RANDOM_3216;
	logic [31:0] _RANDOM_3217;
	logic [31:0] _RANDOM_3218;
	logic [31:0] _RANDOM_3219;
	logic [31:0] _RANDOM_3220;
	logic [31:0] _RANDOM_3221;
	logic [31:0] _RANDOM_3222;
	logic [31:0] _RANDOM_3223;
	logic [31:0] _RANDOM_3224;
	logic [31:0] _RANDOM_3225;
	logic [31:0] _RANDOM_3226;
	logic [31:0] _RANDOM_3227;
	logic [31:0] _RANDOM_3228;
	logic [31:0] _RANDOM_3229;
	logic [31:0] _RANDOM_3230;
	logic [31:0] _RANDOM_3231;
	logic [31:0] _RANDOM_3232;
	logic [31:0] _RANDOM_3233;
	logic [31:0] _RANDOM_3234;
	logic [31:0] _RANDOM_3235;
	logic [31:0] _RANDOM_3236;
	logic [31:0] _RANDOM_3237;
	logic [31:0] _RANDOM_3238;
	logic [31:0] _RANDOM_3239;
	logic [31:0] _RANDOM_3240;
	logic [31:0] _RANDOM_3241;
	logic [31:0] _RANDOM_3242;
	logic [31:0] _RANDOM_3243;
	logic [31:0] _RANDOM_3244;
	logic [31:0] _RANDOM_3245;
	logic [31:0] _RANDOM_3246;
	logic [31:0] _RANDOM_3247;
	logic [31:0] _RANDOM_3248;
	logic [31:0] _RANDOM_3249;
	logic [31:0] _RANDOM_3250;
	logic [31:0] _RANDOM_3251;
	logic [31:0] _RANDOM_3252;
	logic [31:0] _RANDOM_3253;
	logic [31:0] _RANDOM_3254;
	logic [31:0] _RANDOM_3255;
	logic [31:0] _RANDOM_3256;
	logic [31:0] _RANDOM_3257;
	logic [31:0] _RANDOM_3258;
	logic [31:0] _RANDOM_3259;
	logic [31:0] _RANDOM_3260;
	logic [31:0] _RANDOM_3261;
	logic [31:0] _RANDOM_3262;
	logic [31:0] _RANDOM_3263;
	logic [31:0] _RANDOM_3264;
	logic [31:0] _RANDOM_3265;
	logic [31:0] _RANDOM_3266;
	logic [31:0] _RANDOM_3267;
	logic [31:0] _RANDOM_3268;
	logic [31:0] _RANDOM_3269;
	logic [31:0] _RANDOM_3270;
	logic [31:0] _RANDOM_3271;
	logic [31:0] _RANDOM_3272;
	logic [31:0] _RANDOM_3273;
	logic [31:0] _RANDOM_3274;
	logic [31:0] _RANDOM_3275;
	logic [31:0] _RANDOM_3276;
	logic [31:0] _RANDOM_3277;
	logic [31:0] _RANDOM_3278;
	logic [31:0] _RANDOM_3279;
	logic [31:0] _RANDOM_3280;
	logic [31:0] _RANDOM_3281;
	logic [31:0] _RANDOM_3282;
	logic [31:0] _RANDOM_3283;
	logic [31:0] _RANDOM_3284;
	logic [31:0] _RANDOM_3285;
	logic [31:0] _RANDOM_3286;
	logic [31:0] _RANDOM_3287;
	logic [31:0] _RANDOM_3288;
	logic [31:0] _RANDOM_3289;
	logic [31:0] _RANDOM_3290;
	logic [31:0] _RANDOM_3291;
	logic [31:0] _RANDOM_3292;
	logic [31:0] _RANDOM_3293;
	logic [31:0] _RANDOM_3294;
	logic [31:0] _RANDOM_3295;
	logic [31:0] _RANDOM_3296;
	logic [31:0] _RANDOM_3297;
	logic [31:0] _RANDOM_3298;
	logic [31:0] _RANDOM_3299;
	logic [31:0] _RANDOM_3300;
	logic [31:0] _RANDOM_3301;
	logic [31:0] _RANDOM_3302;
	logic [31:0] _RANDOM_3303;
	logic [31:0] _RANDOM_3304;
	logic [31:0] _RANDOM_3305;
	logic [31:0] _RANDOM_3306;
	logic [31:0] _RANDOM_3307;
	logic [31:0] _RANDOM_3308;
	logic [31:0] _RANDOM_3309;
	logic [31:0] _RANDOM_3310;
	logic [31:0] _RANDOM_3311;
	logic [31:0] _RANDOM_3312;
	logic [31:0] _RANDOM_3313;
	logic [31:0] _RANDOM_3314;
	logic [31:0] _RANDOM_3315;
	logic [31:0] _RANDOM_3316;
	logic [31:0] _RANDOM_3317;
	logic [31:0] _RANDOM_3318;
	logic [31:0] _RANDOM_3319;
	logic [31:0] _RANDOM_3320;
	logic [31:0] _RANDOM_3321;
	logic [31:0] _RANDOM_3322;
	logic [31:0] _RANDOM_3323;
	logic [31:0] _RANDOM_3324;
	logic [31:0] _RANDOM_3325;
	logic [31:0] _RANDOM_3326;
	logic [31:0] _RANDOM_3327;
	logic [31:0] _RANDOM_3328;
	logic [31:0] _RANDOM_3329;
	logic [31:0] _RANDOM_3330;
	logic [31:0] _RANDOM_3331;
	logic [31:0] _RANDOM_3332;
	logic [31:0] _RANDOM_3333;
	logic [31:0] _RANDOM_3334;
	logic [31:0] _RANDOM_3335;
	logic [31:0] _RANDOM_3336;
	logic [31:0] _RANDOM_3337;
	logic [31:0] _RANDOM_3338;
	logic [31:0] _RANDOM_3339;
	logic [31:0] _RANDOM_3340;
	logic [31:0] _RANDOM_3341;
	logic [31:0] _RANDOM_3342;
	logic [31:0] _RANDOM_3343;
	logic [31:0] _RANDOM_3344;
	logic [31:0] _RANDOM_3345;
	logic [31:0] _RANDOM_3346;
	logic [31:0] _RANDOM_3347;
	logic [31:0] _RANDOM_3348;
	logic [31:0] _RANDOM_3349;
	logic [31:0] _RANDOM_3350;
	logic [31:0] _RANDOM_3351;
	logic [31:0] _RANDOM_3352;
	logic [31:0] _RANDOM_3353;
	logic [31:0] _RANDOM_3354;
	logic [31:0] _RANDOM_3355;
	logic [31:0] _RANDOM_3356;
	logic [31:0] _RANDOM_3357;
	logic [31:0] _RANDOM_3358;
	logic [31:0] _RANDOM_3359;
	logic [31:0] _RANDOM_3360;
	logic [31:0] _RANDOM_3361;
	logic [31:0] _RANDOM_3362;
	logic [31:0] _RANDOM_3363;
	logic [31:0] _RANDOM_3364;
	logic [31:0] _RANDOM_3365;
	logic [31:0] _RANDOM_3366;
	logic [31:0] _RANDOM_3367;
	logic [31:0] _RANDOM_3368;
	logic [31:0] _RANDOM_3369;
	logic [31:0] _RANDOM_3370;
	logic [31:0] _RANDOM_3371;
	logic [31:0] _RANDOM_3372;
	logic [31:0] _RANDOM_3373;
	logic [31:0] _RANDOM_3374;
	logic [31:0] _RANDOM_3375;
	logic [31:0] _RANDOM_3376;
	logic [31:0] _RANDOM_3377;
	logic [31:0] _RANDOM_3378;
	logic [31:0] _RANDOM_3379;
	logic [31:0] _RANDOM_3380;
	logic [31:0] _RANDOM_3381;
	logic [31:0] _RANDOM_3382;
	logic [31:0] _RANDOM_3383;
	logic [31:0] _RANDOM_3384;
	logic [31:0] _RANDOM_3385;
	logic [31:0] _RANDOM_3386;
	logic [31:0] _RANDOM_3387;
	logic [31:0] _RANDOM_3388;
	logic [31:0] _RANDOM_3389;
	logic [31:0] _RANDOM_3390;
	logic [31:0] _RANDOM_3391;
	logic [31:0] _RANDOM_3392;
	logic [31:0] _RANDOM_3393;
	logic [31:0] _RANDOM_3394;
	logic [31:0] _RANDOM_3395;
	logic [31:0] _RANDOM_3396;
	logic [31:0] _RANDOM_3397;
	logic [31:0] _RANDOM_3398;
	logic [31:0] _RANDOM_3399;
	logic [31:0] _RANDOM_3400;
	logic [31:0] _RANDOM_3401;
	logic [31:0] _RANDOM_3402;
	logic [31:0] _RANDOM_3403;
	logic [31:0] _RANDOM_3404;
	logic [31:0] _RANDOM_3405;
	logic [31:0] _RANDOM_3406;
	logic [31:0] _RANDOM_3407;
	logic [31:0] _RANDOM_3408;
	logic [31:0] _RANDOM_3409;
	logic [31:0] _RANDOM_3410;
	logic [31:0] _RANDOM_3411;
	logic [31:0] _RANDOM_3412;
	logic [31:0] _RANDOM_3413;
	logic [31:0] _RANDOM_3414;
	logic [31:0] _RANDOM_3415;
	logic [31:0] _RANDOM_3416;
	logic [31:0] _RANDOM_3417;
	logic [31:0] _RANDOM_3418;
	logic [31:0] _RANDOM_3419;
	logic [31:0] _RANDOM_3420;
	logic [31:0] _RANDOM_3421;
	logic [31:0] _RANDOM_3422;
	logic [31:0] _RANDOM_3423;
	logic [31:0] _RANDOM_3424;
	logic [31:0] _RANDOM_3425;
	logic [31:0] _RANDOM_3426;
	logic [31:0] _RANDOM_3427;
	logic [31:0] _RANDOM_3428;
	logic [31:0] _RANDOM_3429;
	logic [31:0] _RANDOM_3430;
	logic [31:0] _RANDOM_3431;
	logic [31:0] _RANDOM_3432;
	logic [31:0] _RANDOM_3433;
	logic [31:0] _RANDOM_3434;
	logic [31:0] _RANDOM_3435;
	logic [31:0] _RANDOM_3436;
	logic [31:0] _RANDOM_3437;
	logic [31:0] _RANDOM_3438;
	logic [31:0] _RANDOM_3439;
	logic [31:0] _RANDOM_3440;
	logic [31:0] _RANDOM_3441;
	logic [31:0] _RANDOM_3442;
	logic [31:0] _RANDOM_3443;
	logic [31:0] _RANDOM_3444;
	logic [31:0] _RANDOM_3445;
	logic [31:0] _RANDOM_3446;
	logic [31:0] _RANDOM_3447;
	logic [31:0] _RANDOM_3448;
	logic [31:0] _RANDOM_3449;
	logic [31:0] _RANDOM_3450;
	logic [31:0] _RANDOM_3451;
	logic [31:0] _RANDOM_3452;
	logic [31:0] _RANDOM_3453;
	logic [31:0] _RANDOM_3454;
	logic [31:0] _RANDOM_3455;
	logic [31:0] _RANDOM_3456;
	logic [31:0] _RANDOM_3457;
	logic [31:0] _RANDOM_3458;
	logic [31:0] _RANDOM_3459;
	logic [31:0] _RANDOM_3460;
	logic [31:0] _RANDOM_3461;
	logic [31:0] _RANDOM_3462;
	logic [31:0] _RANDOM_3463;
	logic [31:0] _RANDOM_3464;
	logic [31:0] _RANDOM_3465;
	logic [31:0] _RANDOM_3466;
	logic [31:0] _RANDOM_3467;
	logic [31:0] _RANDOM_3468;
	logic [31:0] _RANDOM_3469;
	logic [31:0] _RANDOM_3470;
	logic [31:0] _RANDOM_3471;
	logic [31:0] _RANDOM_3472;
	logic [31:0] _RANDOM_3473;
	logic [31:0] _RANDOM_3474;
	logic [31:0] _RANDOM_3475;
	logic [31:0] _RANDOM_3476;
	logic [31:0] _RANDOM_3477;
	logic [31:0] _RANDOM_3478;
	logic [31:0] _RANDOM_3479;
	logic [31:0] _RANDOM_3480;
	logic [31:0] _RANDOM_3481;
	logic [31:0] _RANDOM_3482;
	logic [31:0] _RANDOM_3483;
	logic [31:0] _RANDOM_3484;
	logic [31:0] _RANDOM_3485;
	logic [31:0] _RANDOM_3486;
	logic [31:0] _RANDOM_3487;
	logic [31:0] _RANDOM_3488;
	logic [31:0] _RANDOM_3489;
	logic [31:0] _RANDOM_3490;
	logic [31:0] _RANDOM_3491;
	logic [31:0] _RANDOM_3492;
	logic [31:0] _RANDOM_3493;
	logic [31:0] _RANDOM_3494;
	logic [31:0] _RANDOM_3495;
	logic [31:0] _RANDOM_3496;
	logic [31:0] _RANDOM_3497;
	logic [31:0] _RANDOM_3498;
	logic [31:0] _RANDOM_3499;
	logic [31:0] _RANDOM_3500;
	logic [31:0] _RANDOM_3501;
	logic [31:0] _RANDOM_3502;
	logic [31:0] _RANDOM_3503;
	logic [31:0] _RANDOM_3504;
	logic [31:0] _RANDOM_3505;
	logic [31:0] _RANDOM_3506;
	logic [31:0] _RANDOM_3507;
	logic [31:0] _RANDOM_3508;
	logic [31:0] _RANDOM_3509;
	logic [31:0] _RANDOM_3510;
	logic [31:0] _RANDOM_3511;
	logic [31:0] _RANDOM_3512;
	logic [31:0] _RANDOM_3513;
	logic [31:0] _RANDOM_3514;
	logic [31:0] _RANDOM_3515;
	logic [31:0] _RANDOM_3516;
	logic [31:0] _RANDOM_3517;
	logic [31:0] _RANDOM_3518;
	logic [31:0] _RANDOM_3519;
	logic [31:0] _RANDOM_3520;
	logic [31:0] _RANDOM_3521;
	logic [31:0] _RANDOM_3522;
	logic [31:0] _RANDOM_3523;
	logic [31:0] _RANDOM_3524;
	logic [31:0] _RANDOM_3525;
	logic [31:0] _RANDOM_3526;
	logic [31:0] _RANDOM_3527;
	logic [31:0] _RANDOM_3528;
	logic [31:0] _RANDOM_3529;
	logic [31:0] _RANDOM_3530;
	logic [31:0] _RANDOM_3531;
	logic [31:0] _RANDOM_3532;
	logic [31:0] _RANDOM_3533;
	logic [31:0] _RANDOM_3534;
	logic [31:0] _RANDOM_3535;
	logic [31:0] _RANDOM_3536;
	logic [31:0] _RANDOM_3537;
	logic [31:0] _RANDOM_3538;
	logic [31:0] _RANDOM_3539;
	logic [31:0] _RANDOM_3540;
	logic [31:0] _RANDOM_3541;
	logic [31:0] _RANDOM_3542;
	logic [31:0] _RANDOM_3543;
	logic [31:0] _RANDOM_3544;
	logic [31:0] _RANDOM_3545;
	logic [31:0] _RANDOM_3546;
	logic [31:0] _RANDOM_3547;
	logic [31:0] _RANDOM_3548;
	logic [31:0] _RANDOM_3549;
	logic [31:0] _RANDOM_3550;
	logic [31:0] _RANDOM_3551;
	logic [31:0] _RANDOM_3552;
	logic [31:0] _RANDOM_3553;
	logic [31:0] _RANDOM_3554;
	logic [31:0] _RANDOM_3555;
	logic [31:0] _RANDOM_3556;
	logic [31:0] _RANDOM_3557;
	logic [31:0] _RANDOM_3558;
	logic [31:0] _RANDOM_3559;
	logic [31:0] _RANDOM_3560;
	logic [31:0] _RANDOM_3561;
	logic [31:0] _RANDOM_3562;
	logic [31:0] _RANDOM_3563;
	logic [31:0] _RANDOM_3564;
	logic [31:0] _RANDOM_3565;
	logic [31:0] _RANDOM_3566;
	logic [31:0] _RANDOM_3567;
	logic [31:0] _RANDOM_3568;
	logic [31:0] _RANDOM_3569;
	logic [31:0] _RANDOM_3570;
	logic [31:0] _RANDOM_3571;
	logic [31:0] _RANDOM_3572;
	logic [31:0] _RANDOM_3573;
	logic [31:0] _RANDOM_3574;
	logic [31:0] _RANDOM_3575;
	logic [31:0] _RANDOM_3576;
	logic [31:0] _RANDOM_3577;
	logic [31:0] _RANDOM_3578;
	logic [31:0] _RANDOM_3579;
	logic [31:0] _RANDOM_3580;
	logic [31:0] _RANDOM_3581;
	logic [31:0] _RANDOM_3582;
	logic [31:0] _RANDOM_3583;
	logic [31:0] _RANDOM_3584;
	logic [31:0] _RANDOM_3585;
	logic [31:0] _RANDOM_3586;
	logic [31:0] _RANDOM_3587;
	logic [31:0] _RANDOM_3588;
	logic [31:0] _RANDOM_3589;
	logic [31:0] _RANDOM_3590;
	logic [31:0] _RANDOM_3591;
	logic [31:0] _RANDOM_3592;
	logic [31:0] _RANDOM_3593;
	logic [31:0] _RANDOM_3594;
	logic [31:0] _RANDOM_3595;
	logic [31:0] _RANDOM_3596;
	logic [31:0] _RANDOM_3597;
	logic [31:0] _RANDOM_3598;
	logic [31:0] _RANDOM_3599;
	logic [31:0] _RANDOM_3600;
	logic [31:0] _RANDOM_3601;
	logic [31:0] _RANDOM_3602;
	logic [31:0] _RANDOM_3603;
	logic [31:0] _RANDOM_3604;
	logic [31:0] _RANDOM_3605;
	logic [31:0] _RANDOM_3606;
	logic [31:0] _RANDOM_3607;
	logic [31:0] _RANDOM_3608;
	logic [31:0] _RANDOM_3609;
	logic [31:0] _RANDOM_3610;
	logic [31:0] _RANDOM_3611;
	logic [31:0] _RANDOM_3612;
	logic [31:0] _RANDOM_3613;
	logic [31:0] _RANDOM_3614;
	logic [31:0] _RANDOM_3615;
	logic [31:0] _RANDOM_3616;
	logic [31:0] _RANDOM_3617;
	logic [31:0] _RANDOM_3618;
	logic [31:0] _RANDOM_3619;
	logic [31:0] _RANDOM_3620;
	logic [31:0] _RANDOM_3621;
	logic [31:0] _RANDOM_3622;
	logic [31:0] _RANDOM_3623;
	logic [31:0] _RANDOM_3624;
	logic [31:0] _RANDOM_3625;
	logic [31:0] _RANDOM_3626;
	logic [31:0] _RANDOM_3627;
	logic [31:0] _RANDOM_3628;
	logic [31:0] _RANDOM_3629;
	logic [31:0] _RANDOM_3630;
	logic [31:0] _RANDOM_3631;
	logic [31:0] _RANDOM_3632;
	logic [31:0] _RANDOM_3633;
	logic [31:0] _RANDOM_3634;
	logic [31:0] _RANDOM_3635;
	logic [31:0] _RANDOM_3636;
	logic [31:0] _RANDOM_3637;
	logic [31:0] _RANDOM_3638;
	logic [31:0] _RANDOM_3639;
	logic [31:0] _RANDOM_3640;
	logic [31:0] _RANDOM_3641;
	logic [31:0] _RANDOM_3642;
	logic [31:0] _RANDOM_3643;
	logic [31:0] _RANDOM_3644;
	logic [31:0] _RANDOM_3645;
	logic [31:0] _RANDOM_3646;
	logic [31:0] _RANDOM_3647;
	logic [31:0] _RANDOM_3648;
	logic [31:0] _RANDOM_3649;
	logic [31:0] _RANDOM_3650;
	logic [31:0] _RANDOM_3651;
	logic [31:0] _RANDOM_3652;
	logic [31:0] _RANDOM_3653;
	logic [31:0] _RANDOM_3654;
	logic [31:0] _RANDOM_3655;
	logic [31:0] _RANDOM_3656;
	logic [31:0] _RANDOM_3657;
	logic [31:0] _RANDOM_3658;
	logic [31:0] _RANDOM_3659;
	logic [31:0] _RANDOM_3660;
	logic [31:0] _RANDOM_3661;
	logic [31:0] _RANDOM_3662;
	logic [31:0] _RANDOM_3663;
	logic [31:0] _RANDOM_3664;
	logic [31:0] _RANDOM_3665;
	logic [31:0] _RANDOM_3666;
	logic [31:0] _RANDOM_3667;
	logic [31:0] _RANDOM_3668;
	logic [31:0] _RANDOM_3669;
	logic [31:0] _RANDOM_3670;
	logic [31:0] _RANDOM_3671;
	logic [31:0] _RANDOM_3672;
	logic [31:0] _RANDOM_3673;
	logic [31:0] _RANDOM_3674;
	logic [31:0] _RANDOM_3675;
	logic [31:0] _RANDOM_3676;
	logic [31:0] _RANDOM_3677;
	logic [31:0] _RANDOM_3678;
	logic [31:0] _RANDOM_3679;
	logic [31:0] _RANDOM_3680;
	logic [31:0] _RANDOM_3681;
	logic [31:0] _RANDOM_3682;
	logic [31:0] _RANDOM_3683;
	logic [31:0] _RANDOM_3684;
	logic [31:0] _RANDOM_3685;
	logic [31:0] _RANDOM_3686;
	logic [31:0] _RANDOM_3687;
	logic [31:0] _RANDOM_3688;
	logic [31:0] _RANDOM_3689;
	logic [31:0] _RANDOM_3690;
	logic [31:0] _RANDOM_3691;
	Tile mesh_0_0(
		.clock(clock),
		.io_in_a_0(r_0),
		.io_in_b_0(b_0),
		.io_in_d_0(b_1024_0),
		.io_in_control_0_dataflow(mesh_0_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2048_0),
		.io_in_last_0(r_3072_0),
		.io_in_valid_0(r_1024_0),
		.io_out_a_0(_mesh_0_0_io_out_a_0),
		.io_out_c_0(_mesh_0_0_io_out_c_0),
		.io_out_b_0(_mesh_0_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_0_io_out_id_0),
		.io_out_last_0(_mesh_0_0_io_out_last_0),
		.io_out_valid_0(_mesh_0_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9371 == GlobalFiModInstNr[0]) || (9371 == GlobalFiModInstNr[1]) || (9371 == GlobalFiModInstNr[2]) || (9371 == GlobalFiModInstNr[3]))));
	Tile mesh_0_1(
		.clock(clock),
		.io_in_a_0(r_1_0),
		.io_in_b_0(b_32_0),
		.io_in_d_0(b_1056_0),
		.io_in_control_0_dataflow(mesh_0_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2080_0),
		.io_in_last_0(r_3104_0),
		.io_in_valid_0(r_1056_0),
		.io_out_a_0(_mesh_0_1_io_out_a_0),
		.io_out_c_0(_mesh_0_1_io_out_c_0),
		.io_out_b_0(_mesh_0_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_1_io_out_id_0),
		.io_out_last_0(_mesh_0_1_io_out_last_0),
		.io_out_valid_0(_mesh_0_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9372 == GlobalFiModInstNr[0]) || (9372 == GlobalFiModInstNr[1]) || (9372 == GlobalFiModInstNr[2]) || (9372 == GlobalFiModInstNr[3]))));
	Tile mesh_0_2(
		.clock(clock),
		.io_in_a_0(r_2_0),
		.io_in_b_0(b_64_0),
		.io_in_d_0(b_1088_0),
		.io_in_control_0_dataflow(mesh_0_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2112_0),
		.io_in_last_0(r_3136_0),
		.io_in_valid_0(r_1088_0),
		.io_out_a_0(_mesh_0_2_io_out_a_0),
		.io_out_c_0(_mesh_0_2_io_out_c_0),
		.io_out_b_0(_mesh_0_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_2_io_out_id_0),
		.io_out_last_0(_mesh_0_2_io_out_last_0),
		.io_out_valid_0(_mesh_0_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9373 == GlobalFiModInstNr[0]) || (9373 == GlobalFiModInstNr[1]) || (9373 == GlobalFiModInstNr[2]) || (9373 == GlobalFiModInstNr[3]))));
	Tile mesh_0_3(
		.clock(clock),
		.io_in_a_0(r_3_0),
		.io_in_b_0(b_96_0),
		.io_in_d_0(b_1120_0),
		.io_in_control_0_dataflow(mesh_0_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2144_0),
		.io_in_last_0(r_3168_0),
		.io_in_valid_0(r_1120_0),
		.io_out_a_0(_mesh_0_3_io_out_a_0),
		.io_out_c_0(_mesh_0_3_io_out_c_0),
		.io_out_b_0(_mesh_0_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_3_io_out_id_0),
		.io_out_last_0(_mesh_0_3_io_out_last_0),
		.io_out_valid_0(_mesh_0_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9374 == GlobalFiModInstNr[0]) || (9374 == GlobalFiModInstNr[1]) || (9374 == GlobalFiModInstNr[2]) || (9374 == GlobalFiModInstNr[3]))));
	Tile mesh_0_4(
		.clock(clock),
		.io_in_a_0(r_4_0),
		.io_in_b_0(b_128_0),
		.io_in_d_0(b_1152_0),
		.io_in_control_0_dataflow(mesh_0_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2176_0),
		.io_in_last_0(r_3200_0),
		.io_in_valid_0(r_1152_0),
		.io_out_a_0(_mesh_0_4_io_out_a_0),
		.io_out_c_0(_mesh_0_4_io_out_c_0),
		.io_out_b_0(_mesh_0_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_4_io_out_id_0),
		.io_out_last_0(_mesh_0_4_io_out_last_0),
		.io_out_valid_0(_mesh_0_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9375 == GlobalFiModInstNr[0]) || (9375 == GlobalFiModInstNr[1]) || (9375 == GlobalFiModInstNr[2]) || (9375 == GlobalFiModInstNr[3]))));
	Tile mesh_0_5(
		.clock(clock),
		.io_in_a_0(r_5_0),
		.io_in_b_0(b_160_0),
		.io_in_d_0(b_1184_0),
		.io_in_control_0_dataflow(mesh_0_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2208_0),
		.io_in_last_0(r_3232_0),
		.io_in_valid_0(r_1184_0),
		.io_out_a_0(_mesh_0_5_io_out_a_0),
		.io_out_c_0(_mesh_0_5_io_out_c_0),
		.io_out_b_0(_mesh_0_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_5_io_out_id_0),
		.io_out_last_0(_mesh_0_5_io_out_last_0),
		.io_out_valid_0(_mesh_0_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9376 == GlobalFiModInstNr[0]) || (9376 == GlobalFiModInstNr[1]) || (9376 == GlobalFiModInstNr[2]) || (9376 == GlobalFiModInstNr[3]))));
	Tile mesh_0_6(
		.clock(clock),
		.io_in_a_0(r_6_0),
		.io_in_b_0(b_192_0),
		.io_in_d_0(b_1216_0),
		.io_in_control_0_dataflow(mesh_0_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2240_0),
		.io_in_last_0(r_3264_0),
		.io_in_valid_0(r_1216_0),
		.io_out_a_0(_mesh_0_6_io_out_a_0),
		.io_out_c_0(_mesh_0_6_io_out_c_0),
		.io_out_b_0(_mesh_0_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_6_io_out_id_0),
		.io_out_last_0(_mesh_0_6_io_out_last_0),
		.io_out_valid_0(_mesh_0_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9377 == GlobalFiModInstNr[0]) || (9377 == GlobalFiModInstNr[1]) || (9377 == GlobalFiModInstNr[2]) || (9377 == GlobalFiModInstNr[3]))));
	Tile mesh_0_7(
		.clock(clock),
		.io_in_a_0(r_7_0),
		.io_in_b_0(b_224_0),
		.io_in_d_0(b_1248_0),
		.io_in_control_0_dataflow(mesh_0_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2272_0),
		.io_in_last_0(r_3296_0),
		.io_in_valid_0(r_1248_0),
		.io_out_a_0(_mesh_0_7_io_out_a_0),
		.io_out_c_0(_mesh_0_7_io_out_c_0),
		.io_out_b_0(_mesh_0_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_7_io_out_id_0),
		.io_out_last_0(_mesh_0_7_io_out_last_0),
		.io_out_valid_0(_mesh_0_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9378 == GlobalFiModInstNr[0]) || (9378 == GlobalFiModInstNr[1]) || (9378 == GlobalFiModInstNr[2]) || (9378 == GlobalFiModInstNr[3]))));
	Tile mesh_0_8(
		.clock(clock),
		.io_in_a_0(r_8_0),
		.io_in_b_0(b_256_0),
		.io_in_d_0(b_1280_0),
		.io_in_control_0_dataflow(mesh_0_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2304_0),
		.io_in_last_0(r_3328_0),
		.io_in_valid_0(r_1280_0),
		.io_out_a_0(_mesh_0_8_io_out_a_0),
		.io_out_c_0(_mesh_0_8_io_out_c_0),
		.io_out_b_0(_mesh_0_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_8_io_out_id_0),
		.io_out_last_0(_mesh_0_8_io_out_last_0),
		.io_out_valid_0(_mesh_0_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9379 == GlobalFiModInstNr[0]) || (9379 == GlobalFiModInstNr[1]) || (9379 == GlobalFiModInstNr[2]) || (9379 == GlobalFiModInstNr[3]))));
	Tile mesh_0_9(
		.clock(clock),
		.io_in_a_0(r_9_0),
		.io_in_b_0(b_288_0),
		.io_in_d_0(b_1312_0),
		.io_in_control_0_dataflow(mesh_0_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2336_0),
		.io_in_last_0(r_3360_0),
		.io_in_valid_0(r_1312_0),
		.io_out_a_0(_mesh_0_9_io_out_a_0),
		.io_out_c_0(_mesh_0_9_io_out_c_0),
		.io_out_b_0(_mesh_0_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_9_io_out_id_0),
		.io_out_last_0(_mesh_0_9_io_out_last_0),
		.io_out_valid_0(_mesh_0_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9380 == GlobalFiModInstNr[0]) || (9380 == GlobalFiModInstNr[1]) || (9380 == GlobalFiModInstNr[2]) || (9380 == GlobalFiModInstNr[3]))));
	Tile mesh_0_10(
		.clock(clock),
		.io_in_a_0(r_10_0),
		.io_in_b_0(b_320_0),
		.io_in_d_0(b_1344_0),
		.io_in_control_0_dataflow(mesh_0_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2368_0),
		.io_in_last_0(r_3392_0),
		.io_in_valid_0(r_1344_0),
		.io_out_a_0(_mesh_0_10_io_out_a_0),
		.io_out_c_0(_mesh_0_10_io_out_c_0),
		.io_out_b_0(_mesh_0_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_10_io_out_id_0),
		.io_out_last_0(_mesh_0_10_io_out_last_0),
		.io_out_valid_0(_mesh_0_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9381 == GlobalFiModInstNr[0]) || (9381 == GlobalFiModInstNr[1]) || (9381 == GlobalFiModInstNr[2]) || (9381 == GlobalFiModInstNr[3]))));
	Tile mesh_0_11(
		.clock(clock),
		.io_in_a_0(r_11_0),
		.io_in_b_0(b_352_0),
		.io_in_d_0(b_1376_0),
		.io_in_control_0_dataflow(mesh_0_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2400_0),
		.io_in_last_0(r_3424_0),
		.io_in_valid_0(r_1376_0),
		.io_out_a_0(_mesh_0_11_io_out_a_0),
		.io_out_c_0(_mesh_0_11_io_out_c_0),
		.io_out_b_0(_mesh_0_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_11_io_out_id_0),
		.io_out_last_0(_mesh_0_11_io_out_last_0),
		.io_out_valid_0(_mesh_0_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9382 == GlobalFiModInstNr[0]) || (9382 == GlobalFiModInstNr[1]) || (9382 == GlobalFiModInstNr[2]) || (9382 == GlobalFiModInstNr[3]))));
	Tile mesh_0_12(
		.clock(clock),
		.io_in_a_0(r_12_0),
		.io_in_b_0(b_384_0),
		.io_in_d_0(b_1408_0),
		.io_in_control_0_dataflow(mesh_0_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2432_0),
		.io_in_last_0(r_3456_0),
		.io_in_valid_0(r_1408_0),
		.io_out_a_0(_mesh_0_12_io_out_a_0),
		.io_out_c_0(_mesh_0_12_io_out_c_0),
		.io_out_b_0(_mesh_0_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_12_io_out_id_0),
		.io_out_last_0(_mesh_0_12_io_out_last_0),
		.io_out_valid_0(_mesh_0_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9383 == GlobalFiModInstNr[0]) || (9383 == GlobalFiModInstNr[1]) || (9383 == GlobalFiModInstNr[2]) || (9383 == GlobalFiModInstNr[3]))));
	Tile mesh_0_13(
		.clock(clock),
		.io_in_a_0(r_13_0),
		.io_in_b_0(b_416_0),
		.io_in_d_0(b_1440_0),
		.io_in_control_0_dataflow(mesh_0_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2464_0),
		.io_in_last_0(r_3488_0),
		.io_in_valid_0(r_1440_0),
		.io_out_a_0(_mesh_0_13_io_out_a_0),
		.io_out_c_0(_mesh_0_13_io_out_c_0),
		.io_out_b_0(_mesh_0_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_13_io_out_id_0),
		.io_out_last_0(_mesh_0_13_io_out_last_0),
		.io_out_valid_0(_mesh_0_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9384 == GlobalFiModInstNr[0]) || (9384 == GlobalFiModInstNr[1]) || (9384 == GlobalFiModInstNr[2]) || (9384 == GlobalFiModInstNr[3]))));
	Tile mesh_0_14(
		.clock(clock),
		.io_in_a_0(r_14_0),
		.io_in_b_0(b_448_0),
		.io_in_d_0(b_1472_0),
		.io_in_control_0_dataflow(mesh_0_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2496_0),
		.io_in_last_0(r_3520_0),
		.io_in_valid_0(r_1472_0),
		.io_out_a_0(_mesh_0_14_io_out_a_0),
		.io_out_c_0(_mesh_0_14_io_out_c_0),
		.io_out_b_0(_mesh_0_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_14_io_out_id_0),
		.io_out_last_0(_mesh_0_14_io_out_last_0),
		.io_out_valid_0(_mesh_0_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9385 == GlobalFiModInstNr[0]) || (9385 == GlobalFiModInstNr[1]) || (9385 == GlobalFiModInstNr[2]) || (9385 == GlobalFiModInstNr[3]))));
	Tile mesh_0_15(
		.clock(clock),
		.io_in_a_0(r_15_0),
		.io_in_b_0(b_480_0),
		.io_in_d_0(b_1504_0),
		.io_in_control_0_dataflow(mesh_0_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2528_0),
		.io_in_last_0(r_3552_0),
		.io_in_valid_0(r_1504_0),
		.io_out_a_0(_mesh_0_15_io_out_a_0),
		.io_out_c_0(_mesh_0_15_io_out_c_0),
		.io_out_b_0(_mesh_0_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_15_io_out_id_0),
		.io_out_last_0(_mesh_0_15_io_out_last_0),
		.io_out_valid_0(_mesh_0_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9386 == GlobalFiModInstNr[0]) || (9386 == GlobalFiModInstNr[1]) || (9386 == GlobalFiModInstNr[2]) || (9386 == GlobalFiModInstNr[3]))));
	Tile mesh_0_16(
		.clock(clock),
		.io_in_a_0(r_16_0),
		.io_in_b_0(b_512_0),
		.io_in_d_0(b_1536_0),
		.io_in_control_0_dataflow(mesh_0_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2560_0),
		.io_in_last_0(r_3584_0),
		.io_in_valid_0(r_1536_0),
		.io_out_a_0(_mesh_0_16_io_out_a_0),
		.io_out_c_0(_mesh_0_16_io_out_c_0),
		.io_out_b_0(_mesh_0_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_16_io_out_id_0),
		.io_out_last_0(_mesh_0_16_io_out_last_0),
		.io_out_valid_0(_mesh_0_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9387 == GlobalFiModInstNr[0]) || (9387 == GlobalFiModInstNr[1]) || (9387 == GlobalFiModInstNr[2]) || (9387 == GlobalFiModInstNr[3]))));
	Tile mesh_0_17(
		.clock(clock),
		.io_in_a_0(r_17_0),
		.io_in_b_0(b_544_0),
		.io_in_d_0(b_1568_0),
		.io_in_control_0_dataflow(mesh_0_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2592_0),
		.io_in_last_0(r_3616_0),
		.io_in_valid_0(r_1568_0),
		.io_out_a_0(_mesh_0_17_io_out_a_0),
		.io_out_c_0(_mesh_0_17_io_out_c_0),
		.io_out_b_0(_mesh_0_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_17_io_out_id_0),
		.io_out_last_0(_mesh_0_17_io_out_last_0),
		.io_out_valid_0(_mesh_0_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9388 == GlobalFiModInstNr[0]) || (9388 == GlobalFiModInstNr[1]) || (9388 == GlobalFiModInstNr[2]) || (9388 == GlobalFiModInstNr[3]))));
	Tile mesh_0_18(
		.clock(clock),
		.io_in_a_0(r_18_0),
		.io_in_b_0(b_576_0),
		.io_in_d_0(b_1600_0),
		.io_in_control_0_dataflow(mesh_0_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2624_0),
		.io_in_last_0(r_3648_0),
		.io_in_valid_0(r_1600_0),
		.io_out_a_0(_mesh_0_18_io_out_a_0),
		.io_out_c_0(_mesh_0_18_io_out_c_0),
		.io_out_b_0(_mesh_0_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_18_io_out_id_0),
		.io_out_last_0(_mesh_0_18_io_out_last_0),
		.io_out_valid_0(_mesh_0_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9389 == GlobalFiModInstNr[0]) || (9389 == GlobalFiModInstNr[1]) || (9389 == GlobalFiModInstNr[2]) || (9389 == GlobalFiModInstNr[3]))));
	Tile mesh_0_19(
		.clock(clock),
		.io_in_a_0(r_19_0),
		.io_in_b_0(b_608_0),
		.io_in_d_0(b_1632_0),
		.io_in_control_0_dataflow(mesh_0_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2656_0),
		.io_in_last_0(r_3680_0),
		.io_in_valid_0(r_1632_0),
		.io_out_a_0(_mesh_0_19_io_out_a_0),
		.io_out_c_0(_mesh_0_19_io_out_c_0),
		.io_out_b_0(_mesh_0_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_19_io_out_id_0),
		.io_out_last_0(_mesh_0_19_io_out_last_0),
		.io_out_valid_0(_mesh_0_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9390 == GlobalFiModInstNr[0]) || (9390 == GlobalFiModInstNr[1]) || (9390 == GlobalFiModInstNr[2]) || (9390 == GlobalFiModInstNr[3]))));
	Tile mesh_0_20(
		.clock(clock),
		.io_in_a_0(r_20_0),
		.io_in_b_0(b_640_0),
		.io_in_d_0(b_1664_0),
		.io_in_control_0_dataflow(mesh_0_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2688_0),
		.io_in_last_0(r_3712_0),
		.io_in_valid_0(r_1664_0),
		.io_out_a_0(_mesh_0_20_io_out_a_0),
		.io_out_c_0(_mesh_0_20_io_out_c_0),
		.io_out_b_0(_mesh_0_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_20_io_out_id_0),
		.io_out_last_0(_mesh_0_20_io_out_last_0),
		.io_out_valid_0(_mesh_0_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9391 == GlobalFiModInstNr[0]) || (9391 == GlobalFiModInstNr[1]) || (9391 == GlobalFiModInstNr[2]) || (9391 == GlobalFiModInstNr[3]))));
	Tile mesh_0_21(
		.clock(clock),
		.io_in_a_0(r_21_0),
		.io_in_b_0(b_672_0),
		.io_in_d_0(b_1696_0),
		.io_in_control_0_dataflow(mesh_0_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2720_0),
		.io_in_last_0(r_3744_0),
		.io_in_valid_0(r_1696_0),
		.io_out_a_0(_mesh_0_21_io_out_a_0),
		.io_out_c_0(_mesh_0_21_io_out_c_0),
		.io_out_b_0(_mesh_0_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_21_io_out_id_0),
		.io_out_last_0(_mesh_0_21_io_out_last_0),
		.io_out_valid_0(_mesh_0_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9392 == GlobalFiModInstNr[0]) || (9392 == GlobalFiModInstNr[1]) || (9392 == GlobalFiModInstNr[2]) || (9392 == GlobalFiModInstNr[3]))));
	Tile mesh_0_22(
		.clock(clock),
		.io_in_a_0(r_22_0),
		.io_in_b_0(b_704_0),
		.io_in_d_0(b_1728_0),
		.io_in_control_0_dataflow(mesh_0_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2752_0),
		.io_in_last_0(r_3776_0),
		.io_in_valid_0(r_1728_0),
		.io_out_a_0(_mesh_0_22_io_out_a_0),
		.io_out_c_0(_mesh_0_22_io_out_c_0),
		.io_out_b_0(_mesh_0_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_22_io_out_id_0),
		.io_out_last_0(_mesh_0_22_io_out_last_0),
		.io_out_valid_0(_mesh_0_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9393 == GlobalFiModInstNr[0]) || (9393 == GlobalFiModInstNr[1]) || (9393 == GlobalFiModInstNr[2]) || (9393 == GlobalFiModInstNr[3]))));
	Tile mesh_0_23(
		.clock(clock),
		.io_in_a_0(r_23_0),
		.io_in_b_0(b_736_0),
		.io_in_d_0(b_1760_0),
		.io_in_control_0_dataflow(mesh_0_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2784_0),
		.io_in_last_0(r_3808_0),
		.io_in_valid_0(r_1760_0),
		.io_out_a_0(_mesh_0_23_io_out_a_0),
		.io_out_c_0(_mesh_0_23_io_out_c_0),
		.io_out_b_0(_mesh_0_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_23_io_out_id_0),
		.io_out_last_0(_mesh_0_23_io_out_last_0),
		.io_out_valid_0(_mesh_0_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9394 == GlobalFiModInstNr[0]) || (9394 == GlobalFiModInstNr[1]) || (9394 == GlobalFiModInstNr[2]) || (9394 == GlobalFiModInstNr[3]))));
	Tile mesh_0_24(
		.clock(clock),
		.io_in_a_0(r_24_0),
		.io_in_b_0(b_768_0),
		.io_in_d_0(b_1792_0),
		.io_in_control_0_dataflow(mesh_0_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2816_0),
		.io_in_last_0(r_3840_0),
		.io_in_valid_0(r_1792_0),
		.io_out_a_0(_mesh_0_24_io_out_a_0),
		.io_out_c_0(_mesh_0_24_io_out_c_0),
		.io_out_b_0(_mesh_0_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_24_io_out_id_0),
		.io_out_last_0(_mesh_0_24_io_out_last_0),
		.io_out_valid_0(_mesh_0_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9395 == GlobalFiModInstNr[0]) || (9395 == GlobalFiModInstNr[1]) || (9395 == GlobalFiModInstNr[2]) || (9395 == GlobalFiModInstNr[3]))));
	Tile mesh_0_25(
		.clock(clock),
		.io_in_a_0(r_25_0),
		.io_in_b_0(b_800_0),
		.io_in_d_0(b_1824_0),
		.io_in_control_0_dataflow(mesh_0_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2848_0),
		.io_in_last_0(r_3872_0),
		.io_in_valid_0(r_1824_0),
		.io_out_a_0(_mesh_0_25_io_out_a_0),
		.io_out_c_0(_mesh_0_25_io_out_c_0),
		.io_out_b_0(_mesh_0_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_25_io_out_id_0),
		.io_out_last_0(_mesh_0_25_io_out_last_0),
		.io_out_valid_0(_mesh_0_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9396 == GlobalFiModInstNr[0]) || (9396 == GlobalFiModInstNr[1]) || (9396 == GlobalFiModInstNr[2]) || (9396 == GlobalFiModInstNr[3]))));
	Tile mesh_0_26(
		.clock(clock),
		.io_in_a_0(r_26_0),
		.io_in_b_0(b_832_0),
		.io_in_d_0(b_1856_0),
		.io_in_control_0_dataflow(mesh_0_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2880_0),
		.io_in_last_0(r_3904_0),
		.io_in_valid_0(r_1856_0),
		.io_out_a_0(_mesh_0_26_io_out_a_0),
		.io_out_c_0(_mesh_0_26_io_out_c_0),
		.io_out_b_0(_mesh_0_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_26_io_out_id_0),
		.io_out_last_0(_mesh_0_26_io_out_last_0),
		.io_out_valid_0(_mesh_0_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9397 == GlobalFiModInstNr[0]) || (9397 == GlobalFiModInstNr[1]) || (9397 == GlobalFiModInstNr[2]) || (9397 == GlobalFiModInstNr[3]))));
	Tile mesh_0_27(
		.clock(clock),
		.io_in_a_0(r_27_0),
		.io_in_b_0(b_864_0),
		.io_in_d_0(b_1888_0),
		.io_in_control_0_dataflow(mesh_0_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2912_0),
		.io_in_last_0(r_3936_0),
		.io_in_valid_0(r_1888_0),
		.io_out_a_0(_mesh_0_27_io_out_a_0),
		.io_out_c_0(_mesh_0_27_io_out_c_0),
		.io_out_b_0(_mesh_0_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_27_io_out_id_0),
		.io_out_last_0(_mesh_0_27_io_out_last_0),
		.io_out_valid_0(_mesh_0_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9398 == GlobalFiModInstNr[0]) || (9398 == GlobalFiModInstNr[1]) || (9398 == GlobalFiModInstNr[2]) || (9398 == GlobalFiModInstNr[3]))));
	Tile mesh_0_28(
		.clock(clock),
		.io_in_a_0(r_28_0),
		.io_in_b_0(b_896_0),
		.io_in_d_0(b_1920_0),
		.io_in_control_0_dataflow(mesh_0_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2944_0),
		.io_in_last_0(r_3968_0),
		.io_in_valid_0(r_1920_0),
		.io_out_a_0(_mesh_0_28_io_out_a_0),
		.io_out_c_0(_mesh_0_28_io_out_c_0),
		.io_out_b_0(_mesh_0_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_28_io_out_id_0),
		.io_out_last_0(_mesh_0_28_io_out_last_0),
		.io_out_valid_0(_mesh_0_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9399 == GlobalFiModInstNr[0]) || (9399 == GlobalFiModInstNr[1]) || (9399 == GlobalFiModInstNr[2]) || (9399 == GlobalFiModInstNr[3]))));
	Tile mesh_0_29(
		.clock(clock),
		.io_in_a_0(r_29_0),
		.io_in_b_0(b_928_0),
		.io_in_d_0(b_1952_0),
		.io_in_control_0_dataflow(mesh_0_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2976_0),
		.io_in_last_0(r_4000_0),
		.io_in_valid_0(r_1952_0),
		.io_out_a_0(_mesh_0_29_io_out_a_0),
		.io_out_c_0(_mesh_0_29_io_out_c_0),
		.io_out_b_0(_mesh_0_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_29_io_out_id_0),
		.io_out_last_0(_mesh_0_29_io_out_last_0),
		.io_out_valid_0(_mesh_0_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9400 == GlobalFiModInstNr[0]) || (9400 == GlobalFiModInstNr[1]) || (9400 == GlobalFiModInstNr[2]) || (9400 == GlobalFiModInstNr[3]))));
	Tile mesh_0_30(
		.clock(clock),
		.io_in_a_0(r_30_0),
		.io_in_b_0(b_960_0),
		.io_in_d_0(b_1984_0),
		.io_in_control_0_dataflow(mesh_0_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3008_0),
		.io_in_last_0(r_4032_0),
		.io_in_valid_0(r_1984_0),
		.io_out_a_0(_mesh_0_30_io_out_a_0),
		.io_out_c_0(_mesh_0_30_io_out_c_0),
		.io_out_b_0(_mesh_0_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_30_io_out_id_0),
		.io_out_last_0(_mesh_0_30_io_out_last_0),
		.io_out_valid_0(_mesh_0_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9401 == GlobalFiModInstNr[0]) || (9401 == GlobalFiModInstNr[1]) || (9401 == GlobalFiModInstNr[2]) || (9401 == GlobalFiModInstNr[3]))));
	Tile mesh_0_31(
		.clock(clock),
		.io_in_a_0(r_31_0),
		.io_in_b_0(b_992_0),
		.io_in_d_0(b_2016_0),
		.io_in_control_0_dataflow(mesh_0_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3040_0),
		.io_in_last_0(r_4064_0),
		.io_in_valid_0(r_2016_0),
		.io_out_a_0(_mesh_0_31_io_out_a_0),
		.io_out_c_0(_mesh_0_31_io_out_c_0),
		.io_out_b_0(_mesh_0_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_31_io_out_id_0),
		.io_out_last_0(_mesh_0_31_io_out_last_0),
		.io_out_valid_0(_mesh_0_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9402 == GlobalFiModInstNr[0]) || (9402 == GlobalFiModInstNr[1]) || (9402 == GlobalFiModInstNr[2]) || (9402 == GlobalFiModInstNr[3]))));
	Tile mesh_1_0(
		.clock(clock),
		.io_in_a_0(r_32_0),
		.io_in_b_0(b_1_0),
		.io_in_d_0(b_1025_0),
		.io_in_control_0_dataflow(mesh_1_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2049_0),
		.io_in_last_0(r_3073_0),
		.io_in_valid_0(r_1025_0),
		.io_out_a_0(_mesh_1_0_io_out_a_0),
		.io_out_c_0(_mesh_1_0_io_out_c_0),
		.io_out_b_0(_mesh_1_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_0_io_out_id_0),
		.io_out_last_0(_mesh_1_0_io_out_last_0),
		.io_out_valid_0(_mesh_1_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9403 == GlobalFiModInstNr[0]) || (9403 == GlobalFiModInstNr[1]) || (9403 == GlobalFiModInstNr[2]) || (9403 == GlobalFiModInstNr[3]))));
	Tile mesh_1_1(
		.clock(clock),
		.io_in_a_0(r_33_0),
		.io_in_b_0(b_33_0),
		.io_in_d_0(b_1057_0),
		.io_in_control_0_dataflow(mesh_1_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2081_0),
		.io_in_last_0(r_3105_0),
		.io_in_valid_0(r_1057_0),
		.io_out_a_0(_mesh_1_1_io_out_a_0),
		.io_out_c_0(_mesh_1_1_io_out_c_0),
		.io_out_b_0(_mesh_1_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_1_io_out_id_0),
		.io_out_last_0(_mesh_1_1_io_out_last_0),
		.io_out_valid_0(_mesh_1_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9404 == GlobalFiModInstNr[0]) || (9404 == GlobalFiModInstNr[1]) || (9404 == GlobalFiModInstNr[2]) || (9404 == GlobalFiModInstNr[3]))));
	Tile mesh_1_2(
		.clock(clock),
		.io_in_a_0(r_34_0),
		.io_in_b_0(b_65_0),
		.io_in_d_0(b_1089_0),
		.io_in_control_0_dataflow(mesh_1_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2113_0),
		.io_in_last_0(r_3137_0),
		.io_in_valid_0(r_1089_0),
		.io_out_a_0(_mesh_1_2_io_out_a_0),
		.io_out_c_0(_mesh_1_2_io_out_c_0),
		.io_out_b_0(_mesh_1_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_2_io_out_id_0),
		.io_out_last_0(_mesh_1_2_io_out_last_0),
		.io_out_valid_0(_mesh_1_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9405 == GlobalFiModInstNr[0]) || (9405 == GlobalFiModInstNr[1]) || (9405 == GlobalFiModInstNr[2]) || (9405 == GlobalFiModInstNr[3]))));
	Tile mesh_1_3(
		.clock(clock),
		.io_in_a_0(r_35_0),
		.io_in_b_0(b_97_0),
		.io_in_d_0(b_1121_0),
		.io_in_control_0_dataflow(mesh_1_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2145_0),
		.io_in_last_0(r_3169_0),
		.io_in_valid_0(r_1121_0),
		.io_out_a_0(_mesh_1_3_io_out_a_0),
		.io_out_c_0(_mesh_1_3_io_out_c_0),
		.io_out_b_0(_mesh_1_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_3_io_out_id_0),
		.io_out_last_0(_mesh_1_3_io_out_last_0),
		.io_out_valid_0(_mesh_1_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9406 == GlobalFiModInstNr[0]) || (9406 == GlobalFiModInstNr[1]) || (9406 == GlobalFiModInstNr[2]) || (9406 == GlobalFiModInstNr[3]))));
	Tile mesh_1_4(
		.clock(clock),
		.io_in_a_0(r_36_0),
		.io_in_b_0(b_129_0),
		.io_in_d_0(b_1153_0),
		.io_in_control_0_dataflow(mesh_1_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2177_0),
		.io_in_last_0(r_3201_0),
		.io_in_valid_0(r_1153_0),
		.io_out_a_0(_mesh_1_4_io_out_a_0),
		.io_out_c_0(_mesh_1_4_io_out_c_0),
		.io_out_b_0(_mesh_1_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_4_io_out_id_0),
		.io_out_last_0(_mesh_1_4_io_out_last_0),
		.io_out_valid_0(_mesh_1_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9407 == GlobalFiModInstNr[0]) || (9407 == GlobalFiModInstNr[1]) || (9407 == GlobalFiModInstNr[2]) || (9407 == GlobalFiModInstNr[3]))));
	Tile mesh_1_5(
		.clock(clock),
		.io_in_a_0(r_37_0),
		.io_in_b_0(b_161_0),
		.io_in_d_0(b_1185_0),
		.io_in_control_0_dataflow(mesh_1_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2209_0),
		.io_in_last_0(r_3233_0),
		.io_in_valid_0(r_1185_0),
		.io_out_a_0(_mesh_1_5_io_out_a_0),
		.io_out_c_0(_mesh_1_5_io_out_c_0),
		.io_out_b_0(_mesh_1_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_5_io_out_id_0),
		.io_out_last_0(_mesh_1_5_io_out_last_0),
		.io_out_valid_0(_mesh_1_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9408 == GlobalFiModInstNr[0]) || (9408 == GlobalFiModInstNr[1]) || (9408 == GlobalFiModInstNr[2]) || (9408 == GlobalFiModInstNr[3]))));
	Tile mesh_1_6(
		.clock(clock),
		.io_in_a_0(r_38_0),
		.io_in_b_0(b_193_0),
		.io_in_d_0(b_1217_0),
		.io_in_control_0_dataflow(mesh_1_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2241_0),
		.io_in_last_0(r_3265_0),
		.io_in_valid_0(r_1217_0),
		.io_out_a_0(_mesh_1_6_io_out_a_0),
		.io_out_c_0(_mesh_1_6_io_out_c_0),
		.io_out_b_0(_mesh_1_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_6_io_out_id_0),
		.io_out_last_0(_mesh_1_6_io_out_last_0),
		.io_out_valid_0(_mesh_1_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9409 == GlobalFiModInstNr[0]) || (9409 == GlobalFiModInstNr[1]) || (9409 == GlobalFiModInstNr[2]) || (9409 == GlobalFiModInstNr[3]))));
	Tile mesh_1_7(
		.clock(clock),
		.io_in_a_0(r_39_0),
		.io_in_b_0(b_225_0),
		.io_in_d_0(b_1249_0),
		.io_in_control_0_dataflow(mesh_1_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2273_0),
		.io_in_last_0(r_3297_0),
		.io_in_valid_0(r_1249_0),
		.io_out_a_0(_mesh_1_7_io_out_a_0),
		.io_out_c_0(_mesh_1_7_io_out_c_0),
		.io_out_b_0(_mesh_1_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_7_io_out_id_0),
		.io_out_last_0(_mesh_1_7_io_out_last_0),
		.io_out_valid_0(_mesh_1_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9410 == GlobalFiModInstNr[0]) || (9410 == GlobalFiModInstNr[1]) || (9410 == GlobalFiModInstNr[2]) || (9410 == GlobalFiModInstNr[3]))));
	Tile mesh_1_8(
		.clock(clock),
		.io_in_a_0(r_40_0),
		.io_in_b_0(b_257_0),
		.io_in_d_0(b_1281_0),
		.io_in_control_0_dataflow(mesh_1_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2305_0),
		.io_in_last_0(r_3329_0),
		.io_in_valid_0(r_1281_0),
		.io_out_a_0(_mesh_1_8_io_out_a_0),
		.io_out_c_0(_mesh_1_8_io_out_c_0),
		.io_out_b_0(_mesh_1_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_8_io_out_id_0),
		.io_out_last_0(_mesh_1_8_io_out_last_0),
		.io_out_valid_0(_mesh_1_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9411 == GlobalFiModInstNr[0]) || (9411 == GlobalFiModInstNr[1]) || (9411 == GlobalFiModInstNr[2]) || (9411 == GlobalFiModInstNr[3]))));
	Tile mesh_1_9(
		.clock(clock),
		.io_in_a_0(r_41_0),
		.io_in_b_0(b_289_0),
		.io_in_d_0(b_1313_0),
		.io_in_control_0_dataflow(mesh_1_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2337_0),
		.io_in_last_0(r_3361_0),
		.io_in_valid_0(r_1313_0),
		.io_out_a_0(_mesh_1_9_io_out_a_0),
		.io_out_c_0(_mesh_1_9_io_out_c_0),
		.io_out_b_0(_mesh_1_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_9_io_out_id_0),
		.io_out_last_0(_mesh_1_9_io_out_last_0),
		.io_out_valid_0(_mesh_1_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9412 == GlobalFiModInstNr[0]) || (9412 == GlobalFiModInstNr[1]) || (9412 == GlobalFiModInstNr[2]) || (9412 == GlobalFiModInstNr[3]))));
	Tile mesh_1_10(
		.clock(clock),
		.io_in_a_0(r_42_0),
		.io_in_b_0(b_321_0),
		.io_in_d_0(b_1345_0),
		.io_in_control_0_dataflow(mesh_1_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2369_0),
		.io_in_last_0(r_3393_0),
		.io_in_valid_0(r_1345_0),
		.io_out_a_0(_mesh_1_10_io_out_a_0),
		.io_out_c_0(_mesh_1_10_io_out_c_0),
		.io_out_b_0(_mesh_1_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_10_io_out_id_0),
		.io_out_last_0(_mesh_1_10_io_out_last_0),
		.io_out_valid_0(_mesh_1_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9413 == GlobalFiModInstNr[0]) || (9413 == GlobalFiModInstNr[1]) || (9413 == GlobalFiModInstNr[2]) || (9413 == GlobalFiModInstNr[3]))));
	Tile mesh_1_11(
		.clock(clock),
		.io_in_a_0(r_43_0),
		.io_in_b_0(b_353_0),
		.io_in_d_0(b_1377_0),
		.io_in_control_0_dataflow(mesh_1_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2401_0),
		.io_in_last_0(r_3425_0),
		.io_in_valid_0(r_1377_0),
		.io_out_a_0(_mesh_1_11_io_out_a_0),
		.io_out_c_0(_mesh_1_11_io_out_c_0),
		.io_out_b_0(_mesh_1_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_11_io_out_id_0),
		.io_out_last_0(_mesh_1_11_io_out_last_0),
		.io_out_valid_0(_mesh_1_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9414 == GlobalFiModInstNr[0]) || (9414 == GlobalFiModInstNr[1]) || (9414 == GlobalFiModInstNr[2]) || (9414 == GlobalFiModInstNr[3]))));
	Tile mesh_1_12(
		.clock(clock),
		.io_in_a_0(r_44_0),
		.io_in_b_0(b_385_0),
		.io_in_d_0(b_1409_0),
		.io_in_control_0_dataflow(mesh_1_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2433_0),
		.io_in_last_0(r_3457_0),
		.io_in_valid_0(r_1409_0),
		.io_out_a_0(_mesh_1_12_io_out_a_0),
		.io_out_c_0(_mesh_1_12_io_out_c_0),
		.io_out_b_0(_mesh_1_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_12_io_out_id_0),
		.io_out_last_0(_mesh_1_12_io_out_last_0),
		.io_out_valid_0(_mesh_1_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9415 == GlobalFiModInstNr[0]) || (9415 == GlobalFiModInstNr[1]) || (9415 == GlobalFiModInstNr[2]) || (9415 == GlobalFiModInstNr[3]))));
	Tile mesh_1_13(
		.clock(clock),
		.io_in_a_0(r_45_0),
		.io_in_b_0(b_417_0),
		.io_in_d_0(b_1441_0),
		.io_in_control_0_dataflow(mesh_1_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2465_0),
		.io_in_last_0(r_3489_0),
		.io_in_valid_0(r_1441_0),
		.io_out_a_0(_mesh_1_13_io_out_a_0),
		.io_out_c_0(_mesh_1_13_io_out_c_0),
		.io_out_b_0(_mesh_1_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_13_io_out_id_0),
		.io_out_last_0(_mesh_1_13_io_out_last_0),
		.io_out_valid_0(_mesh_1_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9416 == GlobalFiModInstNr[0]) || (9416 == GlobalFiModInstNr[1]) || (9416 == GlobalFiModInstNr[2]) || (9416 == GlobalFiModInstNr[3]))));
	Tile mesh_1_14(
		.clock(clock),
		.io_in_a_0(r_46_0),
		.io_in_b_0(b_449_0),
		.io_in_d_0(b_1473_0),
		.io_in_control_0_dataflow(mesh_1_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2497_0),
		.io_in_last_0(r_3521_0),
		.io_in_valid_0(r_1473_0),
		.io_out_a_0(_mesh_1_14_io_out_a_0),
		.io_out_c_0(_mesh_1_14_io_out_c_0),
		.io_out_b_0(_mesh_1_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_14_io_out_id_0),
		.io_out_last_0(_mesh_1_14_io_out_last_0),
		.io_out_valid_0(_mesh_1_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9417 == GlobalFiModInstNr[0]) || (9417 == GlobalFiModInstNr[1]) || (9417 == GlobalFiModInstNr[2]) || (9417 == GlobalFiModInstNr[3]))));
	Tile mesh_1_15(
		.clock(clock),
		.io_in_a_0(r_47_0),
		.io_in_b_0(b_481_0),
		.io_in_d_0(b_1505_0),
		.io_in_control_0_dataflow(mesh_1_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2529_0),
		.io_in_last_0(r_3553_0),
		.io_in_valid_0(r_1505_0),
		.io_out_a_0(_mesh_1_15_io_out_a_0),
		.io_out_c_0(_mesh_1_15_io_out_c_0),
		.io_out_b_0(_mesh_1_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_15_io_out_id_0),
		.io_out_last_0(_mesh_1_15_io_out_last_0),
		.io_out_valid_0(_mesh_1_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9418 == GlobalFiModInstNr[0]) || (9418 == GlobalFiModInstNr[1]) || (9418 == GlobalFiModInstNr[2]) || (9418 == GlobalFiModInstNr[3]))));
	Tile mesh_1_16(
		.clock(clock),
		.io_in_a_0(r_48_0),
		.io_in_b_0(b_513_0),
		.io_in_d_0(b_1537_0),
		.io_in_control_0_dataflow(mesh_1_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2561_0),
		.io_in_last_0(r_3585_0),
		.io_in_valid_0(r_1537_0),
		.io_out_a_0(_mesh_1_16_io_out_a_0),
		.io_out_c_0(_mesh_1_16_io_out_c_0),
		.io_out_b_0(_mesh_1_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_16_io_out_id_0),
		.io_out_last_0(_mesh_1_16_io_out_last_0),
		.io_out_valid_0(_mesh_1_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9419 == GlobalFiModInstNr[0]) || (9419 == GlobalFiModInstNr[1]) || (9419 == GlobalFiModInstNr[2]) || (9419 == GlobalFiModInstNr[3]))));
	Tile mesh_1_17(
		.clock(clock),
		.io_in_a_0(r_49_0),
		.io_in_b_0(b_545_0),
		.io_in_d_0(b_1569_0),
		.io_in_control_0_dataflow(mesh_1_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2593_0),
		.io_in_last_0(r_3617_0),
		.io_in_valid_0(r_1569_0),
		.io_out_a_0(_mesh_1_17_io_out_a_0),
		.io_out_c_0(_mesh_1_17_io_out_c_0),
		.io_out_b_0(_mesh_1_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_17_io_out_id_0),
		.io_out_last_0(_mesh_1_17_io_out_last_0),
		.io_out_valid_0(_mesh_1_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9420 == GlobalFiModInstNr[0]) || (9420 == GlobalFiModInstNr[1]) || (9420 == GlobalFiModInstNr[2]) || (9420 == GlobalFiModInstNr[3]))));
	Tile mesh_1_18(
		.clock(clock),
		.io_in_a_0(r_50_0),
		.io_in_b_0(b_577_0),
		.io_in_d_0(b_1601_0),
		.io_in_control_0_dataflow(mesh_1_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2625_0),
		.io_in_last_0(r_3649_0),
		.io_in_valid_0(r_1601_0),
		.io_out_a_0(_mesh_1_18_io_out_a_0),
		.io_out_c_0(_mesh_1_18_io_out_c_0),
		.io_out_b_0(_mesh_1_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_18_io_out_id_0),
		.io_out_last_0(_mesh_1_18_io_out_last_0),
		.io_out_valid_0(_mesh_1_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9421 == GlobalFiModInstNr[0]) || (9421 == GlobalFiModInstNr[1]) || (9421 == GlobalFiModInstNr[2]) || (9421 == GlobalFiModInstNr[3]))));
	Tile mesh_1_19(
		.clock(clock),
		.io_in_a_0(r_51_0),
		.io_in_b_0(b_609_0),
		.io_in_d_0(b_1633_0),
		.io_in_control_0_dataflow(mesh_1_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2657_0),
		.io_in_last_0(r_3681_0),
		.io_in_valid_0(r_1633_0),
		.io_out_a_0(_mesh_1_19_io_out_a_0),
		.io_out_c_0(_mesh_1_19_io_out_c_0),
		.io_out_b_0(_mesh_1_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_19_io_out_id_0),
		.io_out_last_0(_mesh_1_19_io_out_last_0),
		.io_out_valid_0(_mesh_1_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9422 == GlobalFiModInstNr[0]) || (9422 == GlobalFiModInstNr[1]) || (9422 == GlobalFiModInstNr[2]) || (9422 == GlobalFiModInstNr[3]))));
	Tile mesh_1_20(
		.clock(clock),
		.io_in_a_0(r_52_0),
		.io_in_b_0(b_641_0),
		.io_in_d_0(b_1665_0),
		.io_in_control_0_dataflow(mesh_1_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2689_0),
		.io_in_last_0(r_3713_0),
		.io_in_valid_0(r_1665_0),
		.io_out_a_0(_mesh_1_20_io_out_a_0),
		.io_out_c_0(_mesh_1_20_io_out_c_0),
		.io_out_b_0(_mesh_1_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_20_io_out_id_0),
		.io_out_last_0(_mesh_1_20_io_out_last_0),
		.io_out_valid_0(_mesh_1_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9423 == GlobalFiModInstNr[0]) || (9423 == GlobalFiModInstNr[1]) || (9423 == GlobalFiModInstNr[2]) || (9423 == GlobalFiModInstNr[3]))));
	Tile mesh_1_21(
		.clock(clock),
		.io_in_a_0(r_53_0),
		.io_in_b_0(b_673_0),
		.io_in_d_0(b_1697_0),
		.io_in_control_0_dataflow(mesh_1_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2721_0),
		.io_in_last_0(r_3745_0),
		.io_in_valid_0(r_1697_0),
		.io_out_a_0(_mesh_1_21_io_out_a_0),
		.io_out_c_0(_mesh_1_21_io_out_c_0),
		.io_out_b_0(_mesh_1_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_21_io_out_id_0),
		.io_out_last_0(_mesh_1_21_io_out_last_0),
		.io_out_valid_0(_mesh_1_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9424 == GlobalFiModInstNr[0]) || (9424 == GlobalFiModInstNr[1]) || (9424 == GlobalFiModInstNr[2]) || (9424 == GlobalFiModInstNr[3]))));
	Tile mesh_1_22(
		.clock(clock),
		.io_in_a_0(r_54_0),
		.io_in_b_0(b_705_0),
		.io_in_d_0(b_1729_0),
		.io_in_control_0_dataflow(mesh_1_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2753_0),
		.io_in_last_0(r_3777_0),
		.io_in_valid_0(r_1729_0),
		.io_out_a_0(_mesh_1_22_io_out_a_0),
		.io_out_c_0(_mesh_1_22_io_out_c_0),
		.io_out_b_0(_mesh_1_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_22_io_out_id_0),
		.io_out_last_0(_mesh_1_22_io_out_last_0),
		.io_out_valid_0(_mesh_1_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9425 == GlobalFiModInstNr[0]) || (9425 == GlobalFiModInstNr[1]) || (9425 == GlobalFiModInstNr[2]) || (9425 == GlobalFiModInstNr[3]))));
	Tile mesh_1_23(
		.clock(clock),
		.io_in_a_0(r_55_0),
		.io_in_b_0(b_737_0),
		.io_in_d_0(b_1761_0),
		.io_in_control_0_dataflow(mesh_1_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2785_0),
		.io_in_last_0(r_3809_0),
		.io_in_valid_0(r_1761_0),
		.io_out_a_0(_mesh_1_23_io_out_a_0),
		.io_out_c_0(_mesh_1_23_io_out_c_0),
		.io_out_b_0(_mesh_1_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_23_io_out_id_0),
		.io_out_last_0(_mesh_1_23_io_out_last_0),
		.io_out_valid_0(_mesh_1_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9426 == GlobalFiModInstNr[0]) || (9426 == GlobalFiModInstNr[1]) || (9426 == GlobalFiModInstNr[2]) || (9426 == GlobalFiModInstNr[3]))));
	Tile mesh_1_24(
		.clock(clock),
		.io_in_a_0(r_56_0),
		.io_in_b_0(b_769_0),
		.io_in_d_0(b_1793_0),
		.io_in_control_0_dataflow(mesh_1_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2817_0),
		.io_in_last_0(r_3841_0),
		.io_in_valid_0(r_1793_0),
		.io_out_a_0(_mesh_1_24_io_out_a_0),
		.io_out_c_0(_mesh_1_24_io_out_c_0),
		.io_out_b_0(_mesh_1_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_24_io_out_id_0),
		.io_out_last_0(_mesh_1_24_io_out_last_0),
		.io_out_valid_0(_mesh_1_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9427 == GlobalFiModInstNr[0]) || (9427 == GlobalFiModInstNr[1]) || (9427 == GlobalFiModInstNr[2]) || (9427 == GlobalFiModInstNr[3]))));
	Tile mesh_1_25(
		.clock(clock),
		.io_in_a_0(r_57_0),
		.io_in_b_0(b_801_0),
		.io_in_d_0(b_1825_0),
		.io_in_control_0_dataflow(mesh_1_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2849_0),
		.io_in_last_0(r_3873_0),
		.io_in_valid_0(r_1825_0),
		.io_out_a_0(_mesh_1_25_io_out_a_0),
		.io_out_c_0(_mesh_1_25_io_out_c_0),
		.io_out_b_0(_mesh_1_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_25_io_out_id_0),
		.io_out_last_0(_mesh_1_25_io_out_last_0),
		.io_out_valid_0(_mesh_1_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9428 == GlobalFiModInstNr[0]) || (9428 == GlobalFiModInstNr[1]) || (9428 == GlobalFiModInstNr[2]) || (9428 == GlobalFiModInstNr[3]))));
	Tile mesh_1_26(
		.clock(clock),
		.io_in_a_0(r_58_0),
		.io_in_b_0(b_833_0),
		.io_in_d_0(b_1857_0),
		.io_in_control_0_dataflow(mesh_1_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2881_0),
		.io_in_last_0(r_3905_0),
		.io_in_valid_0(r_1857_0),
		.io_out_a_0(_mesh_1_26_io_out_a_0),
		.io_out_c_0(_mesh_1_26_io_out_c_0),
		.io_out_b_0(_mesh_1_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_26_io_out_id_0),
		.io_out_last_0(_mesh_1_26_io_out_last_0),
		.io_out_valid_0(_mesh_1_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9429 == GlobalFiModInstNr[0]) || (9429 == GlobalFiModInstNr[1]) || (9429 == GlobalFiModInstNr[2]) || (9429 == GlobalFiModInstNr[3]))));
	Tile mesh_1_27(
		.clock(clock),
		.io_in_a_0(r_59_0),
		.io_in_b_0(b_865_0),
		.io_in_d_0(b_1889_0),
		.io_in_control_0_dataflow(mesh_1_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2913_0),
		.io_in_last_0(r_3937_0),
		.io_in_valid_0(r_1889_0),
		.io_out_a_0(_mesh_1_27_io_out_a_0),
		.io_out_c_0(_mesh_1_27_io_out_c_0),
		.io_out_b_0(_mesh_1_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_27_io_out_id_0),
		.io_out_last_0(_mesh_1_27_io_out_last_0),
		.io_out_valid_0(_mesh_1_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9430 == GlobalFiModInstNr[0]) || (9430 == GlobalFiModInstNr[1]) || (9430 == GlobalFiModInstNr[2]) || (9430 == GlobalFiModInstNr[3]))));
	Tile mesh_1_28(
		.clock(clock),
		.io_in_a_0(r_60_0),
		.io_in_b_0(b_897_0),
		.io_in_d_0(b_1921_0),
		.io_in_control_0_dataflow(mesh_1_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2945_0),
		.io_in_last_0(r_3969_0),
		.io_in_valid_0(r_1921_0),
		.io_out_a_0(_mesh_1_28_io_out_a_0),
		.io_out_c_0(_mesh_1_28_io_out_c_0),
		.io_out_b_0(_mesh_1_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_28_io_out_id_0),
		.io_out_last_0(_mesh_1_28_io_out_last_0),
		.io_out_valid_0(_mesh_1_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9431 == GlobalFiModInstNr[0]) || (9431 == GlobalFiModInstNr[1]) || (9431 == GlobalFiModInstNr[2]) || (9431 == GlobalFiModInstNr[3]))));
	Tile mesh_1_29(
		.clock(clock),
		.io_in_a_0(r_61_0),
		.io_in_b_0(b_929_0),
		.io_in_d_0(b_1953_0),
		.io_in_control_0_dataflow(mesh_1_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2977_0),
		.io_in_last_0(r_4001_0),
		.io_in_valid_0(r_1953_0),
		.io_out_a_0(_mesh_1_29_io_out_a_0),
		.io_out_c_0(_mesh_1_29_io_out_c_0),
		.io_out_b_0(_mesh_1_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_29_io_out_id_0),
		.io_out_last_0(_mesh_1_29_io_out_last_0),
		.io_out_valid_0(_mesh_1_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9432 == GlobalFiModInstNr[0]) || (9432 == GlobalFiModInstNr[1]) || (9432 == GlobalFiModInstNr[2]) || (9432 == GlobalFiModInstNr[3]))));
	Tile mesh_1_30(
		.clock(clock),
		.io_in_a_0(r_62_0),
		.io_in_b_0(b_961_0),
		.io_in_d_0(b_1985_0),
		.io_in_control_0_dataflow(mesh_1_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3009_0),
		.io_in_last_0(r_4033_0),
		.io_in_valid_0(r_1985_0),
		.io_out_a_0(_mesh_1_30_io_out_a_0),
		.io_out_c_0(_mesh_1_30_io_out_c_0),
		.io_out_b_0(_mesh_1_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_30_io_out_id_0),
		.io_out_last_0(_mesh_1_30_io_out_last_0),
		.io_out_valid_0(_mesh_1_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9433 == GlobalFiModInstNr[0]) || (9433 == GlobalFiModInstNr[1]) || (9433 == GlobalFiModInstNr[2]) || (9433 == GlobalFiModInstNr[3]))));
	Tile mesh_1_31(
		.clock(clock),
		.io_in_a_0(r_63_0),
		.io_in_b_0(b_993_0),
		.io_in_d_0(b_2017_0),
		.io_in_control_0_dataflow(mesh_1_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3041_0),
		.io_in_last_0(r_4065_0),
		.io_in_valid_0(r_2017_0),
		.io_out_a_0(_mesh_1_31_io_out_a_0),
		.io_out_c_0(_mesh_1_31_io_out_c_0),
		.io_out_b_0(_mesh_1_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_31_io_out_id_0),
		.io_out_last_0(_mesh_1_31_io_out_last_0),
		.io_out_valid_0(_mesh_1_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9434 == GlobalFiModInstNr[0]) || (9434 == GlobalFiModInstNr[1]) || (9434 == GlobalFiModInstNr[2]) || (9434 == GlobalFiModInstNr[3]))));
	Tile mesh_2_0(
		.clock(clock),
		.io_in_a_0(r_64_0),
		.io_in_b_0(b_2_0),
		.io_in_d_0(b_1026_0),
		.io_in_control_0_dataflow(mesh_2_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2050_0),
		.io_in_last_0(r_3074_0),
		.io_in_valid_0(r_1026_0),
		.io_out_a_0(_mesh_2_0_io_out_a_0),
		.io_out_c_0(_mesh_2_0_io_out_c_0),
		.io_out_b_0(_mesh_2_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_0_io_out_id_0),
		.io_out_last_0(_mesh_2_0_io_out_last_0),
		.io_out_valid_0(_mesh_2_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9435 == GlobalFiModInstNr[0]) || (9435 == GlobalFiModInstNr[1]) || (9435 == GlobalFiModInstNr[2]) || (9435 == GlobalFiModInstNr[3]))));
	Tile mesh_2_1(
		.clock(clock),
		.io_in_a_0(r_65_0),
		.io_in_b_0(b_34_0),
		.io_in_d_0(b_1058_0),
		.io_in_control_0_dataflow(mesh_2_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2082_0),
		.io_in_last_0(r_3106_0),
		.io_in_valid_0(r_1058_0),
		.io_out_a_0(_mesh_2_1_io_out_a_0),
		.io_out_c_0(_mesh_2_1_io_out_c_0),
		.io_out_b_0(_mesh_2_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_1_io_out_id_0),
		.io_out_last_0(_mesh_2_1_io_out_last_0),
		.io_out_valid_0(_mesh_2_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9436 == GlobalFiModInstNr[0]) || (9436 == GlobalFiModInstNr[1]) || (9436 == GlobalFiModInstNr[2]) || (9436 == GlobalFiModInstNr[3]))));
	Tile mesh_2_2(
		.clock(clock),
		.io_in_a_0(r_66_0),
		.io_in_b_0(b_66_0),
		.io_in_d_0(b_1090_0),
		.io_in_control_0_dataflow(mesh_2_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2114_0),
		.io_in_last_0(r_3138_0),
		.io_in_valid_0(r_1090_0),
		.io_out_a_0(_mesh_2_2_io_out_a_0),
		.io_out_c_0(_mesh_2_2_io_out_c_0),
		.io_out_b_0(_mesh_2_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_2_io_out_id_0),
		.io_out_last_0(_mesh_2_2_io_out_last_0),
		.io_out_valid_0(_mesh_2_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9437 == GlobalFiModInstNr[0]) || (9437 == GlobalFiModInstNr[1]) || (9437 == GlobalFiModInstNr[2]) || (9437 == GlobalFiModInstNr[3]))));
	Tile mesh_2_3(
		.clock(clock),
		.io_in_a_0(r_67_0),
		.io_in_b_0(b_98_0),
		.io_in_d_0(b_1122_0),
		.io_in_control_0_dataflow(mesh_2_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2146_0),
		.io_in_last_0(r_3170_0),
		.io_in_valid_0(r_1122_0),
		.io_out_a_0(_mesh_2_3_io_out_a_0),
		.io_out_c_0(_mesh_2_3_io_out_c_0),
		.io_out_b_0(_mesh_2_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_3_io_out_id_0),
		.io_out_last_0(_mesh_2_3_io_out_last_0),
		.io_out_valid_0(_mesh_2_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9438 == GlobalFiModInstNr[0]) || (9438 == GlobalFiModInstNr[1]) || (9438 == GlobalFiModInstNr[2]) || (9438 == GlobalFiModInstNr[3]))));
	Tile mesh_2_4(
		.clock(clock),
		.io_in_a_0(r_68_0),
		.io_in_b_0(b_130_0),
		.io_in_d_0(b_1154_0),
		.io_in_control_0_dataflow(mesh_2_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2178_0),
		.io_in_last_0(r_3202_0),
		.io_in_valid_0(r_1154_0),
		.io_out_a_0(_mesh_2_4_io_out_a_0),
		.io_out_c_0(_mesh_2_4_io_out_c_0),
		.io_out_b_0(_mesh_2_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_4_io_out_id_0),
		.io_out_last_0(_mesh_2_4_io_out_last_0),
		.io_out_valid_0(_mesh_2_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9439 == GlobalFiModInstNr[0]) || (9439 == GlobalFiModInstNr[1]) || (9439 == GlobalFiModInstNr[2]) || (9439 == GlobalFiModInstNr[3]))));
	Tile mesh_2_5(
		.clock(clock),
		.io_in_a_0(r_69_0),
		.io_in_b_0(b_162_0),
		.io_in_d_0(b_1186_0),
		.io_in_control_0_dataflow(mesh_2_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2210_0),
		.io_in_last_0(r_3234_0),
		.io_in_valid_0(r_1186_0),
		.io_out_a_0(_mesh_2_5_io_out_a_0),
		.io_out_c_0(_mesh_2_5_io_out_c_0),
		.io_out_b_0(_mesh_2_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_5_io_out_id_0),
		.io_out_last_0(_mesh_2_5_io_out_last_0),
		.io_out_valid_0(_mesh_2_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9440 == GlobalFiModInstNr[0]) || (9440 == GlobalFiModInstNr[1]) || (9440 == GlobalFiModInstNr[2]) || (9440 == GlobalFiModInstNr[3]))));
	Tile mesh_2_6(
		.clock(clock),
		.io_in_a_0(r_70_0),
		.io_in_b_0(b_194_0),
		.io_in_d_0(b_1218_0),
		.io_in_control_0_dataflow(mesh_2_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2242_0),
		.io_in_last_0(r_3266_0),
		.io_in_valid_0(r_1218_0),
		.io_out_a_0(_mesh_2_6_io_out_a_0),
		.io_out_c_0(_mesh_2_6_io_out_c_0),
		.io_out_b_0(_mesh_2_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_6_io_out_id_0),
		.io_out_last_0(_mesh_2_6_io_out_last_0),
		.io_out_valid_0(_mesh_2_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9441 == GlobalFiModInstNr[0]) || (9441 == GlobalFiModInstNr[1]) || (9441 == GlobalFiModInstNr[2]) || (9441 == GlobalFiModInstNr[3]))));
	Tile mesh_2_7(
		.clock(clock),
		.io_in_a_0(r_71_0),
		.io_in_b_0(b_226_0),
		.io_in_d_0(b_1250_0),
		.io_in_control_0_dataflow(mesh_2_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2274_0),
		.io_in_last_0(r_3298_0),
		.io_in_valid_0(r_1250_0),
		.io_out_a_0(_mesh_2_7_io_out_a_0),
		.io_out_c_0(_mesh_2_7_io_out_c_0),
		.io_out_b_0(_mesh_2_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_7_io_out_id_0),
		.io_out_last_0(_mesh_2_7_io_out_last_0),
		.io_out_valid_0(_mesh_2_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9442 == GlobalFiModInstNr[0]) || (9442 == GlobalFiModInstNr[1]) || (9442 == GlobalFiModInstNr[2]) || (9442 == GlobalFiModInstNr[3]))));
	Tile mesh_2_8(
		.clock(clock),
		.io_in_a_0(r_72_0),
		.io_in_b_0(b_258_0),
		.io_in_d_0(b_1282_0),
		.io_in_control_0_dataflow(mesh_2_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2306_0),
		.io_in_last_0(r_3330_0),
		.io_in_valid_0(r_1282_0),
		.io_out_a_0(_mesh_2_8_io_out_a_0),
		.io_out_c_0(_mesh_2_8_io_out_c_0),
		.io_out_b_0(_mesh_2_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_8_io_out_id_0),
		.io_out_last_0(_mesh_2_8_io_out_last_0),
		.io_out_valid_0(_mesh_2_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9443 == GlobalFiModInstNr[0]) || (9443 == GlobalFiModInstNr[1]) || (9443 == GlobalFiModInstNr[2]) || (9443 == GlobalFiModInstNr[3]))));
	Tile mesh_2_9(
		.clock(clock),
		.io_in_a_0(r_73_0),
		.io_in_b_0(b_290_0),
		.io_in_d_0(b_1314_0),
		.io_in_control_0_dataflow(mesh_2_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2338_0),
		.io_in_last_0(r_3362_0),
		.io_in_valid_0(r_1314_0),
		.io_out_a_0(_mesh_2_9_io_out_a_0),
		.io_out_c_0(_mesh_2_9_io_out_c_0),
		.io_out_b_0(_mesh_2_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_9_io_out_id_0),
		.io_out_last_0(_mesh_2_9_io_out_last_0),
		.io_out_valid_0(_mesh_2_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9444 == GlobalFiModInstNr[0]) || (9444 == GlobalFiModInstNr[1]) || (9444 == GlobalFiModInstNr[2]) || (9444 == GlobalFiModInstNr[3]))));
	Tile mesh_2_10(
		.clock(clock),
		.io_in_a_0(r_74_0),
		.io_in_b_0(b_322_0),
		.io_in_d_0(b_1346_0),
		.io_in_control_0_dataflow(mesh_2_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2370_0),
		.io_in_last_0(r_3394_0),
		.io_in_valid_0(r_1346_0),
		.io_out_a_0(_mesh_2_10_io_out_a_0),
		.io_out_c_0(_mesh_2_10_io_out_c_0),
		.io_out_b_0(_mesh_2_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_10_io_out_id_0),
		.io_out_last_0(_mesh_2_10_io_out_last_0),
		.io_out_valid_0(_mesh_2_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9445 == GlobalFiModInstNr[0]) || (9445 == GlobalFiModInstNr[1]) || (9445 == GlobalFiModInstNr[2]) || (9445 == GlobalFiModInstNr[3]))));
	Tile mesh_2_11(
		.clock(clock),
		.io_in_a_0(r_75_0),
		.io_in_b_0(b_354_0),
		.io_in_d_0(b_1378_0),
		.io_in_control_0_dataflow(mesh_2_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2402_0),
		.io_in_last_0(r_3426_0),
		.io_in_valid_0(r_1378_0),
		.io_out_a_0(_mesh_2_11_io_out_a_0),
		.io_out_c_0(_mesh_2_11_io_out_c_0),
		.io_out_b_0(_mesh_2_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_11_io_out_id_0),
		.io_out_last_0(_mesh_2_11_io_out_last_0),
		.io_out_valid_0(_mesh_2_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9446 == GlobalFiModInstNr[0]) || (9446 == GlobalFiModInstNr[1]) || (9446 == GlobalFiModInstNr[2]) || (9446 == GlobalFiModInstNr[3]))));
	Tile mesh_2_12(
		.clock(clock),
		.io_in_a_0(r_76_0),
		.io_in_b_0(b_386_0),
		.io_in_d_0(b_1410_0),
		.io_in_control_0_dataflow(mesh_2_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2434_0),
		.io_in_last_0(r_3458_0),
		.io_in_valid_0(r_1410_0),
		.io_out_a_0(_mesh_2_12_io_out_a_0),
		.io_out_c_0(_mesh_2_12_io_out_c_0),
		.io_out_b_0(_mesh_2_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_12_io_out_id_0),
		.io_out_last_0(_mesh_2_12_io_out_last_0),
		.io_out_valid_0(_mesh_2_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9447 == GlobalFiModInstNr[0]) || (9447 == GlobalFiModInstNr[1]) || (9447 == GlobalFiModInstNr[2]) || (9447 == GlobalFiModInstNr[3]))));
	Tile mesh_2_13(
		.clock(clock),
		.io_in_a_0(r_77_0),
		.io_in_b_0(b_418_0),
		.io_in_d_0(b_1442_0),
		.io_in_control_0_dataflow(mesh_2_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2466_0),
		.io_in_last_0(r_3490_0),
		.io_in_valid_0(r_1442_0),
		.io_out_a_0(_mesh_2_13_io_out_a_0),
		.io_out_c_0(_mesh_2_13_io_out_c_0),
		.io_out_b_0(_mesh_2_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_13_io_out_id_0),
		.io_out_last_0(_mesh_2_13_io_out_last_0),
		.io_out_valid_0(_mesh_2_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9448 == GlobalFiModInstNr[0]) || (9448 == GlobalFiModInstNr[1]) || (9448 == GlobalFiModInstNr[2]) || (9448 == GlobalFiModInstNr[3]))));
	Tile mesh_2_14(
		.clock(clock),
		.io_in_a_0(r_78_0),
		.io_in_b_0(b_450_0),
		.io_in_d_0(b_1474_0),
		.io_in_control_0_dataflow(mesh_2_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2498_0),
		.io_in_last_0(r_3522_0),
		.io_in_valid_0(r_1474_0),
		.io_out_a_0(_mesh_2_14_io_out_a_0),
		.io_out_c_0(_mesh_2_14_io_out_c_0),
		.io_out_b_0(_mesh_2_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_14_io_out_id_0),
		.io_out_last_0(_mesh_2_14_io_out_last_0),
		.io_out_valid_0(_mesh_2_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9449 == GlobalFiModInstNr[0]) || (9449 == GlobalFiModInstNr[1]) || (9449 == GlobalFiModInstNr[2]) || (9449 == GlobalFiModInstNr[3]))));
	Tile mesh_2_15(
		.clock(clock),
		.io_in_a_0(r_79_0),
		.io_in_b_0(b_482_0),
		.io_in_d_0(b_1506_0),
		.io_in_control_0_dataflow(mesh_2_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2530_0),
		.io_in_last_0(r_3554_0),
		.io_in_valid_0(r_1506_0),
		.io_out_a_0(_mesh_2_15_io_out_a_0),
		.io_out_c_0(_mesh_2_15_io_out_c_0),
		.io_out_b_0(_mesh_2_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_15_io_out_id_0),
		.io_out_last_0(_mesh_2_15_io_out_last_0),
		.io_out_valid_0(_mesh_2_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9450 == GlobalFiModInstNr[0]) || (9450 == GlobalFiModInstNr[1]) || (9450 == GlobalFiModInstNr[2]) || (9450 == GlobalFiModInstNr[3]))));
	Tile mesh_2_16(
		.clock(clock),
		.io_in_a_0(r_80_0),
		.io_in_b_0(b_514_0),
		.io_in_d_0(b_1538_0),
		.io_in_control_0_dataflow(mesh_2_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2562_0),
		.io_in_last_0(r_3586_0),
		.io_in_valid_0(r_1538_0),
		.io_out_a_0(_mesh_2_16_io_out_a_0),
		.io_out_c_0(_mesh_2_16_io_out_c_0),
		.io_out_b_0(_mesh_2_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_16_io_out_id_0),
		.io_out_last_0(_mesh_2_16_io_out_last_0),
		.io_out_valid_0(_mesh_2_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9451 == GlobalFiModInstNr[0]) || (9451 == GlobalFiModInstNr[1]) || (9451 == GlobalFiModInstNr[2]) || (9451 == GlobalFiModInstNr[3]))));
	Tile mesh_2_17(
		.clock(clock),
		.io_in_a_0(r_81_0),
		.io_in_b_0(b_546_0),
		.io_in_d_0(b_1570_0),
		.io_in_control_0_dataflow(mesh_2_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2594_0),
		.io_in_last_0(r_3618_0),
		.io_in_valid_0(r_1570_0),
		.io_out_a_0(_mesh_2_17_io_out_a_0),
		.io_out_c_0(_mesh_2_17_io_out_c_0),
		.io_out_b_0(_mesh_2_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_17_io_out_id_0),
		.io_out_last_0(_mesh_2_17_io_out_last_0),
		.io_out_valid_0(_mesh_2_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9452 == GlobalFiModInstNr[0]) || (9452 == GlobalFiModInstNr[1]) || (9452 == GlobalFiModInstNr[2]) || (9452 == GlobalFiModInstNr[3]))));
	Tile mesh_2_18(
		.clock(clock),
		.io_in_a_0(r_82_0),
		.io_in_b_0(b_578_0),
		.io_in_d_0(b_1602_0),
		.io_in_control_0_dataflow(mesh_2_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2626_0),
		.io_in_last_0(r_3650_0),
		.io_in_valid_0(r_1602_0),
		.io_out_a_0(_mesh_2_18_io_out_a_0),
		.io_out_c_0(_mesh_2_18_io_out_c_0),
		.io_out_b_0(_mesh_2_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_18_io_out_id_0),
		.io_out_last_0(_mesh_2_18_io_out_last_0),
		.io_out_valid_0(_mesh_2_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9453 == GlobalFiModInstNr[0]) || (9453 == GlobalFiModInstNr[1]) || (9453 == GlobalFiModInstNr[2]) || (9453 == GlobalFiModInstNr[3]))));
	Tile mesh_2_19(
		.clock(clock),
		.io_in_a_0(r_83_0),
		.io_in_b_0(b_610_0),
		.io_in_d_0(b_1634_0),
		.io_in_control_0_dataflow(mesh_2_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2658_0),
		.io_in_last_0(r_3682_0),
		.io_in_valid_0(r_1634_0),
		.io_out_a_0(_mesh_2_19_io_out_a_0),
		.io_out_c_0(_mesh_2_19_io_out_c_0),
		.io_out_b_0(_mesh_2_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_19_io_out_id_0),
		.io_out_last_0(_mesh_2_19_io_out_last_0),
		.io_out_valid_0(_mesh_2_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9454 == GlobalFiModInstNr[0]) || (9454 == GlobalFiModInstNr[1]) || (9454 == GlobalFiModInstNr[2]) || (9454 == GlobalFiModInstNr[3]))));
	Tile mesh_2_20(
		.clock(clock),
		.io_in_a_0(r_84_0),
		.io_in_b_0(b_642_0),
		.io_in_d_0(b_1666_0),
		.io_in_control_0_dataflow(mesh_2_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2690_0),
		.io_in_last_0(r_3714_0),
		.io_in_valid_0(r_1666_0),
		.io_out_a_0(_mesh_2_20_io_out_a_0),
		.io_out_c_0(_mesh_2_20_io_out_c_0),
		.io_out_b_0(_mesh_2_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_20_io_out_id_0),
		.io_out_last_0(_mesh_2_20_io_out_last_0),
		.io_out_valid_0(_mesh_2_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9455 == GlobalFiModInstNr[0]) || (9455 == GlobalFiModInstNr[1]) || (9455 == GlobalFiModInstNr[2]) || (9455 == GlobalFiModInstNr[3]))));
	Tile mesh_2_21(
		.clock(clock),
		.io_in_a_0(r_85_0),
		.io_in_b_0(b_674_0),
		.io_in_d_0(b_1698_0),
		.io_in_control_0_dataflow(mesh_2_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2722_0),
		.io_in_last_0(r_3746_0),
		.io_in_valid_0(r_1698_0),
		.io_out_a_0(_mesh_2_21_io_out_a_0),
		.io_out_c_0(_mesh_2_21_io_out_c_0),
		.io_out_b_0(_mesh_2_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_21_io_out_id_0),
		.io_out_last_0(_mesh_2_21_io_out_last_0),
		.io_out_valid_0(_mesh_2_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9456 == GlobalFiModInstNr[0]) || (9456 == GlobalFiModInstNr[1]) || (9456 == GlobalFiModInstNr[2]) || (9456 == GlobalFiModInstNr[3]))));
	Tile mesh_2_22(
		.clock(clock),
		.io_in_a_0(r_86_0),
		.io_in_b_0(b_706_0),
		.io_in_d_0(b_1730_0),
		.io_in_control_0_dataflow(mesh_2_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2754_0),
		.io_in_last_0(r_3778_0),
		.io_in_valid_0(r_1730_0),
		.io_out_a_0(_mesh_2_22_io_out_a_0),
		.io_out_c_0(_mesh_2_22_io_out_c_0),
		.io_out_b_0(_mesh_2_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_22_io_out_id_0),
		.io_out_last_0(_mesh_2_22_io_out_last_0),
		.io_out_valid_0(_mesh_2_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9457 == GlobalFiModInstNr[0]) || (9457 == GlobalFiModInstNr[1]) || (9457 == GlobalFiModInstNr[2]) || (9457 == GlobalFiModInstNr[3]))));
	Tile mesh_2_23(
		.clock(clock),
		.io_in_a_0(r_87_0),
		.io_in_b_0(b_738_0),
		.io_in_d_0(b_1762_0),
		.io_in_control_0_dataflow(mesh_2_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2786_0),
		.io_in_last_0(r_3810_0),
		.io_in_valid_0(r_1762_0),
		.io_out_a_0(_mesh_2_23_io_out_a_0),
		.io_out_c_0(_mesh_2_23_io_out_c_0),
		.io_out_b_0(_mesh_2_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_23_io_out_id_0),
		.io_out_last_0(_mesh_2_23_io_out_last_0),
		.io_out_valid_0(_mesh_2_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9458 == GlobalFiModInstNr[0]) || (9458 == GlobalFiModInstNr[1]) || (9458 == GlobalFiModInstNr[2]) || (9458 == GlobalFiModInstNr[3]))));
	Tile mesh_2_24(
		.clock(clock),
		.io_in_a_0(r_88_0),
		.io_in_b_0(b_770_0),
		.io_in_d_0(b_1794_0),
		.io_in_control_0_dataflow(mesh_2_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2818_0),
		.io_in_last_0(r_3842_0),
		.io_in_valid_0(r_1794_0),
		.io_out_a_0(_mesh_2_24_io_out_a_0),
		.io_out_c_0(_mesh_2_24_io_out_c_0),
		.io_out_b_0(_mesh_2_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_24_io_out_id_0),
		.io_out_last_0(_mesh_2_24_io_out_last_0),
		.io_out_valid_0(_mesh_2_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9459 == GlobalFiModInstNr[0]) || (9459 == GlobalFiModInstNr[1]) || (9459 == GlobalFiModInstNr[2]) || (9459 == GlobalFiModInstNr[3]))));
	Tile mesh_2_25(
		.clock(clock),
		.io_in_a_0(r_89_0),
		.io_in_b_0(b_802_0),
		.io_in_d_0(b_1826_0),
		.io_in_control_0_dataflow(mesh_2_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2850_0),
		.io_in_last_0(r_3874_0),
		.io_in_valid_0(r_1826_0),
		.io_out_a_0(_mesh_2_25_io_out_a_0),
		.io_out_c_0(_mesh_2_25_io_out_c_0),
		.io_out_b_0(_mesh_2_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_25_io_out_id_0),
		.io_out_last_0(_mesh_2_25_io_out_last_0),
		.io_out_valid_0(_mesh_2_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9460 == GlobalFiModInstNr[0]) || (9460 == GlobalFiModInstNr[1]) || (9460 == GlobalFiModInstNr[2]) || (9460 == GlobalFiModInstNr[3]))));
	Tile mesh_2_26(
		.clock(clock),
		.io_in_a_0(r_90_0),
		.io_in_b_0(b_834_0),
		.io_in_d_0(b_1858_0),
		.io_in_control_0_dataflow(mesh_2_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2882_0),
		.io_in_last_0(r_3906_0),
		.io_in_valid_0(r_1858_0),
		.io_out_a_0(_mesh_2_26_io_out_a_0),
		.io_out_c_0(_mesh_2_26_io_out_c_0),
		.io_out_b_0(_mesh_2_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_26_io_out_id_0),
		.io_out_last_0(_mesh_2_26_io_out_last_0),
		.io_out_valid_0(_mesh_2_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9461 == GlobalFiModInstNr[0]) || (9461 == GlobalFiModInstNr[1]) || (9461 == GlobalFiModInstNr[2]) || (9461 == GlobalFiModInstNr[3]))));
	Tile mesh_2_27(
		.clock(clock),
		.io_in_a_0(r_91_0),
		.io_in_b_0(b_866_0),
		.io_in_d_0(b_1890_0),
		.io_in_control_0_dataflow(mesh_2_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2914_0),
		.io_in_last_0(r_3938_0),
		.io_in_valid_0(r_1890_0),
		.io_out_a_0(_mesh_2_27_io_out_a_0),
		.io_out_c_0(_mesh_2_27_io_out_c_0),
		.io_out_b_0(_mesh_2_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_27_io_out_id_0),
		.io_out_last_0(_mesh_2_27_io_out_last_0),
		.io_out_valid_0(_mesh_2_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9462 == GlobalFiModInstNr[0]) || (9462 == GlobalFiModInstNr[1]) || (9462 == GlobalFiModInstNr[2]) || (9462 == GlobalFiModInstNr[3]))));
	Tile mesh_2_28(
		.clock(clock),
		.io_in_a_0(r_92_0),
		.io_in_b_0(b_898_0),
		.io_in_d_0(b_1922_0),
		.io_in_control_0_dataflow(mesh_2_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2946_0),
		.io_in_last_0(r_3970_0),
		.io_in_valid_0(r_1922_0),
		.io_out_a_0(_mesh_2_28_io_out_a_0),
		.io_out_c_0(_mesh_2_28_io_out_c_0),
		.io_out_b_0(_mesh_2_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_28_io_out_id_0),
		.io_out_last_0(_mesh_2_28_io_out_last_0),
		.io_out_valid_0(_mesh_2_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9463 == GlobalFiModInstNr[0]) || (9463 == GlobalFiModInstNr[1]) || (9463 == GlobalFiModInstNr[2]) || (9463 == GlobalFiModInstNr[3]))));
	Tile mesh_2_29(
		.clock(clock),
		.io_in_a_0(r_93_0),
		.io_in_b_0(b_930_0),
		.io_in_d_0(b_1954_0),
		.io_in_control_0_dataflow(mesh_2_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2978_0),
		.io_in_last_0(r_4002_0),
		.io_in_valid_0(r_1954_0),
		.io_out_a_0(_mesh_2_29_io_out_a_0),
		.io_out_c_0(_mesh_2_29_io_out_c_0),
		.io_out_b_0(_mesh_2_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_29_io_out_id_0),
		.io_out_last_0(_mesh_2_29_io_out_last_0),
		.io_out_valid_0(_mesh_2_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9464 == GlobalFiModInstNr[0]) || (9464 == GlobalFiModInstNr[1]) || (9464 == GlobalFiModInstNr[2]) || (9464 == GlobalFiModInstNr[3]))));
	Tile mesh_2_30(
		.clock(clock),
		.io_in_a_0(r_94_0),
		.io_in_b_0(b_962_0),
		.io_in_d_0(b_1986_0),
		.io_in_control_0_dataflow(mesh_2_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3010_0),
		.io_in_last_0(r_4034_0),
		.io_in_valid_0(r_1986_0),
		.io_out_a_0(_mesh_2_30_io_out_a_0),
		.io_out_c_0(_mesh_2_30_io_out_c_0),
		.io_out_b_0(_mesh_2_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_30_io_out_id_0),
		.io_out_last_0(_mesh_2_30_io_out_last_0),
		.io_out_valid_0(_mesh_2_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9465 == GlobalFiModInstNr[0]) || (9465 == GlobalFiModInstNr[1]) || (9465 == GlobalFiModInstNr[2]) || (9465 == GlobalFiModInstNr[3]))));
	Tile mesh_2_31(
		.clock(clock),
		.io_in_a_0(r_95_0),
		.io_in_b_0(b_994_0),
		.io_in_d_0(b_2018_0),
		.io_in_control_0_dataflow(mesh_2_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3042_0),
		.io_in_last_0(r_4066_0),
		.io_in_valid_0(r_2018_0),
		.io_out_a_0(_mesh_2_31_io_out_a_0),
		.io_out_c_0(_mesh_2_31_io_out_c_0),
		.io_out_b_0(_mesh_2_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_31_io_out_id_0),
		.io_out_last_0(_mesh_2_31_io_out_last_0),
		.io_out_valid_0(_mesh_2_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9466 == GlobalFiModInstNr[0]) || (9466 == GlobalFiModInstNr[1]) || (9466 == GlobalFiModInstNr[2]) || (9466 == GlobalFiModInstNr[3]))));
	Tile mesh_3_0(
		.clock(clock),
		.io_in_a_0(r_96_0),
		.io_in_b_0(b_3_0),
		.io_in_d_0(b_1027_0),
		.io_in_control_0_dataflow(mesh_3_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2051_0),
		.io_in_last_0(r_3075_0),
		.io_in_valid_0(r_1027_0),
		.io_out_a_0(_mesh_3_0_io_out_a_0),
		.io_out_c_0(_mesh_3_0_io_out_c_0),
		.io_out_b_0(_mesh_3_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_0_io_out_id_0),
		.io_out_last_0(_mesh_3_0_io_out_last_0),
		.io_out_valid_0(_mesh_3_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9467 == GlobalFiModInstNr[0]) || (9467 == GlobalFiModInstNr[1]) || (9467 == GlobalFiModInstNr[2]) || (9467 == GlobalFiModInstNr[3]))));
	Tile mesh_3_1(
		.clock(clock),
		.io_in_a_0(r_97_0),
		.io_in_b_0(b_35_0),
		.io_in_d_0(b_1059_0),
		.io_in_control_0_dataflow(mesh_3_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2083_0),
		.io_in_last_0(r_3107_0),
		.io_in_valid_0(r_1059_0),
		.io_out_a_0(_mesh_3_1_io_out_a_0),
		.io_out_c_0(_mesh_3_1_io_out_c_0),
		.io_out_b_0(_mesh_3_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_1_io_out_id_0),
		.io_out_last_0(_mesh_3_1_io_out_last_0),
		.io_out_valid_0(_mesh_3_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9468 == GlobalFiModInstNr[0]) || (9468 == GlobalFiModInstNr[1]) || (9468 == GlobalFiModInstNr[2]) || (9468 == GlobalFiModInstNr[3]))));
	Tile mesh_3_2(
		.clock(clock),
		.io_in_a_0(r_98_0),
		.io_in_b_0(b_67_0),
		.io_in_d_0(b_1091_0),
		.io_in_control_0_dataflow(mesh_3_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2115_0),
		.io_in_last_0(r_3139_0),
		.io_in_valid_0(r_1091_0),
		.io_out_a_0(_mesh_3_2_io_out_a_0),
		.io_out_c_0(_mesh_3_2_io_out_c_0),
		.io_out_b_0(_mesh_3_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_2_io_out_id_0),
		.io_out_last_0(_mesh_3_2_io_out_last_0),
		.io_out_valid_0(_mesh_3_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9469 == GlobalFiModInstNr[0]) || (9469 == GlobalFiModInstNr[1]) || (9469 == GlobalFiModInstNr[2]) || (9469 == GlobalFiModInstNr[3]))));
	Tile mesh_3_3(
		.clock(clock),
		.io_in_a_0(r_99_0),
		.io_in_b_0(b_99_0),
		.io_in_d_0(b_1123_0),
		.io_in_control_0_dataflow(mesh_3_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2147_0),
		.io_in_last_0(r_3171_0),
		.io_in_valid_0(r_1123_0),
		.io_out_a_0(_mesh_3_3_io_out_a_0),
		.io_out_c_0(_mesh_3_3_io_out_c_0),
		.io_out_b_0(_mesh_3_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_3_io_out_id_0),
		.io_out_last_0(_mesh_3_3_io_out_last_0),
		.io_out_valid_0(_mesh_3_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9470 == GlobalFiModInstNr[0]) || (9470 == GlobalFiModInstNr[1]) || (9470 == GlobalFiModInstNr[2]) || (9470 == GlobalFiModInstNr[3]))));
	Tile mesh_3_4(
		.clock(clock),
		.io_in_a_0(r_100_0),
		.io_in_b_0(b_131_0),
		.io_in_d_0(b_1155_0),
		.io_in_control_0_dataflow(mesh_3_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2179_0),
		.io_in_last_0(r_3203_0),
		.io_in_valid_0(r_1155_0),
		.io_out_a_0(_mesh_3_4_io_out_a_0),
		.io_out_c_0(_mesh_3_4_io_out_c_0),
		.io_out_b_0(_mesh_3_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_4_io_out_id_0),
		.io_out_last_0(_mesh_3_4_io_out_last_0),
		.io_out_valid_0(_mesh_3_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9471 == GlobalFiModInstNr[0]) || (9471 == GlobalFiModInstNr[1]) || (9471 == GlobalFiModInstNr[2]) || (9471 == GlobalFiModInstNr[3]))));
	Tile mesh_3_5(
		.clock(clock),
		.io_in_a_0(r_101_0),
		.io_in_b_0(b_163_0),
		.io_in_d_0(b_1187_0),
		.io_in_control_0_dataflow(mesh_3_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2211_0),
		.io_in_last_0(r_3235_0),
		.io_in_valid_0(r_1187_0),
		.io_out_a_0(_mesh_3_5_io_out_a_0),
		.io_out_c_0(_mesh_3_5_io_out_c_0),
		.io_out_b_0(_mesh_3_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_5_io_out_id_0),
		.io_out_last_0(_mesh_3_5_io_out_last_0),
		.io_out_valid_0(_mesh_3_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9472 == GlobalFiModInstNr[0]) || (9472 == GlobalFiModInstNr[1]) || (9472 == GlobalFiModInstNr[2]) || (9472 == GlobalFiModInstNr[3]))));
	Tile mesh_3_6(
		.clock(clock),
		.io_in_a_0(r_102_0),
		.io_in_b_0(b_195_0),
		.io_in_d_0(b_1219_0),
		.io_in_control_0_dataflow(mesh_3_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2243_0),
		.io_in_last_0(r_3267_0),
		.io_in_valid_0(r_1219_0),
		.io_out_a_0(_mesh_3_6_io_out_a_0),
		.io_out_c_0(_mesh_3_6_io_out_c_0),
		.io_out_b_0(_mesh_3_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_6_io_out_id_0),
		.io_out_last_0(_mesh_3_6_io_out_last_0),
		.io_out_valid_0(_mesh_3_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9473 == GlobalFiModInstNr[0]) || (9473 == GlobalFiModInstNr[1]) || (9473 == GlobalFiModInstNr[2]) || (9473 == GlobalFiModInstNr[3]))));
	Tile mesh_3_7(
		.clock(clock),
		.io_in_a_0(r_103_0),
		.io_in_b_0(b_227_0),
		.io_in_d_0(b_1251_0),
		.io_in_control_0_dataflow(mesh_3_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2275_0),
		.io_in_last_0(r_3299_0),
		.io_in_valid_0(r_1251_0),
		.io_out_a_0(_mesh_3_7_io_out_a_0),
		.io_out_c_0(_mesh_3_7_io_out_c_0),
		.io_out_b_0(_mesh_3_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_7_io_out_id_0),
		.io_out_last_0(_mesh_3_7_io_out_last_0),
		.io_out_valid_0(_mesh_3_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9474 == GlobalFiModInstNr[0]) || (9474 == GlobalFiModInstNr[1]) || (9474 == GlobalFiModInstNr[2]) || (9474 == GlobalFiModInstNr[3]))));
	Tile mesh_3_8(
		.clock(clock),
		.io_in_a_0(r_104_0),
		.io_in_b_0(b_259_0),
		.io_in_d_0(b_1283_0),
		.io_in_control_0_dataflow(mesh_3_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2307_0),
		.io_in_last_0(r_3331_0),
		.io_in_valid_0(r_1283_0),
		.io_out_a_0(_mesh_3_8_io_out_a_0),
		.io_out_c_0(_mesh_3_8_io_out_c_0),
		.io_out_b_0(_mesh_3_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_8_io_out_id_0),
		.io_out_last_0(_mesh_3_8_io_out_last_0),
		.io_out_valid_0(_mesh_3_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9475 == GlobalFiModInstNr[0]) || (9475 == GlobalFiModInstNr[1]) || (9475 == GlobalFiModInstNr[2]) || (9475 == GlobalFiModInstNr[3]))));
	Tile mesh_3_9(
		.clock(clock),
		.io_in_a_0(r_105_0),
		.io_in_b_0(b_291_0),
		.io_in_d_0(b_1315_0),
		.io_in_control_0_dataflow(mesh_3_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2339_0),
		.io_in_last_0(r_3363_0),
		.io_in_valid_0(r_1315_0),
		.io_out_a_0(_mesh_3_9_io_out_a_0),
		.io_out_c_0(_mesh_3_9_io_out_c_0),
		.io_out_b_0(_mesh_3_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_9_io_out_id_0),
		.io_out_last_0(_mesh_3_9_io_out_last_0),
		.io_out_valid_0(_mesh_3_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9476 == GlobalFiModInstNr[0]) || (9476 == GlobalFiModInstNr[1]) || (9476 == GlobalFiModInstNr[2]) || (9476 == GlobalFiModInstNr[3]))));
	Tile mesh_3_10(
		.clock(clock),
		.io_in_a_0(r_106_0),
		.io_in_b_0(b_323_0),
		.io_in_d_0(b_1347_0),
		.io_in_control_0_dataflow(mesh_3_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2371_0),
		.io_in_last_0(r_3395_0),
		.io_in_valid_0(r_1347_0),
		.io_out_a_0(_mesh_3_10_io_out_a_0),
		.io_out_c_0(_mesh_3_10_io_out_c_0),
		.io_out_b_0(_mesh_3_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_10_io_out_id_0),
		.io_out_last_0(_mesh_3_10_io_out_last_0),
		.io_out_valid_0(_mesh_3_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9477 == GlobalFiModInstNr[0]) || (9477 == GlobalFiModInstNr[1]) || (9477 == GlobalFiModInstNr[2]) || (9477 == GlobalFiModInstNr[3]))));
	Tile mesh_3_11(
		.clock(clock),
		.io_in_a_0(r_107_0),
		.io_in_b_0(b_355_0),
		.io_in_d_0(b_1379_0),
		.io_in_control_0_dataflow(mesh_3_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2403_0),
		.io_in_last_0(r_3427_0),
		.io_in_valid_0(r_1379_0),
		.io_out_a_0(_mesh_3_11_io_out_a_0),
		.io_out_c_0(_mesh_3_11_io_out_c_0),
		.io_out_b_0(_mesh_3_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_11_io_out_id_0),
		.io_out_last_0(_mesh_3_11_io_out_last_0),
		.io_out_valid_0(_mesh_3_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9478 == GlobalFiModInstNr[0]) || (9478 == GlobalFiModInstNr[1]) || (9478 == GlobalFiModInstNr[2]) || (9478 == GlobalFiModInstNr[3]))));
	Tile mesh_3_12(
		.clock(clock),
		.io_in_a_0(r_108_0),
		.io_in_b_0(b_387_0),
		.io_in_d_0(b_1411_0),
		.io_in_control_0_dataflow(mesh_3_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2435_0),
		.io_in_last_0(r_3459_0),
		.io_in_valid_0(r_1411_0),
		.io_out_a_0(_mesh_3_12_io_out_a_0),
		.io_out_c_0(_mesh_3_12_io_out_c_0),
		.io_out_b_0(_mesh_3_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_12_io_out_id_0),
		.io_out_last_0(_mesh_3_12_io_out_last_0),
		.io_out_valid_0(_mesh_3_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9479 == GlobalFiModInstNr[0]) || (9479 == GlobalFiModInstNr[1]) || (9479 == GlobalFiModInstNr[2]) || (9479 == GlobalFiModInstNr[3]))));
	Tile mesh_3_13(
		.clock(clock),
		.io_in_a_0(r_109_0),
		.io_in_b_0(b_419_0),
		.io_in_d_0(b_1443_0),
		.io_in_control_0_dataflow(mesh_3_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2467_0),
		.io_in_last_0(r_3491_0),
		.io_in_valid_0(r_1443_0),
		.io_out_a_0(_mesh_3_13_io_out_a_0),
		.io_out_c_0(_mesh_3_13_io_out_c_0),
		.io_out_b_0(_mesh_3_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_13_io_out_id_0),
		.io_out_last_0(_mesh_3_13_io_out_last_0),
		.io_out_valid_0(_mesh_3_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9480 == GlobalFiModInstNr[0]) || (9480 == GlobalFiModInstNr[1]) || (9480 == GlobalFiModInstNr[2]) || (9480 == GlobalFiModInstNr[3]))));
	Tile mesh_3_14(
		.clock(clock),
		.io_in_a_0(r_110_0),
		.io_in_b_0(b_451_0),
		.io_in_d_0(b_1475_0),
		.io_in_control_0_dataflow(mesh_3_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2499_0),
		.io_in_last_0(r_3523_0),
		.io_in_valid_0(r_1475_0),
		.io_out_a_0(_mesh_3_14_io_out_a_0),
		.io_out_c_0(_mesh_3_14_io_out_c_0),
		.io_out_b_0(_mesh_3_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_14_io_out_id_0),
		.io_out_last_0(_mesh_3_14_io_out_last_0),
		.io_out_valid_0(_mesh_3_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9481 == GlobalFiModInstNr[0]) || (9481 == GlobalFiModInstNr[1]) || (9481 == GlobalFiModInstNr[2]) || (9481 == GlobalFiModInstNr[3]))));
	Tile mesh_3_15(
		.clock(clock),
		.io_in_a_0(r_111_0),
		.io_in_b_0(b_483_0),
		.io_in_d_0(b_1507_0),
		.io_in_control_0_dataflow(mesh_3_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2531_0),
		.io_in_last_0(r_3555_0),
		.io_in_valid_0(r_1507_0),
		.io_out_a_0(_mesh_3_15_io_out_a_0),
		.io_out_c_0(_mesh_3_15_io_out_c_0),
		.io_out_b_0(_mesh_3_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_15_io_out_id_0),
		.io_out_last_0(_mesh_3_15_io_out_last_0),
		.io_out_valid_0(_mesh_3_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9482 == GlobalFiModInstNr[0]) || (9482 == GlobalFiModInstNr[1]) || (9482 == GlobalFiModInstNr[2]) || (9482 == GlobalFiModInstNr[3]))));
	Tile mesh_3_16(
		.clock(clock),
		.io_in_a_0(r_112_0),
		.io_in_b_0(b_515_0),
		.io_in_d_0(b_1539_0),
		.io_in_control_0_dataflow(mesh_3_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2563_0),
		.io_in_last_0(r_3587_0),
		.io_in_valid_0(r_1539_0),
		.io_out_a_0(_mesh_3_16_io_out_a_0),
		.io_out_c_0(_mesh_3_16_io_out_c_0),
		.io_out_b_0(_mesh_3_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_16_io_out_id_0),
		.io_out_last_0(_mesh_3_16_io_out_last_0),
		.io_out_valid_0(_mesh_3_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9483 == GlobalFiModInstNr[0]) || (9483 == GlobalFiModInstNr[1]) || (9483 == GlobalFiModInstNr[2]) || (9483 == GlobalFiModInstNr[3]))));
	Tile mesh_3_17(
		.clock(clock),
		.io_in_a_0(r_113_0),
		.io_in_b_0(b_547_0),
		.io_in_d_0(b_1571_0),
		.io_in_control_0_dataflow(mesh_3_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2595_0),
		.io_in_last_0(r_3619_0),
		.io_in_valid_0(r_1571_0),
		.io_out_a_0(_mesh_3_17_io_out_a_0),
		.io_out_c_0(_mesh_3_17_io_out_c_0),
		.io_out_b_0(_mesh_3_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_17_io_out_id_0),
		.io_out_last_0(_mesh_3_17_io_out_last_0),
		.io_out_valid_0(_mesh_3_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9484 == GlobalFiModInstNr[0]) || (9484 == GlobalFiModInstNr[1]) || (9484 == GlobalFiModInstNr[2]) || (9484 == GlobalFiModInstNr[3]))));
	Tile mesh_3_18(
		.clock(clock),
		.io_in_a_0(r_114_0),
		.io_in_b_0(b_579_0),
		.io_in_d_0(b_1603_0),
		.io_in_control_0_dataflow(mesh_3_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2627_0),
		.io_in_last_0(r_3651_0),
		.io_in_valid_0(r_1603_0),
		.io_out_a_0(_mesh_3_18_io_out_a_0),
		.io_out_c_0(_mesh_3_18_io_out_c_0),
		.io_out_b_0(_mesh_3_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_18_io_out_id_0),
		.io_out_last_0(_mesh_3_18_io_out_last_0),
		.io_out_valid_0(_mesh_3_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9485 == GlobalFiModInstNr[0]) || (9485 == GlobalFiModInstNr[1]) || (9485 == GlobalFiModInstNr[2]) || (9485 == GlobalFiModInstNr[3]))));
	Tile mesh_3_19(
		.clock(clock),
		.io_in_a_0(r_115_0),
		.io_in_b_0(b_611_0),
		.io_in_d_0(b_1635_0),
		.io_in_control_0_dataflow(mesh_3_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2659_0),
		.io_in_last_0(r_3683_0),
		.io_in_valid_0(r_1635_0),
		.io_out_a_0(_mesh_3_19_io_out_a_0),
		.io_out_c_0(_mesh_3_19_io_out_c_0),
		.io_out_b_0(_mesh_3_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_19_io_out_id_0),
		.io_out_last_0(_mesh_3_19_io_out_last_0),
		.io_out_valid_0(_mesh_3_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9486 == GlobalFiModInstNr[0]) || (9486 == GlobalFiModInstNr[1]) || (9486 == GlobalFiModInstNr[2]) || (9486 == GlobalFiModInstNr[3]))));
	Tile mesh_3_20(
		.clock(clock),
		.io_in_a_0(r_116_0),
		.io_in_b_0(b_643_0),
		.io_in_d_0(b_1667_0),
		.io_in_control_0_dataflow(mesh_3_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2691_0),
		.io_in_last_0(r_3715_0),
		.io_in_valid_0(r_1667_0),
		.io_out_a_0(_mesh_3_20_io_out_a_0),
		.io_out_c_0(_mesh_3_20_io_out_c_0),
		.io_out_b_0(_mesh_3_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_20_io_out_id_0),
		.io_out_last_0(_mesh_3_20_io_out_last_0),
		.io_out_valid_0(_mesh_3_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9487 == GlobalFiModInstNr[0]) || (9487 == GlobalFiModInstNr[1]) || (9487 == GlobalFiModInstNr[2]) || (9487 == GlobalFiModInstNr[3]))));
	Tile mesh_3_21(
		.clock(clock),
		.io_in_a_0(r_117_0),
		.io_in_b_0(b_675_0),
		.io_in_d_0(b_1699_0),
		.io_in_control_0_dataflow(mesh_3_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2723_0),
		.io_in_last_0(r_3747_0),
		.io_in_valid_0(r_1699_0),
		.io_out_a_0(_mesh_3_21_io_out_a_0),
		.io_out_c_0(_mesh_3_21_io_out_c_0),
		.io_out_b_0(_mesh_3_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_21_io_out_id_0),
		.io_out_last_0(_mesh_3_21_io_out_last_0),
		.io_out_valid_0(_mesh_3_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9488 == GlobalFiModInstNr[0]) || (9488 == GlobalFiModInstNr[1]) || (9488 == GlobalFiModInstNr[2]) || (9488 == GlobalFiModInstNr[3]))));
	Tile mesh_3_22(
		.clock(clock),
		.io_in_a_0(r_118_0),
		.io_in_b_0(b_707_0),
		.io_in_d_0(b_1731_0),
		.io_in_control_0_dataflow(mesh_3_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2755_0),
		.io_in_last_0(r_3779_0),
		.io_in_valid_0(r_1731_0),
		.io_out_a_0(_mesh_3_22_io_out_a_0),
		.io_out_c_0(_mesh_3_22_io_out_c_0),
		.io_out_b_0(_mesh_3_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_22_io_out_id_0),
		.io_out_last_0(_mesh_3_22_io_out_last_0),
		.io_out_valid_0(_mesh_3_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9489 == GlobalFiModInstNr[0]) || (9489 == GlobalFiModInstNr[1]) || (9489 == GlobalFiModInstNr[2]) || (9489 == GlobalFiModInstNr[3]))));
	Tile mesh_3_23(
		.clock(clock),
		.io_in_a_0(r_119_0),
		.io_in_b_0(b_739_0),
		.io_in_d_0(b_1763_0),
		.io_in_control_0_dataflow(mesh_3_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2787_0),
		.io_in_last_0(r_3811_0),
		.io_in_valid_0(r_1763_0),
		.io_out_a_0(_mesh_3_23_io_out_a_0),
		.io_out_c_0(_mesh_3_23_io_out_c_0),
		.io_out_b_0(_mesh_3_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_23_io_out_id_0),
		.io_out_last_0(_mesh_3_23_io_out_last_0),
		.io_out_valid_0(_mesh_3_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9490 == GlobalFiModInstNr[0]) || (9490 == GlobalFiModInstNr[1]) || (9490 == GlobalFiModInstNr[2]) || (9490 == GlobalFiModInstNr[3]))));
	Tile mesh_3_24(
		.clock(clock),
		.io_in_a_0(r_120_0),
		.io_in_b_0(b_771_0),
		.io_in_d_0(b_1795_0),
		.io_in_control_0_dataflow(mesh_3_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2819_0),
		.io_in_last_0(r_3843_0),
		.io_in_valid_0(r_1795_0),
		.io_out_a_0(_mesh_3_24_io_out_a_0),
		.io_out_c_0(_mesh_3_24_io_out_c_0),
		.io_out_b_0(_mesh_3_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_24_io_out_id_0),
		.io_out_last_0(_mesh_3_24_io_out_last_0),
		.io_out_valid_0(_mesh_3_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9491 == GlobalFiModInstNr[0]) || (9491 == GlobalFiModInstNr[1]) || (9491 == GlobalFiModInstNr[2]) || (9491 == GlobalFiModInstNr[3]))));
	Tile mesh_3_25(
		.clock(clock),
		.io_in_a_0(r_121_0),
		.io_in_b_0(b_803_0),
		.io_in_d_0(b_1827_0),
		.io_in_control_0_dataflow(mesh_3_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2851_0),
		.io_in_last_0(r_3875_0),
		.io_in_valid_0(r_1827_0),
		.io_out_a_0(_mesh_3_25_io_out_a_0),
		.io_out_c_0(_mesh_3_25_io_out_c_0),
		.io_out_b_0(_mesh_3_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_25_io_out_id_0),
		.io_out_last_0(_mesh_3_25_io_out_last_0),
		.io_out_valid_0(_mesh_3_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9492 == GlobalFiModInstNr[0]) || (9492 == GlobalFiModInstNr[1]) || (9492 == GlobalFiModInstNr[2]) || (9492 == GlobalFiModInstNr[3]))));
	Tile mesh_3_26(
		.clock(clock),
		.io_in_a_0(r_122_0),
		.io_in_b_0(b_835_0),
		.io_in_d_0(b_1859_0),
		.io_in_control_0_dataflow(mesh_3_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2883_0),
		.io_in_last_0(r_3907_0),
		.io_in_valid_0(r_1859_0),
		.io_out_a_0(_mesh_3_26_io_out_a_0),
		.io_out_c_0(_mesh_3_26_io_out_c_0),
		.io_out_b_0(_mesh_3_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_26_io_out_id_0),
		.io_out_last_0(_mesh_3_26_io_out_last_0),
		.io_out_valid_0(_mesh_3_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9493 == GlobalFiModInstNr[0]) || (9493 == GlobalFiModInstNr[1]) || (9493 == GlobalFiModInstNr[2]) || (9493 == GlobalFiModInstNr[3]))));
	Tile mesh_3_27(
		.clock(clock),
		.io_in_a_0(r_123_0),
		.io_in_b_0(b_867_0),
		.io_in_d_0(b_1891_0),
		.io_in_control_0_dataflow(mesh_3_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2915_0),
		.io_in_last_0(r_3939_0),
		.io_in_valid_0(r_1891_0),
		.io_out_a_0(_mesh_3_27_io_out_a_0),
		.io_out_c_0(_mesh_3_27_io_out_c_0),
		.io_out_b_0(_mesh_3_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_27_io_out_id_0),
		.io_out_last_0(_mesh_3_27_io_out_last_0),
		.io_out_valid_0(_mesh_3_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9494 == GlobalFiModInstNr[0]) || (9494 == GlobalFiModInstNr[1]) || (9494 == GlobalFiModInstNr[2]) || (9494 == GlobalFiModInstNr[3]))));
	Tile mesh_3_28(
		.clock(clock),
		.io_in_a_0(r_124_0),
		.io_in_b_0(b_899_0),
		.io_in_d_0(b_1923_0),
		.io_in_control_0_dataflow(mesh_3_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2947_0),
		.io_in_last_0(r_3971_0),
		.io_in_valid_0(r_1923_0),
		.io_out_a_0(_mesh_3_28_io_out_a_0),
		.io_out_c_0(_mesh_3_28_io_out_c_0),
		.io_out_b_0(_mesh_3_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_28_io_out_id_0),
		.io_out_last_0(_mesh_3_28_io_out_last_0),
		.io_out_valid_0(_mesh_3_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9495 == GlobalFiModInstNr[0]) || (9495 == GlobalFiModInstNr[1]) || (9495 == GlobalFiModInstNr[2]) || (9495 == GlobalFiModInstNr[3]))));
	Tile mesh_3_29(
		.clock(clock),
		.io_in_a_0(r_125_0),
		.io_in_b_0(b_931_0),
		.io_in_d_0(b_1955_0),
		.io_in_control_0_dataflow(mesh_3_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2979_0),
		.io_in_last_0(r_4003_0),
		.io_in_valid_0(r_1955_0),
		.io_out_a_0(_mesh_3_29_io_out_a_0),
		.io_out_c_0(_mesh_3_29_io_out_c_0),
		.io_out_b_0(_mesh_3_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_29_io_out_id_0),
		.io_out_last_0(_mesh_3_29_io_out_last_0),
		.io_out_valid_0(_mesh_3_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9496 == GlobalFiModInstNr[0]) || (9496 == GlobalFiModInstNr[1]) || (9496 == GlobalFiModInstNr[2]) || (9496 == GlobalFiModInstNr[3]))));
	Tile mesh_3_30(
		.clock(clock),
		.io_in_a_0(r_126_0),
		.io_in_b_0(b_963_0),
		.io_in_d_0(b_1987_0),
		.io_in_control_0_dataflow(mesh_3_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3011_0),
		.io_in_last_0(r_4035_0),
		.io_in_valid_0(r_1987_0),
		.io_out_a_0(_mesh_3_30_io_out_a_0),
		.io_out_c_0(_mesh_3_30_io_out_c_0),
		.io_out_b_0(_mesh_3_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_30_io_out_id_0),
		.io_out_last_0(_mesh_3_30_io_out_last_0),
		.io_out_valid_0(_mesh_3_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9497 == GlobalFiModInstNr[0]) || (9497 == GlobalFiModInstNr[1]) || (9497 == GlobalFiModInstNr[2]) || (9497 == GlobalFiModInstNr[3]))));
	Tile mesh_3_31(
		.clock(clock),
		.io_in_a_0(r_127_0),
		.io_in_b_0(b_995_0),
		.io_in_d_0(b_2019_0),
		.io_in_control_0_dataflow(mesh_3_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3043_0),
		.io_in_last_0(r_4067_0),
		.io_in_valid_0(r_2019_0),
		.io_out_a_0(_mesh_3_31_io_out_a_0),
		.io_out_c_0(_mesh_3_31_io_out_c_0),
		.io_out_b_0(_mesh_3_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_31_io_out_id_0),
		.io_out_last_0(_mesh_3_31_io_out_last_0),
		.io_out_valid_0(_mesh_3_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9498 == GlobalFiModInstNr[0]) || (9498 == GlobalFiModInstNr[1]) || (9498 == GlobalFiModInstNr[2]) || (9498 == GlobalFiModInstNr[3]))));
	Tile mesh_4_0(
		.clock(clock),
		.io_in_a_0(r_128_0),
		.io_in_b_0(b_4_0),
		.io_in_d_0(b_1028_0),
		.io_in_control_0_dataflow(mesh_4_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2052_0),
		.io_in_last_0(r_3076_0),
		.io_in_valid_0(r_1028_0),
		.io_out_a_0(_mesh_4_0_io_out_a_0),
		.io_out_c_0(_mesh_4_0_io_out_c_0),
		.io_out_b_0(_mesh_4_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_0_io_out_id_0),
		.io_out_last_0(_mesh_4_0_io_out_last_0),
		.io_out_valid_0(_mesh_4_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9499 == GlobalFiModInstNr[0]) || (9499 == GlobalFiModInstNr[1]) || (9499 == GlobalFiModInstNr[2]) || (9499 == GlobalFiModInstNr[3]))));
	Tile mesh_4_1(
		.clock(clock),
		.io_in_a_0(r_129_0),
		.io_in_b_0(b_36_0),
		.io_in_d_0(b_1060_0),
		.io_in_control_0_dataflow(mesh_4_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2084_0),
		.io_in_last_0(r_3108_0),
		.io_in_valid_0(r_1060_0),
		.io_out_a_0(_mesh_4_1_io_out_a_0),
		.io_out_c_0(_mesh_4_1_io_out_c_0),
		.io_out_b_0(_mesh_4_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_1_io_out_id_0),
		.io_out_last_0(_mesh_4_1_io_out_last_0),
		.io_out_valid_0(_mesh_4_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9500 == GlobalFiModInstNr[0]) || (9500 == GlobalFiModInstNr[1]) || (9500 == GlobalFiModInstNr[2]) || (9500 == GlobalFiModInstNr[3]))));
	Tile mesh_4_2(
		.clock(clock),
		.io_in_a_0(r_130_0),
		.io_in_b_0(b_68_0),
		.io_in_d_0(b_1092_0),
		.io_in_control_0_dataflow(mesh_4_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2116_0),
		.io_in_last_0(r_3140_0),
		.io_in_valid_0(r_1092_0),
		.io_out_a_0(_mesh_4_2_io_out_a_0),
		.io_out_c_0(_mesh_4_2_io_out_c_0),
		.io_out_b_0(_mesh_4_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_2_io_out_id_0),
		.io_out_last_0(_mesh_4_2_io_out_last_0),
		.io_out_valid_0(_mesh_4_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9501 == GlobalFiModInstNr[0]) || (9501 == GlobalFiModInstNr[1]) || (9501 == GlobalFiModInstNr[2]) || (9501 == GlobalFiModInstNr[3]))));
	Tile mesh_4_3(
		.clock(clock),
		.io_in_a_0(r_131_0),
		.io_in_b_0(b_100_0),
		.io_in_d_0(b_1124_0),
		.io_in_control_0_dataflow(mesh_4_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2148_0),
		.io_in_last_0(r_3172_0),
		.io_in_valid_0(r_1124_0),
		.io_out_a_0(_mesh_4_3_io_out_a_0),
		.io_out_c_0(_mesh_4_3_io_out_c_0),
		.io_out_b_0(_mesh_4_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_3_io_out_id_0),
		.io_out_last_0(_mesh_4_3_io_out_last_0),
		.io_out_valid_0(_mesh_4_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9502 == GlobalFiModInstNr[0]) || (9502 == GlobalFiModInstNr[1]) || (9502 == GlobalFiModInstNr[2]) || (9502 == GlobalFiModInstNr[3]))));
	Tile mesh_4_4(
		.clock(clock),
		.io_in_a_0(r_132_0),
		.io_in_b_0(b_132_0),
		.io_in_d_0(b_1156_0),
		.io_in_control_0_dataflow(mesh_4_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2180_0),
		.io_in_last_0(r_3204_0),
		.io_in_valid_0(r_1156_0),
		.io_out_a_0(_mesh_4_4_io_out_a_0),
		.io_out_c_0(_mesh_4_4_io_out_c_0),
		.io_out_b_0(_mesh_4_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_4_io_out_id_0),
		.io_out_last_0(_mesh_4_4_io_out_last_0),
		.io_out_valid_0(_mesh_4_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9503 == GlobalFiModInstNr[0]) || (9503 == GlobalFiModInstNr[1]) || (9503 == GlobalFiModInstNr[2]) || (9503 == GlobalFiModInstNr[3]))));
	Tile mesh_4_5(
		.clock(clock),
		.io_in_a_0(r_133_0),
		.io_in_b_0(b_164_0),
		.io_in_d_0(b_1188_0),
		.io_in_control_0_dataflow(mesh_4_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2212_0),
		.io_in_last_0(r_3236_0),
		.io_in_valid_0(r_1188_0),
		.io_out_a_0(_mesh_4_5_io_out_a_0),
		.io_out_c_0(_mesh_4_5_io_out_c_0),
		.io_out_b_0(_mesh_4_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_5_io_out_id_0),
		.io_out_last_0(_mesh_4_5_io_out_last_0),
		.io_out_valid_0(_mesh_4_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9504 == GlobalFiModInstNr[0]) || (9504 == GlobalFiModInstNr[1]) || (9504 == GlobalFiModInstNr[2]) || (9504 == GlobalFiModInstNr[3]))));
	Tile mesh_4_6(
		.clock(clock),
		.io_in_a_0(r_134_0),
		.io_in_b_0(b_196_0),
		.io_in_d_0(b_1220_0),
		.io_in_control_0_dataflow(mesh_4_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2244_0),
		.io_in_last_0(r_3268_0),
		.io_in_valid_0(r_1220_0),
		.io_out_a_0(_mesh_4_6_io_out_a_0),
		.io_out_c_0(_mesh_4_6_io_out_c_0),
		.io_out_b_0(_mesh_4_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_6_io_out_id_0),
		.io_out_last_0(_mesh_4_6_io_out_last_0),
		.io_out_valid_0(_mesh_4_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9505 == GlobalFiModInstNr[0]) || (9505 == GlobalFiModInstNr[1]) || (9505 == GlobalFiModInstNr[2]) || (9505 == GlobalFiModInstNr[3]))));
	Tile mesh_4_7(
		.clock(clock),
		.io_in_a_0(r_135_0),
		.io_in_b_0(b_228_0),
		.io_in_d_0(b_1252_0),
		.io_in_control_0_dataflow(mesh_4_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2276_0),
		.io_in_last_0(r_3300_0),
		.io_in_valid_0(r_1252_0),
		.io_out_a_0(_mesh_4_7_io_out_a_0),
		.io_out_c_0(_mesh_4_7_io_out_c_0),
		.io_out_b_0(_mesh_4_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_7_io_out_id_0),
		.io_out_last_0(_mesh_4_7_io_out_last_0),
		.io_out_valid_0(_mesh_4_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9506 == GlobalFiModInstNr[0]) || (9506 == GlobalFiModInstNr[1]) || (9506 == GlobalFiModInstNr[2]) || (9506 == GlobalFiModInstNr[3]))));
	Tile mesh_4_8(
		.clock(clock),
		.io_in_a_0(r_136_0),
		.io_in_b_0(b_260_0),
		.io_in_d_0(b_1284_0),
		.io_in_control_0_dataflow(mesh_4_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2308_0),
		.io_in_last_0(r_3332_0),
		.io_in_valid_0(r_1284_0),
		.io_out_a_0(_mesh_4_8_io_out_a_0),
		.io_out_c_0(_mesh_4_8_io_out_c_0),
		.io_out_b_0(_mesh_4_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_8_io_out_id_0),
		.io_out_last_0(_mesh_4_8_io_out_last_0),
		.io_out_valid_0(_mesh_4_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9507 == GlobalFiModInstNr[0]) || (9507 == GlobalFiModInstNr[1]) || (9507 == GlobalFiModInstNr[2]) || (9507 == GlobalFiModInstNr[3]))));
	Tile mesh_4_9(
		.clock(clock),
		.io_in_a_0(r_137_0),
		.io_in_b_0(b_292_0),
		.io_in_d_0(b_1316_0),
		.io_in_control_0_dataflow(mesh_4_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2340_0),
		.io_in_last_0(r_3364_0),
		.io_in_valid_0(r_1316_0),
		.io_out_a_0(_mesh_4_9_io_out_a_0),
		.io_out_c_0(_mesh_4_9_io_out_c_0),
		.io_out_b_0(_mesh_4_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_9_io_out_id_0),
		.io_out_last_0(_mesh_4_9_io_out_last_0),
		.io_out_valid_0(_mesh_4_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9508 == GlobalFiModInstNr[0]) || (9508 == GlobalFiModInstNr[1]) || (9508 == GlobalFiModInstNr[2]) || (9508 == GlobalFiModInstNr[3]))));
	Tile mesh_4_10(
		.clock(clock),
		.io_in_a_0(r_138_0),
		.io_in_b_0(b_324_0),
		.io_in_d_0(b_1348_0),
		.io_in_control_0_dataflow(mesh_4_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2372_0),
		.io_in_last_0(r_3396_0),
		.io_in_valid_0(r_1348_0),
		.io_out_a_0(_mesh_4_10_io_out_a_0),
		.io_out_c_0(_mesh_4_10_io_out_c_0),
		.io_out_b_0(_mesh_4_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_10_io_out_id_0),
		.io_out_last_0(_mesh_4_10_io_out_last_0),
		.io_out_valid_0(_mesh_4_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9509 == GlobalFiModInstNr[0]) || (9509 == GlobalFiModInstNr[1]) || (9509 == GlobalFiModInstNr[2]) || (9509 == GlobalFiModInstNr[3]))));
	Tile mesh_4_11(
		.clock(clock),
		.io_in_a_0(r_139_0),
		.io_in_b_0(b_356_0),
		.io_in_d_0(b_1380_0),
		.io_in_control_0_dataflow(mesh_4_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2404_0),
		.io_in_last_0(r_3428_0),
		.io_in_valid_0(r_1380_0),
		.io_out_a_0(_mesh_4_11_io_out_a_0),
		.io_out_c_0(_mesh_4_11_io_out_c_0),
		.io_out_b_0(_mesh_4_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_11_io_out_id_0),
		.io_out_last_0(_mesh_4_11_io_out_last_0),
		.io_out_valid_0(_mesh_4_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9510 == GlobalFiModInstNr[0]) || (9510 == GlobalFiModInstNr[1]) || (9510 == GlobalFiModInstNr[2]) || (9510 == GlobalFiModInstNr[3]))));
	Tile mesh_4_12(
		.clock(clock),
		.io_in_a_0(r_140_0),
		.io_in_b_0(b_388_0),
		.io_in_d_0(b_1412_0),
		.io_in_control_0_dataflow(mesh_4_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2436_0),
		.io_in_last_0(r_3460_0),
		.io_in_valid_0(r_1412_0),
		.io_out_a_0(_mesh_4_12_io_out_a_0),
		.io_out_c_0(_mesh_4_12_io_out_c_0),
		.io_out_b_0(_mesh_4_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_12_io_out_id_0),
		.io_out_last_0(_mesh_4_12_io_out_last_0),
		.io_out_valid_0(_mesh_4_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9511 == GlobalFiModInstNr[0]) || (9511 == GlobalFiModInstNr[1]) || (9511 == GlobalFiModInstNr[2]) || (9511 == GlobalFiModInstNr[3]))));
	Tile mesh_4_13(
		.clock(clock),
		.io_in_a_0(r_141_0),
		.io_in_b_0(b_420_0),
		.io_in_d_0(b_1444_0),
		.io_in_control_0_dataflow(mesh_4_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2468_0),
		.io_in_last_0(r_3492_0),
		.io_in_valid_0(r_1444_0),
		.io_out_a_0(_mesh_4_13_io_out_a_0),
		.io_out_c_0(_mesh_4_13_io_out_c_0),
		.io_out_b_0(_mesh_4_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_13_io_out_id_0),
		.io_out_last_0(_mesh_4_13_io_out_last_0),
		.io_out_valid_0(_mesh_4_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9512 == GlobalFiModInstNr[0]) || (9512 == GlobalFiModInstNr[1]) || (9512 == GlobalFiModInstNr[2]) || (9512 == GlobalFiModInstNr[3]))));
	Tile mesh_4_14(
		.clock(clock),
		.io_in_a_0(r_142_0),
		.io_in_b_0(b_452_0),
		.io_in_d_0(b_1476_0),
		.io_in_control_0_dataflow(mesh_4_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2500_0),
		.io_in_last_0(r_3524_0),
		.io_in_valid_0(r_1476_0),
		.io_out_a_0(_mesh_4_14_io_out_a_0),
		.io_out_c_0(_mesh_4_14_io_out_c_0),
		.io_out_b_0(_mesh_4_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_14_io_out_id_0),
		.io_out_last_0(_mesh_4_14_io_out_last_0),
		.io_out_valid_0(_mesh_4_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9513 == GlobalFiModInstNr[0]) || (9513 == GlobalFiModInstNr[1]) || (9513 == GlobalFiModInstNr[2]) || (9513 == GlobalFiModInstNr[3]))));
	Tile mesh_4_15(
		.clock(clock),
		.io_in_a_0(r_143_0),
		.io_in_b_0(b_484_0),
		.io_in_d_0(b_1508_0),
		.io_in_control_0_dataflow(mesh_4_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2532_0),
		.io_in_last_0(r_3556_0),
		.io_in_valid_0(r_1508_0),
		.io_out_a_0(_mesh_4_15_io_out_a_0),
		.io_out_c_0(_mesh_4_15_io_out_c_0),
		.io_out_b_0(_mesh_4_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_15_io_out_id_0),
		.io_out_last_0(_mesh_4_15_io_out_last_0),
		.io_out_valid_0(_mesh_4_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9514 == GlobalFiModInstNr[0]) || (9514 == GlobalFiModInstNr[1]) || (9514 == GlobalFiModInstNr[2]) || (9514 == GlobalFiModInstNr[3]))));
	Tile mesh_4_16(
		.clock(clock),
		.io_in_a_0(r_144_0),
		.io_in_b_0(b_516_0),
		.io_in_d_0(b_1540_0),
		.io_in_control_0_dataflow(mesh_4_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2564_0),
		.io_in_last_0(r_3588_0),
		.io_in_valid_0(r_1540_0),
		.io_out_a_0(_mesh_4_16_io_out_a_0),
		.io_out_c_0(_mesh_4_16_io_out_c_0),
		.io_out_b_0(_mesh_4_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_16_io_out_id_0),
		.io_out_last_0(_mesh_4_16_io_out_last_0),
		.io_out_valid_0(_mesh_4_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9515 == GlobalFiModInstNr[0]) || (9515 == GlobalFiModInstNr[1]) || (9515 == GlobalFiModInstNr[2]) || (9515 == GlobalFiModInstNr[3]))));
	Tile mesh_4_17(
		.clock(clock),
		.io_in_a_0(r_145_0),
		.io_in_b_0(b_548_0),
		.io_in_d_0(b_1572_0),
		.io_in_control_0_dataflow(mesh_4_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2596_0),
		.io_in_last_0(r_3620_0),
		.io_in_valid_0(r_1572_0),
		.io_out_a_0(_mesh_4_17_io_out_a_0),
		.io_out_c_0(_mesh_4_17_io_out_c_0),
		.io_out_b_0(_mesh_4_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_17_io_out_id_0),
		.io_out_last_0(_mesh_4_17_io_out_last_0),
		.io_out_valid_0(_mesh_4_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9516 == GlobalFiModInstNr[0]) || (9516 == GlobalFiModInstNr[1]) || (9516 == GlobalFiModInstNr[2]) || (9516 == GlobalFiModInstNr[3]))));
	Tile mesh_4_18(
		.clock(clock),
		.io_in_a_0(r_146_0),
		.io_in_b_0(b_580_0),
		.io_in_d_0(b_1604_0),
		.io_in_control_0_dataflow(mesh_4_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2628_0),
		.io_in_last_0(r_3652_0),
		.io_in_valid_0(r_1604_0),
		.io_out_a_0(_mesh_4_18_io_out_a_0),
		.io_out_c_0(_mesh_4_18_io_out_c_0),
		.io_out_b_0(_mesh_4_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_18_io_out_id_0),
		.io_out_last_0(_mesh_4_18_io_out_last_0),
		.io_out_valid_0(_mesh_4_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9517 == GlobalFiModInstNr[0]) || (9517 == GlobalFiModInstNr[1]) || (9517 == GlobalFiModInstNr[2]) || (9517 == GlobalFiModInstNr[3]))));
	Tile mesh_4_19(
		.clock(clock),
		.io_in_a_0(r_147_0),
		.io_in_b_0(b_612_0),
		.io_in_d_0(b_1636_0),
		.io_in_control_0_dataflow(mesh_4_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2660_0),
		.io_in_last_0(r_3684_0),
		.io_in_valid_0(r_1636_0),
		.io_out_a_0(_mesh_4_19_io_out_a_0),
		.io_out_c_0(_mesh_4_19_io_out_c_0),
		.io_out_b_0(_mesh_4_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_19_io_out_id_0),
		.io_out_last_0(_mesh_4_19_io_out_last_0),
		.io_out_valid_0(_mesh_4_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9518 == GlobalFiModInstNr[0]) || (9518 == GlobalFiModInstNr[1]) || (9518 == GlobalFiModInstNr[2]) || (9518 == GlobalFiModInstNr[3]))));
	Tile mesh_4_20(
		.clock(clock),
		.io_in_a_0(r_148_0),
		.io_in_b_0(b_644_0),
		.io_in_d_0(b_1668_0),
		.io_in_control_0_dataflow(mesh_4_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2692_0),
		.io_in_last_0(r_3716_0),
		.io_in_valid_0(r_1668_0),
		.io_out_a_0(_mesh_4_20_io_out_a_0),
		.io_out_c_0(_mesh_4_20_io_out_c_0),
		.io_out_b_0(_mesh_4_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_20_io_out_id_0),
		.io_out_last_0(_mesh_4_20_io_out_last_0),
		.io_out_valid_0(_mesh_4_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9519 == GlobalFiModInstNr[0]) || (9519 == GlobalFiModInstNr[1]) || (9519 == GlobalFiModInstNr[2]) || (9519 == GlobalFiModInstNr[3]))));
	Tile mesh_4_21(
		.clock(clock),
		.io_in_a_0(r_149_0),
		.io_in_b_0(b_676_0),
		.io_in_d_0(b_1700_0),
		.io_in_control_0_dataflow(mesh_4_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2724_0),
		.io_in_last_0(r_3748_0),
		.io_in_valid_0(r_1700_0),
		.io_out_a_0(_mesh_4_21_io_out_a_0),
		.io_out_c_0(_mesh_4_21_io_out_c_0),
		.io_out_b_0(_mesh_4_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_21_io_out_id_0),
		.io_out_last_0(_mesh_4_21_io_out_last_0),
		.io_out_valid_0(_mesh_4_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9520 == GlobalFiModInstNr[0]) || (9520 == GlobalFiModInstNr[1]) || (9520 == GlobalFiModInstNr[2]) || (9520 == GlobalFiModInstNr[3]))));
	Tile mesh_4_22(
		.clock(clock),
		.io_in_a_0(r_150_0),
		.io_in_b_0(b_708_0),
		.io_in_d_0(b_1732_0),
		.io_in_control_0_dataflow(mesh_4_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2756_0),
		.io_in_last_0(r_3780_0),
		.io_in_valid_0(r_1732_0),
		.io_out_a_0(_mesh_4_22_io_out_a_0),
		.io_out_c_0(_mesh_4_22_io_out_c_0),
		.io_out_b_0(_mesh_4_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_22_io_out_id_0),
		.io_out_last_0(_mesh_4_22_io_out_last_0),
		.io_out_valid_0(_mesh_4_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9521 == GlobalFiModInstNr[0]) || (9521 == GlobalFiModInstNr[1]) || (9521 == GlobalFiModInstNr[2]) || (9521 == GlobalFiModInstNr[3]))));
	Tile mesh_4_23(
		.clock(clock),
		.io_in_a_0(r_151_0),
		.io_in_b_0(b_740_0),
		.io_in_d_0(b_1764_0),
		.io_in_control_0_dataflow(mesh_4_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2788_0),
		.io_in_last_0(r_3812_0),
		.io_in_valid_0(r_1764_0),
		.io_out_a_0(_mesh_4_23_io_out_a_0),
		.io_out_c_0(_mesh_4_23_io_out_c_0),
		.io_out_b_0(_mesh_4_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_23_io_out_id_0),
		.io_out_last_0(_mesh_4_23_io_out_last_0),
		.io_out_valid_0(_mesh_4_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9522 == GlobalFiModInstNr[0]) || (9522 == GlobalFiModInstNr[1]) || (9522 == GlobalFiModInstNr[2]) || (9522 == GlobalFiModInstNr[3]))));
	Tile mesh_4_24(
		.clock(clock),
		.io_in_a_0(r_152_0),
		.io_in_b_0(b_772_0),
		.io_in_d_0(b_1796_0),
		.io_in_control_0_dataflow(mesh_4_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2820_0),
		.io_in_last_0(r_3844_0),
		.io_in_valid_0(r_1796_0),
		.io_out_a_0(_mesh_4_24_io_out_a_0),
		.io_out_c_0(_mesh_4_24_io_out_c_0),
		.io_out_b_0(_mesh_4_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_24_io_out_id_0),
		.io_out_last_0(_mesh_4_24_io_out_last_0),
		.io_out_valid_0(_mesh_4_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9523 == GlobalFiModInstNr[0]) || (9523 == GlobalFiModInstNr[1]) || (9523 == GlobalFiModInstNr[2]) || (9523 == GlobalFiModInstNr[3]))));
	Tile mesh_4_25(
		.clock(clock),
		.io_in_a_0(r_153_0),
		.io_in_b_0(b_804_0),
		.io_in_d_0(b_1828_0),
		.io_in_control_0_dataflow(mesh_4_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2852_0),
		.io_in_last_0(r_3876_0),
		.io_in_valid_0(r_1828_0),
		.io_out_a_0(_mesh_4_25_io_out_a_0),
		.io_out_c_0(_mesh_4_25_io_out_c_0),
		.io_out_b_0(_mesh_4_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_25_io_out_id_0),
		.io_out_last_0(_mesh_4_25_io_out_last_0),
		.io_out_valid_0(_mesh_4_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9524 == GlobalFiModInstNr[0]) || (9524 == GlobalFiModInstNr[1]) || (9524 == GlobalFiModInstNr[2]) || (9524 == GlobalFiModInstNr[3]))));
	Tile mesh_4_26(
		.clock(clock),
		.io_in_a_0(r_154_0),
		.io_in_b_0(b_836_0),
		.io_in_d_0(b_1860_0),
		.io_in_control_0_dataflow(mesh_4_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2884_0),
		.io_in_last_0(r_3908_0),
		.io_in_valid_0(r_1860_0),
		.io_out_a_0(_mesh_4_26_io_out_a_0),
		.io_out_c_0(_mesh_4_26_io_out_c_0),
		.io_out_b_0(_mesh_4_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_26_io_out_id_0),
		.io_out_last_0(_mesh_4_26_io_out_last_0),
		.io_out_valid_0(_mesh_4_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9525 == GlobalFiModInstNr[0]) || (9525 == GlobalFiModInstNr[1]) || (9525 == GlobalFiModInstNr[2]) || (9525 == GlobalFiModInstNr[3]))));
	Tile mesh_4_27(
		.clock(clock),
		.io_in_a_0(r_155_0),
		.io_in_b_0(b_868_0),
		.io_in_d_0(b_1892_0),
		.io_in_control_0_dataflow(mesh_4_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2916_0),
		.io_in_last_0(r_3940_0),
		.io_in_valid_0(r_1892_0),
		.io_out_a_0(_mesh_4_27_io_out_a_0),
		.io_out_c_0(_mesh_4_27_io_out_c_0),
		.io_out_b_0(_mesh_4_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_27_io_out_id_0),
		.io_out_last_0(_mesh_4_27_io_out_last_0),
		.io_out_valid_0(_mesh_4_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9526 == GlobalFiModInstNr[0]) || (9526 == GlobalFiModInstNr[1]) || (9526 == GlobalFiModInstNr[2]) || (9526 == GlobalFiModInstNr[3]))));
	Tile mesh_4_28(
		.clock(clock),
		.io_in_a_0(r_156_0),
		.io_in_b_0(b_900_0),
		.io_in_d_0(b_1924_0),
		.io_in_control_0_dataflow(mesh_4_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2948_0),
		.io_in_last_0(r_3972_0),
		.io_in_valid_0(r_1924_0),
		.io_out_a_0(_mesh_4_28_io_out_a_0),
		.io_out_c_0(_mesh_4_28_io_out_c_0),
		.io_out_b_0(_mesh_4_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_28_io_out_id_0),
		.io_out_last_0(_mesh_4_28_io_out_last_0),
		.io_out_valid_0(_mesh_4_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9527 == GlobalFiModInstNr[0]) || (9527 == GlobalFiModInstNr[1]) || (9527 == GlobalFiModInstNr[2]) || (9527 == GlobalFiModInstNr[3]))));
	Tile mesh_4_29(
		.clock(clock),
		.io_in_a_0(r_157_0),
		.io_in_b_0(b_932_0),
		.io_in_d_0(b_1956_0),
		.io_in_control_0_dataflow(mesh_4_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2980_0),
		.io_in_last_0(r_4004_0),
		.io_in_valid_0(r_1956_0),
		.io_out_a_0(_mesh_4_29_io_out_a_0),
		.io_out_c_0(_mesh_4_29_io_out_c_0),
		.io_out_b_0(_mesh_4_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_29_io_out_id_0),
		.io_out_last_0(_mesh_4_29_io_out_last_0),
		.io_out_valid_0(_mesh_4_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9528 == GlobalFiModInstNr[0]) || (9528 == GlobalFiModInstNr[1]) || (9528 == GlobalFiModInstNr[2]) || (9528 == GlobalFiModInstNr[3]))));
	Tile mesh_4_30(
		.clock(clock),
		.io_in_a_0(r_158_0),
		.io_in_b_0(b_964_0),
		.io_in_d_0(b_1988_0),
		.io_in_control_0_dataflow(mesh_4_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3012_0),
		.io_in_last_0(r_4036_0),
		.io_in_valid_0(r_1988_0),
		.io_out_a_0(_mesh_4_30_io_out_a_0),
		.io_out_c_0(_mesh_4_30_io_out_c_0),
		.io_out_b_0(_mesh_4_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_30_io_out_id_0),
		.io_out_last_0(_mesh_4_30_io_out_last_0),
		.io_out_valid_0(_mesh_4_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9529 == GlobalFiModInstNr[0]) || (9529 == GlobalFiModInstNr[1]) || (9529 == GlobalFiModInstNr[2]) || (9529 == GlobalFiModInstNr[3]))));
	Tile mesh_4_31(
		.clock(clock),
		.io_in_a_0(r_159_0),
		.io_in_b_0(b_996_0),
		.io_in_d_0(b_2020_0),
		.io_in_control_0_dataflow(mesh_4_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3044_0),
		.io_in_last_0(r_4068_0),
		.io_in_valid_0(r_2020_0),
		.io_out_a_0(_mesh_4_31_io_out_a_0),
		.io_out_c_0(_mesh_4_31_io_out_c_0),
		.io_out_b_0(_mesh_4_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_31_io_out_id_0),
		.io_out_last_0(_mesh_4_31_io_out_last_0),
		.io_out_valid_0(_mesh_4_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9530 == GlobalFiModInstNr[0]) || (9530 == GlobalFiModInstNr[1]) || (9530 == GlobalFiModInstNr[2]) || (9530 == GlobalFiModInstNr[3]))));
	Tile mesh_5_0(
		.clock(clock),
		.io_in_a_0(r_160_0),
		.io_in_b_0(b_5_0),
		.io_in_d_0(b_1029_0),
		.io_in_control_0_dataflow(mesh_5_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2053_0),
		.io_in_last_0(r_3077_0),
		.io_in_valid_0(r_1029_0),
		.io_out_a_0(_mesh_5_0_io_out_a_0),
		.io_out_c_0(_mesh_5_0_io_out_c_0),
		.io_out_b_0(_mesh_5_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_0_io_out_id_0),
		.io_out_last_0(_mesh_5_0_io_out_last_0),
		.io_out_valid_0(_mesh_5_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9531 == GlobalFiModInstNr[0]) || (9531 == GlobalFiModInstNr[1]) || (9531 == GlobalFiModInstNr[2]) || (9531 == GlobalFiModInstNr[3]))));
	Tile mesh_5_1(
		.clock(clock),
		.io_in_a_0(r_161_0),
		.io_in_b_0(b_37_0),
		.io_in_d_0(b_1061_0),
		.io_in_control_0_dataflow(mesh_5_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2085_0),
		.io_in_last_0(r_3109_0),
		.io_in_valid_0(r_1061_0),
		.io_out_a_0(_mesh_5_1_io_out_a_0),
		.io_out_c_0(_mesh_5_1_io_out_c_0),
		.io_out_b_0(_mesh_5_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_1_io_out_id_0),
		.io_out_last_0(_mesh_5_1_io_out_last_0),
		.io_out_valid_0(_mesh_5_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9532 == GlobalFiModInstNr[0]) || (9532 == GlobalFiModInstNr[1]) || (9532 == GlobalFiModInstNr[2]) || (9532 == GlobalFiModInstNr[3]))));
	Tile mesh_5_2(
		.clock(clock),
		.io_in_a_0(r_162_0),
		.io_in_b_0(b_69_0),
		.io_in_d_0(b_1093_0),
		.io_in_control_0_dataflow(mesh_5_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2117_0),
		.io_in_last_0(r_3141_0),
		.io_in_valid_0(r_1093_0),
		.io_out_a_0(_mesh_5_2_io_out_a_0),
		.io_out_c_0(_mesh_5_2_io_out_c_0),
		.io_out_b_0(_mesh_5_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_2_io_out_id_0),
		.io_out_last_0(_mesh_5_2_io_out_last_0),
		.io_out_valid_0(_mesh_5_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9533 == GlobalFiModInstNr[0]) || (9533 == GlobalFiModInstNr[1]) || (9533 == GlobalFiModInstNr[2]) || (9533 == GlobalFiModInstNr[3]))));
	Tile mesh_5_3(
		.clock(clock),
		.io_in_a_0(r_163_0),
		.io_in_b_0(b_101_0),
		.io_in_d_0(b_1125_0),
		.io_in_control_0_dataflow(mesh_5_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2149_0),
		.io_in_last_0(r_3173_0),
		.io_in_valid_0(r_1125_0),
		.io_out_a_0(_mesh_5_3_io_out_a_0),
		.io_out_c_0(_mesh_5_3_io_out_c_0),
		.io_out_b_0(_mesh_5_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_3_io_out_id_0),
		.io_out_last_0(_mesh_5_3_io_out_last_0),
		.io_out_valid_0(_mesh_5_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9534 == GlobalFiModInstNr[0]) || (9534 == GlobalFiModInstNr[1]) || (9534 == GlobalFiModInstNr[2]) || (9534 == GlobalFiModInstNr[3]))));
	Tile mesh_5_4(
		.clock(clock),
		.io_in_a_0(r_164_0),
		.io_in_b_0(b_133_0),
		.io_in_d_0(b_1157_0),
		.io_in_control_0_dataflow(mesh_5_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2181_0),
		.io_in_last_0(r_3205_0),
		.io_in_valid_0(r_1157_0),
		.io_out_a_0(_mesh_5_4_io_out_a_0),
		.io_out_c_0(_mesh_5_4_io_out_c_0),
		.io_out_b_0(_mesh_5_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_4_io_out_id_0),
		.io_out_last_0(_mesh_5_4_io_out_last_0),
		.io_out_valid_0(_mesh_5_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9535 == GlobalFiModInstNr[0]) || (9535 == GlobalFiModInstNr[1]) || (9535 == GlobalFiModInstNr[2]) || (9535 == GlobalFiModInstNr[3]))));
	Tile mesh_5_5(
		.clock(clock),
		.io_in_a_0(r_165_0),
		.io_in_b_0(b_165_0),
		.io_in_d_0(b_1189_0),
		.io_in_control_0_dataflow(mesh_5_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2213_0),
		.io_in_last_0(r_3237_0),
		.io_in_valid_0(r_1189_0),
		.io_out_a_0(_mesh_5_5_io_out_a_0),
		.io_out_c_0(_mesh_5_5_io_out_c_0),
		.io_out_b_0(_mesh_5_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_5_io_out_id_0),
		.io_out_last_0(_mesh_5_5_io_out_last_0),
		.io_out_valid_0(_mesh_5_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9536 == GlobalFiModInstNr[0]) || (9536 == GlobalFiModInstNr[1]) || (9536 == GlobalFiModInstNr[2]) || (9536 == GlobalFiModInstNr[3]))));
	Tile mesh_5_6(
		.clock(clock),
		.io_in_a_0(r_166_0),
		.io_in_b_0(b_197_0),
		.io_in_d_0(b_1221_0),
		.io_in_control_0_dataflow(mesh_5_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2245_0),
		.io_in_last_0(r_3269_0),
		.io_in_valid_0(r_1221_0),
		.io_out_a_0(_mesh_5_6_io_out_a_0),
		.io_out_c_0(_mesh_5_6_io_out_c_0),
		.io_out_b_0(_mesh_5_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_6_io_out_id_0),
		.io_out_last_0(_mesh_5_6_io_out_last_0),
		.io_out_valid_0(_mesh_5_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9537 == GlobalFiModInstNr[0]) || (9537 == GlobalFiModInstNr[1]) || (9537 == GlobalFiModInstNr[2]) || (9537 == GlobalFiModInstNr[3]))));
	Tile mesh_5_7(
		.clock(clock),
		.io_in_a_0(r_167_0),
		.io_in_b_0(b_229_0),
		.io_in_d_0(b_1253_0),
		.io_in_control_0_dataflow(mesh_5_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2277_0),
		.io_in_last_0(r_3301_0),
		.io_in_valid_0(r_1253_0),
		.io_out_a_0(_mesh_5_7_io_out_a_0),
		.io_out_c_0(_mesh_5_7_io_out_c_0),
		.io_out_b_0(_mesh_5_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_7_io_out_id_0),
		.io_out_last_0(_mesh_5_7_io_out_last_0),
		.io_out_valid_0(_mesh_5_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9538 == GlobalFiModInstNr[0]) || (9538 == GlobalFiModInstNr[1]) || (9538 == GlobalFiModInstNr[2]) || (9538 == GlobalFiModInstNr[3]))));
	Tile mesh_5_8(
		.clock(clock),
		.io_in_a_0(r_168_0),
		.io_in_b_0(b_261_0),
		.io_in_d_0(b_1285_0),
		.io_in_control_0_dataflow(mesh_5_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2309_0),
		.io_in_last_0(r_3333_0),
		.io_in_valid_0(r_1285_0),
		.io_out_a_0(_mesh_5_8_io_out_a_0),
		.io_out_c_0(_mesh_5_8_io_out_c_0),
		.io_out_b_0(_mesh_5_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_8_io_out_id_0),
		.io_out_last_0(_mesh_5_8_io_out_last_0),
		.io_out_valid_0(_mesh_5_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9539 == GlobalFiModInstNr[0]) || (9539 == GlobalFiModInstNr[1]) || (9539 == GlobalFiModInstNr[2]) || (9539 == GlobalFiModInstNr[3]))));
	Tile mesh_5_9(
		.clock(clock),
		.io_in_a_0(r_169_0),
		.io_in_b_0(b_293_0),
		.io_in_d_0(b_1317_0),
		.io_in_control_0_dataflow(mesh_5_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2341_0),
		.io_in_last_0(r_3365_0),
		.io_in_valid_0(r_1317_0),
		.io_out_a_0(_mesh_5_9_io_out_a_0),
		.io_out_c_0(_mesh_5_9_io_out_c_0),
		.io_out_b_0(_mesh_5_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_9_io_out_id_0),
		.io_out_last_0(_mesh_5_9_io_out_last_0),
		.io_out_valid_0(_mesh_5_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9540 == GlobalFiModInstNr[0]) || (9540 == GlobalFiModInstNr[1]) || (9540 == GlobalFiModInstNr[2]) || (9540 == GlobalFiModInstNr[3]))));
	Tile mesh_5_10(
		.clock(clock),
		.io_in_a_0(r_170_0),
		.io_in_b_0(b_325_0),
		.io_in_d_0(b_1349_0),
		.io_in_control_0_dataflow(mesh_5_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2373_0),
		.io_in_last_0(r_3397_0),
		.io_in_valid_0(r_1349_0),
		.io_out_a_0(_mesh_5_10_io_out_a_0),
		.io_out_c_0(_mesh_5_10_io_out_c_0),
		.io_out_b_0(_mesh_5_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_10_io_out_id_0),
		.io_out_last_0(_mesh_5_10_io_out_last_0),
		.io_out_valid_0(_mesh_5_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9541 == GlobalFiModInstNr[0]) || (9541 == GlobalFiModInstNr[1]) || (9541 == GlobalFiModInstNr[2]) || (9541 == GlobalFiModInstNr[3]))));
	Tile mesh_5_11(
		.clock(clock),
		.io_in_a_0(r_171_0),
		.io_in_b_0(b_357_0),
		.io_in_d_0(b_1381_0),
		.io_in_control_0_dataflow(mesh_5_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2405_0),
		.io_in_last_0(r_3429_0),
		.io_in_valid_0(r_1381_0),
		.io_out_a_0(_mesh_5_11_io_out_a_0),
		.io_out_c_0(_mesh_5_11_io_out_c_0),
		.io_out_b_0(_mesh_5_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_11_io_out_id_0),
		.io_out_last_0(_mesh_5_11_io_out_last_0),
		.io_out_valid_0(_mesh_5_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9542 == GlobalFiModInstNr[0]) || (9542 == GlobalFiModInstNr[1]) || (9542 == GlobalFiModInstNr[2]) || (9542 == GlobalFiModInstNr[3]))));
	Tile mesh_5_12(
		.clock(clock),
		.io_in_a_0(r_172_0),
		.io_in_b_0(b_389_0),
		.io_in_d_0(b_1413_0),
		.io_in_control_0_dataflow(mesh_5_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2437_0),
		.io_in_last_0(r_3461_0),
		.io_in_valid_0(r_1413_0),
		.io_out_a_0(_mesh_5_12_io_out_a_0),
		.io_out_c_0(_mesh_5_12_io_out_c_0),
		.io_out_b_0(_mesh_5_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_12_io_out_id_0),
		.io_out_last_0(_mesh_5_12_io_out_last_0),
		.io_out_valid_0(_mesh_5_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9543 == GlobalFiModInstNr[0]) || (9543 == GlobalFiModInstNr[1]) || (9543 == GlobalFiModInstNr[2]) || (9543 == GlobalFiModInstNr[3]))));
	Tile mesh_5_13(
		.clock(clock),
		.io_in_a_0(r_173_0),
		.io_in_b_0(b_421_0),
		.io_in_d_0(b_1445_0),
		.io_in_control_0_dataflow(mesh_5_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2469_0),
		.io_in_last_0(r_3493_0),
		.io_in_valid_0(r_1445_0),
		.io_out_a_0(_mesh_5_13_io_out_a_0),
		.io_out_c_0(_mesh_5_13_io_out_c_0),
		.io_out_b_0(_mesh_5_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_13_io_out_id_0),
		.io_out_last_0(_mesh_5_13_io_out_last_0),
		.io_out_valid_0(_mesh_5_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9544 == GlobalFiModInstNr[0]) || (9544 == GlobalFiModInstNr[1]) || (9544 == GlobalFiModInstNr[2]) || (9544 == GlobalFiModInstNr[3]))));
	Tile mesh_5_14(
		.clock(clock),
		.io_in_a_0(r_174_0),
		.io_in_b_0(b_453_0),
		.io_in_d_0(b_1477_0),
		.io_in_control_0_dataflow(mesh_5_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2501_0),
		.io_in_last_0(r_3525_0),
		.io_in_valid_0(r_1477_0),
		.io_out_a_0(_mesh_5_14_io_out_a_0),
		.io_out_c_0(_mesh_5_14_io_out_c_0),
		.io_out_b_0(_mesh_5_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_14_io_out_id_0),
		.io_out_last_0(_mesh_5_14_io_out_last_0),
		.io_out_valid_0(_mesh_5_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9545 == GlobalFiModInstNr[0]) || (9545 == GlobalFiModInstNr[1]) || (9545 == GlobalFiModInstNr[2]) || (9545 == GlobalFiModInstNr[3]))));
	Tile mesh_5_15(
		.clock(clock),
		.io_in_a_0(r_175_0),
		.io_in_b_0(b_485_0),
		.io_in_d_0(b_1509_0),
		.io_in_control_0_dataflow(mesh_5_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2533_0),
		.io_in_last_0(r_3557_0),
		.io_in_valid_0(r_1509_0),
		.io_out_a_0(_mesh_5_15_io_out_a_0),
		.io_out_c_0(_mesh_5_15_io_out_c_0),
		.io_out_b_0(_mesh_5_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_15_io_out_id_0),
		.io_out_last_0(_mesh_5_15_io_out_last_0),
		.io_out_valid_0(_mesh_5_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9546 == GlobalFiModInstNr[0]) || (9546 == GlobalFiModInstNr[1]) || (9546 == GlobalFiModInstNr[2]) || (9546 == GlobalFiModInstNr[3]))));
	Tile mesh_5_16(
		.clock(clock),
		.io_in_a_0(r_176_0),
		.io_in_b_0(b_517_0),
		.io_in_d_0(b_1541_0),
		.io_in_control_0_dataflow(mesh_5_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2565_0),
		.io_in_last_0(r_3589_0),
		.io_in_valid_0(r_1541_0),
		.io_out_a_0(_mesh_5_16_io_out_a_0),
		.io_out_c_0(_mesh_5_16_io_out_c_0),
		.io_out_b_0(_mesh_5_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_16_io_out_id_0),
		.io_out_last_0(_mesh_5_16_io_out_last_0),
		.io_out_valid_0(_mesh_5_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9547 == GlobalFiModInstNr[0]) || (9547 == GlobalFiModInstNr[1]) || (9547 == GlobalFiModInstNr[2]) || (9547 == GlobalFiModInstNr[3]))));
	Tile mesh_5_17(
		.clock(clock),
		.io_in_a_0(r_177_0),
		.io_in_b_0(b_549_0),
		.io_in_d_0(b_1573_0),
		.io_in_control_0_dataflow(mesh_5_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2597_0),
		.io_in_last_0(r_3621_0),
		.io_in_valid_0(r_1573_0),
		.io_out_a_0(_mesh_5_17_io_out_a_0),
		.io_out_c_0(_mesh_5_17_io_out_c_0),
		.io_out_b_0(_mesh_5_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_17_io_out_id_0),
		.io_out_last_0(_mesh_5_17_io_out_last_0),
		.io_out_valid_0(_mesh_5_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9548 == GlobalFiModInstNr[0]) || (9548 == GlobalFiModInstNr[1]) || (9548 == GlobalFiModInstNr[2]) || (9548 == GlobalFiModInstNr[3]))));
	Tile mesh_5_18(
		.clock(clock),
		.io_in_a_0(r_178_0),
		.io_in_b_0(b_581_0),
		.io_in_d_0(b_1605_0),
		.io_in_control_0_dataflow(mesh_5_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2629_0),
		.io_in_last_0(r_3653_0),
		.io_in_valid_0(r_1605_0),
		.io_out_a_0(_mesh_5_18_io_out_a_0),
		.io_out_c_0(_mesh_5_18_io_out_c_0),
		.io_out_b_0(_mesh_5_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_18_io_out_id_0),
		.io_out_last_0(_mesh_5_18_io_out_last_0),
		.io_out_valid_0(_mesh_5_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9549 == GlobalFiModInstNr[0]) || (9549 == GlobalFiModInstNr[1]) || (9549 == GlobalFiModInstNr[2]) || (9549 == GlobalFiModInstNr[3]))));
	Tile mesh_5_19(
		.clock(clock),
		.io_in_a_0(r_179_0),
		.io_in_b_0(b_613_0),
		.io_in_d_0(b_1637_0),
		.io_in_control_0_dataflow(mesh_5_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2661_0),
		.io_in_last_0(r_3685_0),
		.io_in_valid_0(r_1637_0),
		.io_out_a_0(_mesh_5_19_io_out_a_0),
		.io_out_c_0(_mesh_5_19_io_out_c_0),
		.io_out_b_0(_mesh_5_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_19_io_out_id_0),
		.io_out_last_0(_mesh_5_19_io_out_last_0),
		.io_out_valid_0(_mesh_5_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9550 == GlobalFiModInstNr[0]) || (9550 == GlobalFiModInstNr[1]) || (9550 == GlobalFiModInstNr[2]) || (9550 == GlobalFiModInstNr[3]))));
	Tile mesh_5_20(
		.clock(clock),
		.io_in_a_0(r_180_0),
		.io_in_b_0(b_645_0),
		.io_in_d_0(b_1669_0),
		.io_in_control_0_dataflow(mesh_5_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2693_0),
		.io_in_last_0(r_3717_0),
		.io_in_valid_0(r_1669_0),
		.io_out_a_0(_mesh_5_20_io_out_a_0),
		.io_out_c_0(_mesh_5_20_io_out_c_0),
		.io_out_b_0(_mesh_5_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_20_io_out_id_0),
		.io_out_last_0(_mesh_5_20_io_out_last_0),
		.io_out_valid_0(_mesh_5_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9551 == GlobalFiModInstNr[0]) || (9551 == GlobalFiModInstNr[1]) || (9551 == GlobalFiModInstNr[2]) || (9551 == GlobalFiModInstNr[3]))));
	Tile mesh_5_21(
		.clock(clock),
		.io_in_a_0(r_181_0),
		.io_in_b_0(b_677_0),
		.io_in_d_0(b_1701_0),
		.io_in_control_0_dataflow(mesh_5_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2725_0),
		.io_in_last_0(r_3749_0),
		.io_in_valid_0(r_1701_0),
		.io_out_a_0(_mesh_5_21_io_out_a_0),
		.io_out_c_0(_mesh_5_21_io_out_c_0),
		.io_out_b_0(_mesh_5_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_21_io_out_id_0),
		.io_out_last_0(_mesh_5_21_io_out_last_0),
		.io_out_valid_0(_mesh_5_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9552 == GlobalFiModInstNr[0]) || (9552 == GlobalFiModInstNr[1]) || (9552 == GlobalFiModInstNr[2]) || (9552 == GlobalFiModInstNr[3]))));
	Tile mesh_5_22(
		.clock(clock),
		.io_in_a_0(r_182_0),
		.io_in_b_0(b_709_0),
		.io_in_d_0(b_1733_0),
		.io_in_control_0_dataflow(mesh_5_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2757_0),
		.io_in_last_0(r_3781_0),
		.io_in_valid_0(r_1733_0),
		.io_out_a_0(_mesh_5_22_io_out_a_0),
		.io_out_c_0(_mesh_5_22_io_out_c_0),
		.io_out_b_0(_mesh_5_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_22_io_out_id_0),
		.io_out_last_0(_mesh_5_22_io_out_last_0),
		.io_out_valid_0(_mesh_5_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9553 == GlobalFiModInstNr[0]) || (9553 == GlobalFiModInstNr[1]) || (9553 == GlobalFiModInstNr[2]) || (9553 == GlobalFiModInstNr[3]))));
	Tile mesh_5_23(
		.clock(clock),
		.io_in_a_0(r_183_0),
		.io_in_b_0(b_741_0),
		.io_in_d_0(b_1765_0),
		.io_in_control_0_dataflow(mesh_5_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2789_0),
		.io_in_last_0(r_3813_0),
		.io_in_valid_0(r_1765_0),
		.io_out_a_0(_mesh_5_23_io_out_a_0),
		.io_out_c_0(_mesh_5_23_io_out_c_0),
		.io_out_b_0(_mesh_5_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_23_io_out_id_0),
		.io_out_last_0(_mesh_5_23_io_out_last_0),
		.io_out_valid_0(_mesh_5_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9554 == GlobalFiModInstNr[0]) || (9554 == GlobalFiModInstNr[1]) || (9554 == GlobalFiModInstNr[2]) || (9554 == GlobalFiModInstNr[3]))));
	Tile mesh_5_24(
		.clock(clock),
		.io_in_a_0(r_184_0),
		.io_in_b_0(b_773_0),
		.io_in_d_0(b_1797_0),
		.io_in_control_0_dataflow(mesh_5_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2821_0),
		.io_in_last_0(r_3845_0),
		.io_in_valid_0(r_1797_0),
		.io_out_a_0(_mesh_5_24_io_out_a_0),
		.io_out_c_0(_mesh_5_24_io_out_c_0),
		.io_out_b_0(_mesh_5_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_24_io_out_id_0),
		.io_out_last_0(_mesh_5_24_io_out_last_0),
		.io_out_valid_0(_mesh_5_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9555 == GlobalFiModInstNr[0]) || (9555 == GlobalFiModInstNr[1]) || (9555 == GlobalFiModInstNr[2]) || (9555 == GlobalFiModInstNr[3]))));
	Tile mesh_5_25(
		.clock(clock),
		.io_in_a_0(r_185_0),
		.io_in_b_0(b_805_0),
		.io_in_d_0(b_1829_0),
		.io_in_control_0_dataflow(mesh_5_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2853_0),
		.io_in_last_0(r_3877_0),
		.io_in_valid_0(r_1829_0),
		.io_out_a_0(_mesh_5_25_io_out_a_0),
		.io_out_c_0(_mesh_5_25_io_out_c_0),
		.io_out_b_0(_mesh_5_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_25_io_out_id_0),
		.io_out_last_0(_mesh_5_25_io_out_last_0),
		.io_out_valid_0(_mesh_5_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9556 == GlobalFiModInstNr[0]) || (9556 == GlobalFiModInstNr[1]) || (9556 == GlobalFiModInstNr[2]) || (9556 == GlobalFiModInstNr[3]))));
	Tile mesh_5_26(
		.clock(clock),
		.io_in_a_0(r_186_0),
		.io_in_b_0(b_837_0),
		.io_in_d_0(b_1861_0),
		.io_in_control_0_dataflow(mesh_5_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2885_0),
		.io_in_last_0(r_3909_0),
		.io_in_valid_0(r_1861_0),
		.io_out_a_0(_mesh_5_26_io_out_a_0),
		.io_out_c_0(_mesh_5_26_io_out_c_0),
		.io_out_b_0(_mesh_5_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_26_io_out_id_0),
		.io_out_last_0(_mesh_5_26_io_out_last_0),
		.io_out_valid_0(_mesh_5_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9557 == GlobalFiModInstNr[0]) || (9557 == GlobalFiModInstNr[1]) || (9557 == GlobalFiModInstNr[2]) || (9557 == GlobalFiModInstNr[3]))));
	Tile mesh_5_27(
		.clock(clock),
		.io_in_a_0(r_187_0),
		.io_in_b_0(b_869_0),
		.io_in_d_0(b_1893_0),
		.io_in_control_0_dataflow(mesh_5_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2917_0),
		.io_in_last_0(r_3941_0),
		.io_in_valid_0(r_1893_0),
		.io_out_a_0(_mesh_5_27_io_out_a_0),
		.io_out_c_0(_mesh_5_27_io_out_c_0),
		.io_out_b_0(_mesh_5_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_27_io_out_id_0),
		.io_out_last_0(_mesh_5_27_io_out_last_0),
		.io_out_valid_0(_mesh_5_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9558 == GlobalFiModInstNr[0]) || (9558 == GlobalFiModInstNr[1]) || (9558 == GlobalFiModInstNr[2]) || (9558 == GlobalFiModInstNr[3]))));
	Tile mesh_5_28(
		.clock(clock),
		.io_in_a_0(r_188_0),
		.io_in_b_0(b_901_0),
		.io_in_d_0(b_1925_0),
		.io_in_control_0_dataflow(mesh_5_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2949_0),
		.io_in_last_0(r_3973_0),
		.io_in_valid_0(r_1925_0),
		.io_out_a_0(_mesh_5_28_io_out_a_0),
		.io_out_c_0(_mesh_5_28_io_out_c_0),
		.io_out_b_0(_mesh_5_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_28_io_out_id_0),
		.io_out_last_0(_mesh_5_28_io_out_last_0),
		.io_out_valid_0(_mesh_5_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9559 == GlobalFiModInstNr[0]) || (9559 == GlobalFiModInstNr[1]) || (9559 == GlobalFiModInstNr[2]) || (9559 == GlobalFiModInstNr[3]))));
	Tile mesh_5_29(
		.clock(clock),
		.io_in_a_0(r_189_0),
		.io_in_b_0(b_933_0),
		.io_in_d_0(b_1957_0),
		.io_in_control_0_dataflow(mesh_5_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2981_0),
		.io_in_last_0(r_4005_0),
		.io_in_valid_0(r_1957_0),
		.io_out_a_0(_mesh_5_29_io_out_a_0),
		.io_out_c_0(_mesh_5_29_io_out_c_0),
		.io_out_b_0(_mesh_5_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_29_io_out_id_0),
		.io_out_last_0(_mesh_5_29_io_out_last_0),
		.io_out_valid_0(_mesh_5_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9560 == GlobalFiModInstNr[0]) || (9560 == GlobalFiModInstNr[1]) || (9560 == GlobalFiModInstNr[2]) || (9560 == GlobalFiModInstNr[3]))));
	Tile mesh_5_30(
		.clock(clock),
		.io_in_a_0(r_190_0),
		.io_in_b_0(b_965_0),
		.io_in_d_0(b_1989_0),
		.io_in_control_0_dataflow(mesh_5_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3013_0),
		.io_in_last_0(r_4037_0),
		.io_in_valid_0(r_1989_0),
		.io_out_a_0(_mesh_5_30_io_out_a_0),
		.io_out_c_0(_mesh_5_30_io_out_c_0),
		.io_out_b_0(_mesh_5_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_30_io_out_id_0),
		.io_out_last_0(_mesh_5_30_io_out_last_0),
		.io_out_valid_0(_mesh_5_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9561 == GlobalFiModInstNr[0]) || (9561 == GlobalFiModInstNr[1]) || (9561 == GlobalFiModInstNr[2]) || (9561 == GlobalFiModInstNr[3]))));
	Tile mesh_5_31(
		.clock(clock),
		.io_in_a_0(r_191_0),
		.io_in_b_0(b_997_0),
		.io_in_d_0(b_2021_0),
		.io_in_control_0_dataflow(mesh_5_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3045_0),
		.io_in_last_0(r_4069_0),
		.io_in_valid_0(r_2021_0),
		.io_out_a_0(_mesh_5_31_io_out_a_0),
		.io_out_c_0(_mesh_5_31_io_out_c_0),
		.io_out_b_0(_mesh_5_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_31_io_out_id_0),
		.io_out_last_0(_mesh_5_31_io_out_last_0),
		.io_out_valid_0(_mesh_5_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9562 == GlobalFiModInstNr[0]) || (9562 == GlobalFiModInstNr[1]) || (9562 == GlobalFiModInstNr[2]) || (9562 == GlobalFiModInstNr[3]))));
	Tile mesh_6_0(
		.clock(clock),
		.io_in_a_0(r_192_0),
		.io_in_b_0(b_6_0),
		.io_in_d_0(b_1030_0),
		.io_in_control_0_dataflow(mesh_6_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2054_0),
		.io_in_last_0(r_3078_0),
		.io_in_valid_0(r_1030_0),
		.io_out_a_0(_mesh_6_0_io_out_a_0),
		.io_out_c_0(_mesh_6_0_io_out_c_0),
		.io_out_b_0(_mesh_6_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_0_io_out_id_0),
		.io_out_last_0(_mesh_6_0_io_out_last_0),
		.io_out_valid_0(_mesh_6_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9563 == GlobalFiModInstNr[0]) || (9563 == GlobalFiModInstNr[1]) || (9563 == GlobalFiModInstNr[2]) || (9563 == GlobalFiModInstNr[3]))));
	Tile mesh_6_1(
		.clock(clock),
		.io_in_a_0(r_193_0),
		.io_in_b_0(b_38_0),
		.io_in_d_0(b_1062_0),
		.io_in_control_0_dataflow(mesh_6_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2086_0),
		.io_in_last_0(r_3110_0),
		.io_in_valid_0(r_1062_0),
		.io_out_a_0(_mesh_6_1_io_out_a_0),
		.io_out_c_0(_mesh_6_1_io_out_c_0),
		.io_out_b_0(_mesh_6_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_1_io_out_id_0),
		.io_out_last_0(_mesh_6_1_io_out_last_0),
		.io_out_valid_0(_mesh_6_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9564 == GlobalFiModInstNr[0]) || (9564 == GlobalFiModInstNr[1]) || (9564 == GlobalFiModInstNr[2]) || (9564 == GlobalFiModInstNr[3]))));
	Tile mesh_6_2(
		.clock(clock),
		.io_in_a_0(r_194_0),
		.io_in_b_0(b_70_0),
		.io_in_d_0(b_1094_0),
		.io_in_control_0_dataflow(mesh_6_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2118_0),
		.io_in_last_0(r_3142_0),
		.io_in_valid_0(r_1094_0),
		.io_out_a_0(_mesh_6_2_io_out_a_0),
		.io_out_c_0(_mesh_6_2_io_out_c_0),
		.io_out_b_0(_mesh_6_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_2_io_out_id_0),
		.io_out_last_0(_mesh_6_2_io_out_last_0),
		.io_out_valid_0(_mesh_6_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9565 == GlobalFiModInstNr[0]) || (9565 == GlobalFiModInstNr[1]) || (9565 == GlobalFiModInstNr[2]) || (9565 == GlobalFiModInstNr[3]))));
	Tile mesh_6_3(
		.clock(clock),
		.io_in_a_0(r_195_0),
		.io_in_b_0(b_102_0),
		.io_in_d_0(b_1126_0),
		.io_in_control_0_dataflow(mesh_6_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2150_0),
		.io_in_last_0(r_3174_0),
		.io_in_valid_0(r_1126_0),
		.io_out_a_0(_mesh_6_3_io_out_a_0),
		.io_out_c_0(_mesh_6_3_io_out_c_0),
		.io_out_b_0(_mesh_6_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_3_io_out_id_0),
		.io_out_last_0(_mesh_6_3_io_out_last_0),
		.io_out_valid_0(_mesh_6_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9566 == GlobalFiModInstNr[0]) || (9566 == GlobalFiModInstNr[1]) || (9566 == GlobalFiModInstNr[2]) || (9566 == GlobalFiModInstNr[3]))));
	Tile mesh_6_4(
		.clock(clock),
		.io_in_a_0(r_196_0),
		.io_in_b_0(b_134_0),
		.io_in_d_0(b_1158_0),
		.io_in_control_0_dataflow(mesh_6_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2182_0),
		.io_in_last_0(r_3206_0),
		.io_in_valid_0(r_1158_0),
		.io_out_a_0(_mesh_6_4_io_out_a_0),
		.io_out_c_0(_mesh_6_4_io_out_c_0),
		.io_out_b_0(_mesh_6_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_4_io_out_id_0),
		.io_out_last_0(_mesh_6_4_io_out_last_0),
		.io_out_valid_0(_mesh_6_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9567 == GlobalFiModInstNr[0]) || (9567 == GlobalFiModInstNr[1]) || (9567 == GlobalFiModInstNr[2]) || (9567 == GlobalFiModInstNr[3]))));
	Tile mesh_6_5(
		.clock(clock),
		.io_in_a_0(r_197_0),
		.io_in_b_0(b_166_0),
		.io_in_d_0(b_1190_0),
		.io_in_control_0_dataflow(mesh_6_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2214_0),
		.io_in_last_0(r_3238_0),
		.io_in_valid_0(r_1190_0),
		.io_out_a_0(_mesh_6_5_io_out_a_0),
		.io_out_c_0(_mesh_6_5_io_out_c_0),
		.io_out_b_0(_mesh_6_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_5_io_out_id_0),
		.io_out_last_0(_mesh_6_5_io_out_last_0),
		.io_out_valid_0(_mesh_6_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9568 == GlobalFiModInstNr[0]) || (9568 == GlobalFiModInstNr[1]) || (9568 == GlobalFiModInstNr[2]) || (9568 == GlobalFiModInstNr[3]))));
	Tile mesh_6_6(
		.clock(clock),
		.io_in_a_0(r_198_0),
		.io_in_b_0(b_198_0),
		.io_in_d_0(b_1222_0),
		.io_in_control_0_dataflow(mesh_6_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2246_0),
		.io_in_last_0(r_3270_0),
		.io_in_valid_0(r_1222_0),
		.io_out_a_0(_mesh_6_6_io_out_a_0),
		.io_out_c_0(_mesh_6_6_io_out_c_0),
		.io_out_b_0(_mesh_6_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_6_io_out_id_0),
		.io_out_last_0(_mesh_6_6_io_out_last_0),
		.io_out_valid_0(_mesh_6_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9569 == GlobalFiModInstNr[0]) || (9569 == GlobalFiModInstNr[1]) || (9569 == GlobalFiModInstNr[2]) || (9569 == GlobalFiModInstNr[3]))));
	Tile mesh_6_7(
		.clock(clock),
		.io_in_a_0(r_199_0),
		.io_in_b_0(b_230_0),
		.io_in_d_0(b_1254_0),
		.io_in_control_0_dataflow(mesh_6_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2278_0),
		.io_in_last_0(r_3302_0),
		.io_in_valid_0(r_1254_0),
		.io_out_a_0(_mesh_6_7_io_out_a_0),
		.io_out_c_0(_mesh_6_7_io_out_c_0),
		.io_out_b_0(_mesh_6_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_7_io_out_id_0),
		.io_out_last_0(_mesh_6_7_io_out_last_0),
		.io_out_valid_0(_mesh_6_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9570 == GlobalFiModInstNr[0]) || (9570 == GlobalFiModInstNr[1]) || (9570 == GlobalFiModInstNr[2]) || (9570 == GlobalFiModInstNr[3]))));
	Tile mesh_6_8(
		.clock(clock),
		.io_in_a_0(r_200_0),
		.io_in_b_0(b_262_0),
		.io_in_d_0(b_1286_0),
		.io_in_control_0_dataflow(mesh_6_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2310_0),
		.io_in_last_0(r_3334_0),
		.io_in_valid_0(r_1286_0),
		.io_out_a_0(_mesh_6_8_io_out_a_0),
		.io_out_c_0(_mesh_6_8_io_out_c_0),
		.io_out_b_0(_mesh_6_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_8_io_out_id_0),
		.io_out_last_0(_mesh_6_8_io_out_last_0),
		.io_out_valid_0(_mesh_6_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9571 == GlobalFiModInstNr[0]) || (9571 == GlobalFiModInstNr[1]) || (9571 == GlobalFiModInstNr[2]) || (9571 == GlobalFiModInstNr[3]))));
	Tile mesh_6_9(
		.clock(clock),
		.io_in_a_0(r_201_0),
		.io_in_b_0(b_294_0),
		.io_in_d_0(b_1318_0),
		.io_in_control_0_dataflow(mesh_6_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2342_0),
		.io_in_last_0(r_3366_0),
		.io_in_valid_0(r_1318_0),
		.io_out_a_0(_mesh_6_9_io_out_a_0),
		.io_out_c_0(_mesh_6_9_io_out_c_0),
		.io_out_b_0(_mesh_6_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_9_io_out_id_0),
		.io_out_last_0(_mesh_6_9_io_out_last_0),
		.io_out_valid_0(_mesh_6_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9572 == GlobalFiModInstNr[0]) || (9572 == GlobalFiModInstNr[1]) || (9572 == GlobalFiModInstNr[2]) || (9572 == GlobalFiModInstNr[3]))));
	Tile mesh_6_10(
		.clock(clock),
		.io_in_a_0(r_202_0),
		.io_in_b_0(b_326_0),
		.io_in_d_0(b_1350_0),
		.io_in_control_0_dataflow(mesh_6_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2374_0),
		.io_in_last_0(r_3398_0),
		.io_in_valid_0(r_1350_0),
		.io_out_a_0(_mesh_6_10_io_out_a_0),
		.io_out_c_0(_mesh_6_10_io_out_c_0),
		.io_out_b_0(_mesh_6_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_10_io_out_id_0),
		.io_out_last_0(_mesh_6_10_io_out_last_0),
		.io_out_valid_0(_mesh_6_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9573 == GlobalFiModInstNr[0]) || (9573 == GlobalFiModInstNr[1]) || (9573 == GlobalFiModInstNr[2]) || (9573 == GlobalFiModInstNr[3]))));
	Tile mesh_6_11(
		.clock(clock),
		.io_in_a_0(r_203_0),
		.io_in_b_0(b_358_0),
		.io_in_d_0(b_1382_0),
		.io_in_control_0_dataflow(mesh_6_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2406_0),
		.io_in_last_0(r_3430_0),
		.io_in_valid_0(r_1382_0),
		.io_out_a_0(_mesh_6_11_io_out_a_0),
		.io_out_c_0(_mesh_6_11_io_out_c_0),
		.io_out_b_0(_mesh_6_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_11_io_out_id_0),
		.io_out_last_0(_mesh_6_11_io_out_last_0),
		.io_out_valid_0(_mesh_6_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9574 == GlobalFiModInstNr[0]) || (9574 == GlobalFiModInstNr[1]) || (9574 == GlobalFiModInstNr[2]) || (9574 == GlobalFiModInstNr[3]))));
	Tile mesh_6_12(
		.clock(clock),
		.io_in_a_0(r_204_0),
		.io_in_b_0(b_390_0),
		.io_in_d_0(b_1414_0),
		.io_in_control_0_dataflow(mesh_6_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2438_0),
		.io_in_last_0(r_3462_0),
		.io_in_valid_0(r_1414_0),
		.io_out_a_0(_mesh_6_12_io_out_a_0),
		.io_out_c_0(_mesh_6_12_io_out_c_0),
		.io_out_b_0(_mesh_6_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_12_io_out_id_0),
		.io_out_last_0(_mesh_6_12_io_out_last_0),
		.io_out_valid_0(_mesh_6_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9575 == GlobalFiModInstNr[0]) || (9575 == GlobalFiModInstNr[1]) || (9575 == GlobalFiModInstNr[2]) || (9575 == GlobalFiModInstNr[3]))));
	Tile mesh_6_13(
		.clock(clock),
		.io_in_a_0(r_205_0),
		.io_in_b_0(b_422_0),
		.io_in_d_0(b_1446_0),
		.io_in_control_0_dataflow(mesh_6_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2470_0),
		.io_in_last_0(r_3494_0),
		.io_in_valid_0(r_1446_0),
		.io_out_a_0(_mesh_6_13_io_out_a_0),
		.io_out_c_0(_mesh_6_13_io_out_c_0),
		.io_out_b_0(_mesh_6_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_13_io_out_id_0),
		.io_out_last_0(_mesh_6_13_io_out_last_0),
		.io_out_valid_0(_mesh_6_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9576 == GlobalFiModInstNr[0]) || (9576 == GlobalFiModInstNr[1]) || (9576 == GlobalFiModInstNr[2]) || (9576 == GlobalFiModInstNr[3]))));
	Tile mesh_6_14(
		.clock(clock),
		.io_in_a_0(r_206_0),
		.io_in_b_0(b_454_0),
		.io_in_d_0(b_1478_0),
		.io_in_control_0_dataflow(mesh_6_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2502_0),
		.io_in_last_0(r_3526_0),
		.io_in_valid_0(r_1478_0),
		.io_out_a_0(_mesh_6_14_io_out_a_0),
		.io_out_c_0(_mesh_6_14_io_out_c_0),
		.io_out_b_0(_mesh_6_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_14_io_out_id_0),
		.io_out_last_0(_mesh_6_14_io_out_last_0),
		.io_out_valid_0(_mesh_6_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9577 == GlobalFiModInstNr[0]) || (9577 == GlobalFiModInstNr[1]) || (9577 == GlobalFiModInstNr[2]) || (9577 == GlobalFiModInstNr[3]))));
	Tile mesh_6_15(
		.clock(clock),
		.io_in_a_0(r_207_0),
		.io_in_b_0(b_486_0),
		.io_in_d_0(b_1510_0),
		.io_in_control_0_dataflow(mesh_6_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2534_0),
		.io_in_last_0(r_3558_0),
		.io_in_valid_0(r_1510_0),
		.io_out_a_0(_mesh_6_15_io_out_a_0),
		.io_out_c_0(_mesh_6_15_io_out_c_0),
		.io_out_b_0(_mesh_6_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_15_io_out_id_0),
		.io_out_last_0(_mesh_6_15_io_out_last_0),
		.io_out_valid_0(_mesh_6_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9578 == GlobalFiModInstNr[0]) || (9578 == GlobalFiModInstNr[1]) || (9578 == GlobalFiModInstNr[2]) || (9578 == GlobalFiModInstNr[3]))));
	Tile mesh_6_16(
		.clock(clock),
		.io_in_a_0(r_208_0),
		.io_in_b_0(b_518_0),
		.io_in_d_0(b_1542_0),
		.io_in_control_0_dataflow(mesh_6_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2566_0),
		.io_in_last_0(r_3590_0),
		.io_in_valid_0(r_1542_0),
		.io_out_a_0(_mesh_6_16_io_out_a_0),
		.io_out_c_0(_mesh_6_16_io_out_c_0),
		.io_out_b_0(_mesh_6_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_16_io_out_id_0),
		.io_out_last_0(_mesh_6_16_io_out_last_0),
		.io_out_valid_0(_mesh_6_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9579 == GlobalFiModInstNr[0]) || (9579 == GlobalFiModInstNr[1]) || (9579 == GlobalFiModInstNr[2]) || (9579 == GlobalFiModInstNr[3]))));
	Tile mesh_6_17(
		.clock(clock),
		.io_in_a_0(r_209_0),
		.io_in_b_0(b_550_0),
		.io_in_d_0(b_1574_0),
		.io_in_control_0_dataflow(mesh_6_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2598_0),
		.io_in_last_0(r_3622_0),
		.io_in_valid_0(r_1574_0),
		.io_out_a_0(_mesh_6_17_io_out_a_0),
		.io_out_c_0(_mesh_6_17_io_out_c_0),
		.io_out_b_0(_mesh_6_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_17_io_out_id_0),
		.io_out_last_0(_mesh_6_17_io_out_last_0),
		.io_out_valid_0(_mesh_6_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9580 == GlobalFiModInstNr[0]) || (9580 == GlobalFiModInstNr[1]) || (9580 == GlobalFiModInstNr[2]) || (9580 == GlobalFiModInstNr[3]))));
	Tile mesh_6_18(
		.clock(clock),
		.io_in_a_0(r_210_0),
		.io_in_b_0(b_582_0),
		.io_in_d_0(b_1606_0),
		.io_in_control_0_dataflow(mesh_6_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2630_0),
		.io_in_last_0(r_3654_0),
		.io_in_valid_0(r_1606_0),
		.io_out_a_0(_mesh_6_18_io_out_a_0),
		.io_out_c_0(_mesh_6_18_io_out_c_0),
		.io_out_b_0(_mesh_6_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_18_io_out_id_0),
		.io_out_last_0(_mesh_6_18_io_out_last_0),
		.io_out_valid_0(_mesh_6_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9581 == GlobalFiModInstNr[0]) || (9581 == GlobalFiModInstNr[1]) || (9581 == GlobalFiModInstNr[2]) || (9581 == GlobalFiModInstNr[3]))));
	Tile mesh_6_19(
		.clock(clock),
		.io_in_a_0(r_211_0),
		.io_in_b_0(b_614_0),
		.io_in_d_0(b_1638_0),
		.io_in_control_0_dataflow(mesh_6_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2662_0),
		.io_in_last_0(r_3686_0),
		.io_in_valid_0(r_1638_0),
		.io_out_a_0(_mesh_6_19_io_out_a_0),
		.io_out_c_0(_mesh_6_19_io_out_c_0),
		.io_out_b_0(_mesh_6_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_19_io_out_id_0),
		.io_out_last_0(_mesh_6_19_io_out_last_0),
		.io_out_valid_0(_mesh_6_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9582 == GlobalFiModInstNr[0]) || (9582 == GlobalFiModInstNr[1]) || (9582 == GlobalFiModInstNr[2]) || (9582 == GlobalFiModInstNr[3]))));
	Tile mesh_6_20(
		.clock(clock),
		.io_in_a_0(r_212_0),
		.io_in_b_0(b_646_0),
		.io_in_d_0(b_1670_0),
		.io_in_control_0_dataflow(mesh_6_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2694_0),
		.io_in_last_0(r_3718_0),
		.io_in_valid_0(r_1670_0),
		.io_out_a_0(_mesh_6_20_io_out_a_0),
		.io_out_c_0(_mesh_6_20_io_out_c_0),
		.io_out_b_0(_mesh_6_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_20_io_out_id_0),
		.io_out_last_0(_mesh_6_20_io_out_last_0),
		.io_out_valid_0(_mesh_6_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9583 == GlobalFiModInstNr[0]) || (9583 == GlobalFiModInstNr[1]) || (9583 == GlobalFiModInstNr[2]) || (9583 == GlobalFiModInstNr[3]))));
	Tile mesh_6_21(
		.clock(clock),
		.io_in_a_0(r_213_0),
		.io_in_b_0(b_678_0),
		.io_in_d_0(b_1702_0),
		.io_in_control_0_dataflow(mesh_6_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2726_0),
		.io_in_last_0(r_3750_0),
		.io_in_valid_0(r_1702_0),
		.io_out_a_0(_mesh_6_21_io_out_a_0),
		.io_out_c_0(_mesh_6_21_io_out_c_0),
		.io_out_b_0(_mesh_6_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_21_io_out_id_0),
		.io_out_last_0(_mesh_6_21_io_out_last_0),
		.io_out_valid_0(_mesh_6_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9584 == GlobalFiModInstNr[0]) || (9584 == GlobalFiModInstNr[1]) || (9584 == GlobalFiModInstNr[2]) || (9584 == GlobalFiModInstNr[3]))));
	Tile mesh_6_22(
		.clock(clock),
		.io_in_a_0(r_214_0),
		.io_in_b_0(b_710_0),
		.io_in_d_0(b_1734_0),
		.io_in_control_0_dataflow(mesh_6_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2758_0),
		.io_in_last_0(r_3782_0),
		.io_in_valid_0(r_1734_0),
		.io_out_a_0(_mesh_6_22_io_out_a_0),
		.io_out_c_0(_mesh_6_22_io_out_c_0),
		.io_out_b_0(_mesh_6_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_22_io_out_id_0),
		.io_out_last_0(_mesh_6_22_io_out_last_0),
		.io_out_valid_0(_mesh_6_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9585 == GlobalFiModInstNr[0]) || (9585 == GlobalFiModInstNr[1]) || (9585 == GlobalFiModInstNr[2]) || (9585 == GlobalFiModInstNr[3]))));
	Tile mesh_6_23(
		.clock(clock),
		.io_in_a_0(r_215_0),
		.io_in_b_0(b_742_0),
		.io_in_d_0(b_1766_0),
		.io_in_control_0_dataflow(mesh_6_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2790_0),
		.io_in_last_0(r_3814_0),
		.io_in_valid_0(r_1766_0),
		.io_out_a_0(_mesh_6_23_io_out_a_0),
		.io_out_c_0(_mesh_6_23_io_out_c_0),
		.io_out_b_0(_mesh_6_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_23_io_out_id_0),
		.io_out_last_0(_mesh_6_23_io_out_last_0),
		.io_out_valid_0(_mesh_6_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9586 == GlobalFiModInstNr[0]) || (9586 == GlobalFiModInstNr[1]) || (9586 == GlobalFiModInstNr[2]) || (9586 == GlobalFiModInstNr[3]))));
	Tile mesh_6_24(
		.clock(clock),
		.io_in_a_0(r_216_0),
		.io_in_b_0(b_774_0),
		.io_in_d_0(b_1798_0),
		.io_in_control_0_dataflow(mesh_6_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2822_0),
		.io_in_last_0(r_3846_0),
		.io_in_valid_0(r_1798_0),
		.io_out_a_0(_mesh_6_24_io_out_a_0),
		.io_out_c_0(_mesh_6_24_io_out_c_0),
		.io_out_b_0(_mesh_6_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_24_io_out_id_0),
		.io_out_last_0(_mesh_6_24_io_out_last_0),
		.io_out_valid_0(_mesh_6_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9587 == GlobalFiModInstNr[0]) || (9587 == GlobalFiModInstNr[1]) || (9587 == GlobalFiModInstNr[2]) || (9587 == GlobalFiModInstNr[3]))));
	Tile mesh_6_25(
		.clock(clock),
		.io_in_a_0(r_217_0),
		.io_in_b_0(b_806_0),
		.io_in_d_0(b_1830_0),
		.io_in_control_0_dataflow(mesh_6_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2854_0),
		.io_in_last_0(r_3878_0),
		.io_in_valid_0(r_1830_0),
		.io_out_a_0(_mesh_6_25_io_out_a_0),
		.io_out_c_0(_mesh_6_25_io_out_c_0),
		.io_out_b_0(_mesh_6_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_25_io_out_id_0),
		.io_out_last_0(_mesh_6_25_io_out_last_0),
		.io_out_valid_0(_mesh_6_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9588 == GlobalFiModInstNr[0]) || (9588 == GlobalFiModInstNr[1]) || (9588 == GlobalFiModInstNr[2]) || (9588 == GlobalFiModInstNr[3]))));
	Tile mesh_6_26(
		.clock(clock),
		.io_in_a_0(r_218_0),
		.io_in_b_0(b_838_0),
		.io_in_d_0(b_1862_0),
		.io_in_control_0_dataflow(mesh_6_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2886_0),
		.io_in_last_0(r_3910_0),
		.io_in_valid_0(r_1862_0),
		.io_out_a_0(_mesh_6_26_io_out_a_0),
		.io_out_c_0(_mesh_6_26_io_out_c_0),
		.io_out_b_0(_mesh_6_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_26_io_out_id_0),
		.io_out_last_0(_mesh_6_26_io_out_last_0),
		.io_out_valid_0(_mesh_6_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9589 == GlobalFiModInstNr[0]) || (9589 == GlobalFiModInstNr[1]) || (9589 == GlobalFiModInstNr[2]) || (9589 == GlobalFiModInstNr[3]))));
	Tile mesh_6_27(
		.clock(clock),
		.io_in_a_0(r_219_0),
		.io_in_b_0(b_870_0),
		.io_in_d_0(b_1894_0),
		.io_in_control_0_dataflow(mesh_6_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2918_0),
		.io_in_last_0(r_3942_0),
		.io_in_valid_0(r_1894_0),
		.io_out_a_0(_mesh_6_27_io_out_a_0),
		.io_out_c_0(_mesh_6_27_io_out_c_0),
		.io_out_b_0(_mesh_6_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_27_io_out_id_0),
		.io_out_last_0(_mesh_6_27_io_out_last_0),
		.io_out_valid_0(_mesh_6_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9590 == GlobalFiModInstNr[0]) || (9590 == GlobalFiModInstNr[1]) || (9590 == GlobalFiModInstNr[2]) || (9590 == GlobalFiModInstNr[3]))));
	Tile mesh_6_28(
		.clock(clock),
		.io_in_a_0(r_220_0),
		.io_in_b_0(b_902_0),
		.io_in_d_0(b_1926_0),
		.io_in_control_0_dataflow(mesh_6_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2950_0),
		.io_in_last_0(r_3974_0),
		.io_in_valid_0(r_1926_0),
		.io_out_a_0(_mesh_6_28_io_out_a_0),
		.io_out_c_0(_mesh_6_28_io_out_c_0),
		.io_out_b_0(_mesh_6_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_28_io_out_id_0),
		.io_out_last_0(_mesh_6_28_io_out_last_0),
		.io_out_valid_0(_mesh_6_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9591 == GlobalFiModInstNr[0]) || (9591 == GlobalFiModInstNr[1]) || (9591 == GlobalFiModInstNr[2]) || (9591 == GlobalFiModInstNr[3]))));
	Tile mesh_6_29(
		.clock(clock),
		.io_in_a_0(r_221_0),
		.io_in_b_0(b_934_0),
		.io_in_d_0(b_1958_0),
		.io_in_control_0_dataflow(mesh_6_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2982_0),
		.io_in_last_0(r_4006_0),
		.io_in_valid_0(r_1958_0),
		.io_out_a_0(_mesh_6_29_io_out_a_0),
		.io_out_c_0(_mesh_6_29_io_out_c_0),
		.io_out_b_0(_mesh_6_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_29_io_out_id_0),
		.io_out_last_0(_mesh_6_29_io_out_last_0),
		.io_out_valid_0(_mesh_6_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9592 == GlobalFiModInstNr[0]) || (9592 == GlobalFiModInstNr[1]) || (9592 == GlobalFiModInstNr[2]) || (9592 == GlobalFiModInstNr[3]))));
	Tile mesh_6_30(
		.clock(clock),
		.io_in_a_0(r_222_0),
		.io_in_b_0(b_966_0),
		.io_in_d_0(b_1990_0),
		.io_in_control_0_dataflow(mesh_6_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3014_0),
		.io_in_last_0(r_4038_0),
		.io_in_valid_0(r_1990_0),
		.io_out_a_0(_mesh_6_30_io_out_a_0),
		.io_out_c_0(_mesh_6_30_io_out_c_0),
		.io_out_b_0(_mesh_6_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_30_io_out_id_0),
		.io_out_last_0(_mesh_6_30_io_out_last_0),
		.io_out_valid_0(_mesh_6_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9593 == GlobalFiModInstNr[0]) || (9593 == GlobalFiModInstNr[1]) || (9593 == GlobalFiModInstNr[2]) || (9593 == GlobalFiModInstNr[3]))));
	Tile mesh_6_31(
		.clock(clock),
		.io_in_a_0(r_223_0),
		.io_in_b_0(b_998_0),
		.io_in_d_0(b_2022_0),
		.io_in_control_0_dataflow(mesh_6_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3046_0),
		.io_in_last_0(r_4070_0),
		.io_in_valid_0(r_2022_0),
		.io_out_a_0(_mesh_6_31_io_out_a_0),
		.io_out_c_0(_mesh_6_31_io_out_c_0),
		.io_out_b_0(_mesh_6_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_31_io_out_id_0),
		.io_out_last_0(_mesh_6_31_io_out_last_0),
		.io_out_valid_0(_mesh_6_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9594 == GlobalFiModInstNr[0]) || (9594 == GlobalFiModInstNr[1]) || (9594 == GlobalFiModInstNr[2]) || (9594 == GlobalFiModInstNr[3]))));
	Tile mesh_7_0(
		.clock(clock),
		.io_in_a_0(r_224_0),
		.io_in_b_0(b_7_0),
		.io_in_d_0(b_1031_0),
		.io_in_control_0_dataflow(mesh_7_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2055_0),
		.io_in_last_0(r_3079_0),
		.io_in_valid_0(r_1031_0),
		.io_out_a_0(_mesh_7_0_io_out_a_0),
		.io_out_c_0(_mesh_7_0_io_out_c_0),
		.io_out_b_0(_mesh_7_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_0_io_out_id_0),
		.io_out_last_0(_mesh_7_0_io_out_last_0),
		.io_out_valid_0(_mesh_7_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9595 == GlobalFiModInstNr[0]) || (9595 == GlobalFiModInstNr[1]) || (9595 == GlobalFiModInstNr[2]) || (9595 == GlobalFiModInstNr[3]))));
	Tile mesh_7_1(
		.clock(clock),
		.io_in_a_0(r_225_0),
		.io_in_b_0(b_39_0),
		.io_in_d_0(b_1063_0),
		.io_in_control_0_dataflow(mesh_7_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2087_0),
		.io_in_last_0(r_3111_0),
		.io_in_valid_0(r_1063_0),
		.io_out_a_0(_mesh_7_1_io_out_a_0),
		.io_out_c_0(_mesh_7_1_io_out_c_0),
		.io_out_b_0(_mesh_7_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_1_io_out_id_0),
		.io_out_last_0(_mesh_7_1_io_out_last_0),
		.io_out_valid_0(_mesh_7_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9596 == GlobalFiModInstNr[0]) || (9596 == GlobalFiModInstNr[1]) || (9596 == GlobalFiModInstNr[2]) || (9596 == GlobalFiModInstNr[3]))));
	Tile mesh_7_2(
		.clock(clock),
		.io_in_a_0(r_226_0),
		.io_in_b_0(b_71_0),
		.io_in_d_0(b_1095_0),
		.io_in_control_0_dataflow(mesh_7_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2119_0),
		.io_in_last_0(r_3143_0),
		.io_in_valid_0(r_1095_0),
		.io_out_a_0(_mesh_7_2_io_out_a_0),
		.io_out_c_0(_mesh_7_2_io_out_c_0),
		.io_out_b_0(_mesh_7_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_2_io_out_id_0),
		.io_out_last_0(_mesh_7_2_io_out_last_0),
		.io_out_valid_0(_mesh_7_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9597 == GlobalFiModInstNr[0]) || (9597 == GlobalFiModInstNr[1]) || (9597 == GlobalFiModInstNr[2]) || (9597 == GlobalFiModInstNr[3]))));
	Tile mesh_7_3(
		.clock(clock),
		.io_in_a_0(r_227_0),
		.io_in_b_0(b_103_0),
		.io_in_d_0(b_1127_0),
		.io_in_control_0_dataflow(mesh_7_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2151_0),
		.io_in_last_0(r_3175_0),
		.io_in_valid_0(r_1127_0),
		.io_out_a_0(_mesh_7_3_io_out_a_0),
		.io_out_c_0(_mesh_7_3_io_out_c_0),
		.io_out_b_0(_mesh_7_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_3_io_out_id_0),
		.io_out_last_0(_mesh_7_3_io_out_last_0),
		.io_out_valid_0(_mesh_7_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9598 == GlobalFiModInstNr[0]) || (9598 == GlobalFiModInstNr[1]) || (9598 == GlobalFiModInstNr[2]) || (9598 == GlobalFiModInstNr[3]))));
	Tile mesh_7_4(
		.clock(clock),
		.io_in_a_0(r_228_0),
		.io_in_b_0(b_135_0),
		.io_in_d_0(b_1159_0),
		.io_in_control_0_dataflow(mesh_7_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2183_0),
		.io_in_last_0(r_3207_0),
		.io_in_valid_0(r_1159_0),
		.io_out_a_0(_mesh_7_4_io_out_a_0),
		.io_out_c_0(_mesh_7_4_io_out_c_0),
		.io_out_b_0(_mesh_7_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_4_io_out_id_0),
		.io_out_last_0(_mesh_7_4_io_out_last_0),
		.io_out_valid_0(_mesh_7_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9599 == GlobalFiModInstNr[0]) || (9599 == GlobalFiModInstNr[1]) || (9599 == GlobalFiModInstNr[2]) || (9599 == GlobalFiModInstNr[3]))));
	Tile mesh_7_5(
		.clock(clock),
		.io_in_a_0(r_229_0),
		.io_in_b_0(b_167_0),
		.io_in_d_0(b_1191_0),
		.io_in_control_0_dataflow(mesh_7_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2215_0),
		.io_in_last_0(r_3239_0),
		.io_in_valid_0(r_1191_0),
		.io_out_a_0(_mesh_7_5_io_out_a_0),
		.io_out_c_0(_mesh_7_5_io_out_c_0),
		.io_out_b_0(_mesh_7_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_5_io_out_id_0),
		.io_out_last_0(_mesh_7_5_io_out_last_0),
		.io_out_valid_0(_mesh_7_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9600 == GlobalFiModInstNr[0]) || (9600 == GlobalFiModInstNr[1]) || (9600 == GlobalFiModInstNr[2]) || (9600 == GlobalFiModInstNr[3]))));
	Tile mesh_7_6(
		.clock(clock),
		.io_in_a_0(r_230_0),
		.io_in_b_0(b_199_0),
		.io_in_d_0(b_1223_0),
		.io_in_control_0_dataflow(mesh_7_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2247_0),
		.io_in_last_0(r_3271_0),
		.io_in_valid_0(r_1223_0),
		.io_out_a_0(_mesh_7_6_io_out_a_0),
		.io_out_c_0(_mesh_7_6_io_out_c_0),
		.io_out_b_0(_mesh_7_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_6_io_out_id_0),
		.io_out_last_0(_mesh_7_6_io_out_last_0),
		.io_out_valid_0(_mesh_7_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9601 == GlobalFiModInstNr[0]) || (9601 == GlobalFiModInstNr[1]) || (9601 == GlobalFiModInstNr[2]) || (9601 == GlobalFiModInstNr[3]))));
	Tile mesh_7_7(
		.clock(clock),
		.io_in_a_0(r_231_0),
		.io_in_b_0(b_231_0),
		.io_in_d_0(b_1255_0),
		.io_in_control_0_dataflow(mesh_7_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2279_0),
		.io_in_last_0(r_3303_0),
		.io_in_valid_0(r_1255_0),
		.io_out_a_0(_mesh_7_7_io_out_a_0),
		.io_out_c_0(_mesh_7_7_io_out_c_0),
		.io_out_b_0(_mesh_7_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_7_io_out_id_0),
		.io_out_last_0(_mesh_7_7_io_out_last_0),
		.io_out_valid_0(_mesh_7_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9602 == GlobalFiModInstNr[0]) || (9602 == GlobalFiModInstNr[1]) || (9602 == GlobalFiModInstNr[2]) || (9602 == GlobalFiModInstNr[3]))));
	Tile mesh_7_8(
		.clock(clock),
		.io_in_a_0(r_232_0),
		.io_in_b_0(b_263_0),
		.io_in_d_0(b_1287_0),
		.io_in_control_0_dataflow(mesh_7_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2311_0),
		.io_in_last_0(r_3335_0),
		.io_in_valid_0(r_1287_0),
		.io_out_a_0(_mesh_7_8_io_out_a_0),
		.io_out_c_0(_mesh_7_8_io_out_c_0),
		.io_out_b_0(_mesh_7_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_8_io_out_id_0),
		.io_out_last_0(_mesh_7_8_io_out_last_0),
		.io_out_valid_0(_mesh_7_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9603 == GlobalFiModInstNr[0]) || (9603 == GlobalFiModInstNr[1]) || (9603 == GlobalFiModInstNr[2]) || (9603 == GlobalFiModInstNr[3]))));
	Tile mesh_7_9(
		.clock(clock),
		.io_in_a_0(r_233_0),
		.io_in_b_0(b_295_0),
		.io_in_d_0(b_1319_0),
		.io_in_control_0_dataflow(mesh_7_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2343_0),
		.io_in_last_0(r_3367_0),
		.io_in_valid_0(r_1319_0),
		.io_out_a_0(_mesh_7_9_io_out_a_0),
		.io_out_c_0(_mesh_7_9_io_out_c_0),
		.io_out_b_0(_mesh_7_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_9_io_out_id_0),
		.io_out_last_0(_mesh_7_9_io_out_last_0),
		.io_out_valid_0(_mesh_7_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9604 == GlobalFiModInstNr[0]) || (9604 == GlobalFiModInstNr[1]) || (9604 == GlobalFiModInstNr[2]) || (9604 == GlobalFiModInstNr[3]))));
	Tile mesh_7_10(
		.clock(clock),
		.io_in_a_0(r_234_0),
		.io_in_b_0(b_327_0),
		.io_in_d_0(b_1351_0),
		.io_in_control_0_dataflow(mesh_7_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2375_0),
		.io_in_last_0(r_3399_0),
		.io_in_valid_0(r_1351_0),
		.io_out_a_0(_mesh_7_10_io_out_a_0),
		.io_out_c_0(_mesh_7_10_io_out_c_0),
		.io_out_b_0(_mesh_7_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_10_io_out_id_0),
		.io_out_last_0(_mesh_7_10_io_out_last_0),
		.io_out_valid_0(_mesh_7_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9605 == GlobalFiModInstNr[0]) || (9605 == GlobalFiModInstNr[1]) || (9605 == GlobalFiModInstNr[2]) || (9605 == GlobalFiModInstNr[3]))));
	Tile mesh_7_11(
		.clock(clock),
		.io_in_a_0(r_235_0),
		.io_in_b_0(b_359_0),
		.io_in_d_0(b_1383_0),
		.io_in_control_0_dataflow(mesh_7_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2407_0),
		.io_in_last_0(r_3431_0),
		.io_in_valid_0(r_1383_0),
		.io_out_a_0(_mesh_7_11_io_out_a_0),
		.io_out_c_0(_mesh_7_11_io_out_c_0),
		.io_out_b_0(_mesh_7_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_11_io_out_id_0),
		.io_out_last_0(_mesh_7_11_io_out_last_0),
		.io_out_valid_0(_mesh_7_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9606 == GlobalFiModInstNr[0]) || (9606 == GlobalFiModInstNr[1]) || (9606 == GlobalFiModInstNr[2]) || (9606 == GlobalFiModInstNr[3]))));
	Tile mesh_7_12(
		.clock(clock),
		.io_in_a_0(r_236_0),
		.io_in_b_0(b_391_0),
		.io_in_d_0(b_1415_0),
		.io_in_control_0_dataflow(mesh_7_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2439_0),
		.io_in_last_0(r_3463_0),
		.io_in_valid_0(r_1415_0),
		.io_out_a_0(_mesh_7_12_io_out_a_0),
		.io_out_c_0(_mesh_7_12_io_out_c_0),
		.io_out_b_0(_mesh_7_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_12_io_out_id_0),
		.io_out_last_0(_mesh_7_12_io_out_last_0),
		.io_out_valid_0(_mesh_7_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9607 == GlobalFiModInstNr[0]) || (9607 == GlobalFiModInstNr[1]) || (9607 == GlobalFiModInstNr[2]) || (9607 == GlobalFiModInstNr[3]))));
	Tile mesh_7_13(
		.clock(clock),
		.io_in_a_0(r_237_0),
		.io_in_b_0(b_423_0),
		.io_in_d_0(b_1447_0),
		.io_in_control_0_dataflow(mesh_7_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2471_0),
		.io_in_last_0(r_3495_0),
		.io_in_valid_0(r_1447_0),
		.io_out_a_0(_mesh_7_13_io_out_a_0),
		.io_out_c_0(_mesh_7_13_io_out_c_0),
		.io_out_b_0(_mesh_7_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_13_io_out_id_0),
		.io_out_last_0(_mesh_7_13_io_out_last_0),
		.io_out_valid_0(_mesh_7_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9608 == GlobalFiModInstNr[0]) || (9608 == GlobalFiModInstNr[1]) || (9608 == GlobalFiModInstNr[2]) || (9608 == GlobalFiModInstNr[3]))));
	Tile mesh_7_14(
		.clock(clock),
		.io_in_a_0(r_238_0),
		.io_in_b_0(b_455_0),
		.io_in_d_0(b_1479_0),
		.io_in_control_0_dataflow(mesh_7_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2503_0),
		.io_in_last_0(r_3527_0),
		.io_in_valid_0(r_1479_0),
		.io_out_a_0(_mesh_7_14_io_out_a_0),
		.io_out_c_0(_mesh_7_14_io_out_c_0),
		.io_out_b_0(_mesh_7_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_14_io_out_id_0),
		.io_out_last_0(_mesh_7_14_io_out_last_0),
		.io_out_valid_0(_mesh_7_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9609 == GlobalFiModInstNr[0]) || (9609 == GlobalFiModInstNr[1]) || (9609 == GlobalFiModInstNr[2]) || (9609 == GlobalFiModInstNr[3]))));
	Tile mesh_7_15(
		.clock(clock),
		.io_in_a_0(r_239_0),
		.io_in_b_0(b_487_0),
		.io_in_d_0(b_1511_0),
		.io_in_control_0_dataflow(mesh_7_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2535_0),
		.io_in_last_0(r_3559_0),
		.io_in_valid_0(r_1511_0),
		.io_out_a_0(_mesh_7_15_io_out_a_0),
		.io_out_c_0(_mesh_7_15_io_out_c_0),
		.io_out_b_0(_mesh_7_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_15_io_out_id_0),
		.io_out_last_0(_mesh_7_15_io_out_last_0),
		.io_out_valid_0(_mesh_7_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9610 == GlobalFiModInstNr[0]) || (9610 == GlobalFiModInstNr[1]) || (9610 == GlobalFiModInstNr[2]) || (9610 == GlobalFiModInstNr[3]))));
	Tile mesh_7_16(
		.clock(clock),
		.io_in_a_0(r_240_0),
		.io_in_b_0(b_519_0),
		.io_in_d_0(b_1543_0),
		.io_in_control_0_dataflow(mesh_7_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2567_0),
		.io_in_last_0(r_3591_0),
		.io_in_valid_0(r_1543_0),
		.io_out_a_0(_mesh_7_16_io_out_a_0),
		.io_out_c_0(_mesh_7_16_io_out_c_0),
		.io_out_b_0(_mesh_7_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_16_io_out_id_0),
		.io_out_last_0(_mesh_7_16_io_out_last_0),
		.io_out_valid_0(_mesh_7_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9611 == GlobalFiModInstNr[0]) || (9611 == GlobalFiModInstNr[1]) || (9611 == GlobalFiModInstNr[2]) || (9611 == GlobalFiModInstNr[3]))));
	Tile mesh_7_17(
		.clock(clock),
		.io_in_a_0(r_241_0),
		.io_in_b_0(b_551_0),
		.io_in_d_0(b_1575_0),
		.io_in_control_0_dataflow(mesh_7_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2599_0),
		.io_in_last_0(r_3623_0),
		.io_in_valid_0(r_1575_0),
		.io_out_a_0(_mesh_7_17_io_out_a_0),
		.io_out_c_0(_mesh_7_17_io_out_c_0),
		.io_out_b_0(_mesh_7_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_17_io_out_id_0),
		.io_out_last_0(_mesh_7_17_io_out_last_0),
		.io_out_valid_0(_mesh_7_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9612 == GlobalFiModInstNr[0]) || (9612 == GlobalFiModInstNr[1]) || (9612 == GlobalFiModInstNr[2]) || (9612 == GlobalFiModInstNr[3]))));
	Tile mesh_7_18(
		.clock(clock),
		.io_in_a_0(r_242_0),
		.io_in_b_0(b_583_0),
		.io_in_d_0(b_1607_0),
		.io_in_control_0_dataflow(mesh_7_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2631_0),
		.io_in_last_0(r_3655_0),
		.io_in_valid_0(r_1607_0),
		.io_out_a_0(_mesh_7_18_io_out_a_0),
		.io_out_c_0(_mesh_7_18_io_out_c_0),
		.io_out_b_0(_mesh_7_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_18_io_out_id_0),
		.io_out_last_0(_mesh_7_18_io_out_last_0),
		.io_out_valid_0(_mesh_7_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9613 == GlobalFiModInstNr[0]) || (9613 == GlobalFiModInstNr[1]) || (9613 == GlobalFiModInstNr[2]) || (9613 == GlobalFiModInstNr[3]))));
	Tile mesh_7_19(
		.clock(clock),
		.io_in_a_0(r_243_0),
		.io_in_b_0(b_615_0),
		.io_in_d_0(b_1639_0),
		.io_in_control_0_dataflow(mesh_7_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2663_0),
		.io_in_last_0(r_3687_0),
		.io_in_valid_0(r_1639_0),
		.io_out_a_0(_mesh_7_19_io_out_a_0),
		.io_out_c_0(_mesh_7_19_io_out_c_0),
		.io_out_b_0(_mesh_7_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_19_io_out_id_0),
		.io_out_last_0(_mesh_7_19_io_out_last_0),
		.io_out_valid_0(_mesh_7_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9614 == GlobalFiModInstNr[0]) || (9614 == GlobalFiModInstNr[1]) || (9614 == GlobalFiModInstNr[2]) || (9614 == GlobalFiModInstNr[3]))));
	Tile mesh_7_20(
		.clock(clock),
		.io_in_a_0(r_244_0),
		.io_in_b_0(b_647_0),
		.io_in_d_0(b_1671_0),
		.io_in_control_0_dataflow(mesh_7_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2695_0),
		.io_in_last_0(r_3719_0),
		.io_in_valid_0(r_1671_0),
		.io_out_a_0(_mesh_7_20_io_out_a_0),
		.io_out_c_0(_mesh_7_20_io_out_c_0),
		.io_out_b_0(_mesh_7_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_20_io_out_id_0),
		.io_out_last_0(_mesh_7_20_io_out_last_0),
		.io_out_valid_0(_mesh_7_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9615 == GlobalFiModInstNr[0]) || (9615 == GlobalFiModInstNr[1]) || (9615 == GlobalFiModInstNr[2]) || (9615 == GlobalFiModInstNr[3]))));
	Tile mesh_7_21(
		.clock(clock),
		.io_in_a_0(r_245_0),
		.io_in_b_0(b_679_0),
		.io_in_d_0(b_1703_0),
		.io_in_control_0_dataflow(mesh_7_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2727_0),
		.io_in_last_0(r_3751_0),
		.io_in_valid_0(r_1703_0),
		.io_out_a_0(_mesh_7_21_io_out_a_0),
		.io_out_c_0(_mesh_7_21_io_out_c_0),
		.io_out_b_0(_mesh_7_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_21_io_out_id_0),
		.io_out_last_0(_mesh_7_21_io_out_last_0),
		.io_out_valid_0(_mesh_7_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9616 == GlobalFiModInstNr[0]) || (9616 == GlobalFiModInstNr[1]) || (9616 == GlobalFiModInstNr[2]) || (9616 == GlobalFiModInstNr[3]))));
	Tile mesh_7_22(
		.clock(clock),
		.io_in_a_0(r_246_0),
		.io_in_b_0(b_711_0),
		.io_in_d_0(b_1735_0),
		.io_in_control_0_dataflow(mesh_7_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2759_0),
		.io_in_last_0(r_3783_0),
		.io_in_valid_0(r_1735_0),
		.io_out_a_0(_mesh_7_22_io_out_a_0),
		.io_out_c_0(_mesh_7_22_io_out_c_0),
		.io_out_b_0(_mesh_7_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_22_io_out_id_0),
		.io_out_last_0(_mesh_7_22_io_out_last_0),
		.io_out_valid_0(_mesh_7_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9617 == GlobalFiModInstNr[0]) || (9617 == GlobalFiModInstNr[1]) || (9617 == GlobalFiModInstNr[2]) || (9617 == GlobalFiModInstNr[3]))));
	Tile mesh_7_23(
		.clock(clock),
		.io_in_a_0(r_247_0),
		.io_in_b_0(b_743_0),
		.io_in_d_0(b_1767_0),
		.io_in_control_0_dataflow(mesh_7_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2791_0),
		.io_in_last_0(r_3815_0),
		.io_in_valid_0(r_1767_0),
		.io_out_a_0(_mesh_7_23_io_out_a_0),
		.io_out_c_0(_mesh_7_23_io_out_c_0),
		.io_out_b_0(_mesh_7_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_23_io_out_id_0),
		.io_out_last_0(_mesh_7_23_io_out_last_0),
		.io_out_valid_0(_mesh_7_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9618 == GlobalFiModInstNr[0]) || (9618 == GlobalFiModInstNr[1]) || (9618 == GlobalFiModInstNr[2]) || (9618 == GlobalFiModInstNr[3]))));
	Tile mesh_7_24(
		.clock(clock),
		.io_in_a_0(r_248_0),
		.io_in_b_0(b_775_0),
		.io_in_d_0(b_1799_0),
		.io_in_control_0_dataflow(mesh_7_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2823_0),
		.io_in_last_0(r_3847_0),
		.io_in_valid_0(r_1799_0),
		.io_out_a_0(_mesh_7_24_io_out_a_0),
		.io_out_c_0(_mesh_7_24_io_out_c_0),
		.io_out_b_0(_mesh_7_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_24_io_out_id_0),
		.io_out_last_0(_mesh_7_24_io_out_last_0),
		.io_out_valid_0(_mesh_7_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9619 == GlobalFiModInstNr[0]) || (9619 == GlobalFiModInstNr[1]) || (9619 == GlobalFiModInstNr[2]) || (9619 == GlobalFiModInstNr[3]))));
	Tile mesh_7_25(
		.clock(clock),
		.io_in_a_0(r_249_0),
		.io_in_b_0(b_807_0),
		.io_in_d_0(b_1831_0),
		.io_in_control_0_dataflow(mesh_7_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2855_0),
		.io_in_last_0(r_3879_0),
		.io_in_valid_0(r_1831_0),
		.io_out_a_0(_mesh_7_25_io_out_a_0),
		.io_out_c_0(_mesh_7_25_io_out_c_0),
		.io_out_b_0(_mesh_7_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_25_io_out_id_0),
		.io_out_last_0(_mesh_7_25_io_out_last_0),
		.io_out_valid_0(_mesh_7_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9620 == GlobalFiModInstNr[0]) || (9620 == GlobalFiModInstNr[1]) || (9620 == GlobalFiModInstNr[2]) || (9620 == GlobalFiModInstNr[3]))));
	Tile mesh_7_26(
		.clock(clock),
		.io_in_a_0(r_250_0),
		.io_in_b_0(b_839_0),
		.io_in_d_0(b_1863_0),
		.io_in_control_0_dataflow(mesh_7_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2887_0),
		.io_in_last_0(r_3911_0),
		.io_in_valid_0(r_1863_0),
		.io_out_a_0(_mesh_7_26_io_out_a_0),
		.io_out_c_0(_mesh_7_26_io_out_c_0),
		.io_out_b_0(_mesh_7_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_26_io_out_id_0),
		.io_out_last_0(_mesh_7_26_io_out_last_0),
		.io_out_valid_0(_mesh_7_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9621 == GlobalFiModInstNr[0]) || (9621 == GlobalFiModInstNr[1]) || (9621 == GlobalFiModInstNr[2]) || (9621 == GlobalFiModInstNr[3]))));
	Tile mesh_7_27(
		.clock(clock),
		.io_in_a_0(r_251_0),
		.io_in_b_0(b_871_0),
		.io_in_d_0(b_1895_0),
		.io_in_control_0_dataflow(mesh_7_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2919_0),
		.io_in_last_0(r_3943_0),
		.io_in_valid_0(r_1895_0),
		.io_out_a_0(_mesh_7_27_io_out_a_0),
		.io_out_c_0(_mesh_7_27_io_out_c_0),
		.io_out_b_0(_mesh_7_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_27_io_out_id_0),
		.io_out_last_0(_mesh_7_27_io_out_last_0),
		.io_out_valid_0(_mesh_7_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9622 == GlobalFiModInstNr[0]) || (9622 == GlobalFiModInstNr[1]) || (9622 == GlobalFiModInstNr[2]) || (9622 == GlobalFiModInstNr[3]))));
	Tile mesh_7_28(
		.clock(clock),
		.io_in_a_0(r_252_0),
		.io_in_b_0(b_903_0),
		.io_in_d_0(b_1927_0),
		.io_in_control_0_dataflow(mesh_7_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2951_0),
		.io_in_last_0(r_3975_0),
		.io_in_valid_0(r_1927_0),
		.io_out_a_0(_mesh_7_28_io_out_a_0),
		.io_out_c_0(_mesh_7_28_io_out_c_0),
		.io_out_b_0(_mesh_7_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_28_io_out_id_0),
		.io_out_last_0(_mesh_7_28_io_out_last_0),
		.io_out_valid_0(_mesh_7_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9623 == GlobalFiModInstNr[0]) || (9623 == GlobalFiModInstNr[1]) || (9623 == GlobalFiModInstNr[2]) || (9623 == GlobalFiModInstNr[3]))));
	Tile mesh_7_29(
		.clock(clock),
		.io_in_a_0(r_253_0),
		.io_in_b_0(b_935_0),
		.io_in_d_0(b_1959_0),
		.io_in_control_0_dataflow(mesh_7_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2983_0),
		.io_in_last_0(r_4007_0),
		.io_in_valid_0(r_1959_0),
		.io_out_a_0(_mesh_7_29_io_out_a_0),
		.io_out_c_0(_mesh_7_29_io_out_c_0),
		.io_out_b_0(_mesh_7_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_29_io_out_id_0),
		.io_out_last_0(_mesh_7_29_io_out_last_0),
		.io_out_valid_0(_mesh_7_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9624 == GlobalFiModInstNr[0]) || (9624 == GlobalFiModInstNr[1]) || (9624 == GlobalFiModInstNr[2]) || (9624 == GlobalFiModInstNr[3]))));
	Tile mesh_7_30(
		.clock(clock),
		.io_in_a_0(r_254_0),
		.io_in_b_0(b_967_0),
		.io_in_d_0(b_1991_0),
		.io_in_control_0_dataflow(mesh_7_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3015_0),
		.io_in_last_0(r_4039_0),
		.io_in_valid_0(r_1991_0),
		.io_out_a_0(_mesh_7_30_io_out_a_0),
		.io_out_c_0(_mesh_7_30_io_out_c_0),
		.io_out_b_0(_mesh_7_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_30_io_out_id_0),
		.io_out_last_0(_mesh_7_30_io_out_last_0),
		.io_out_valid_0(_mesh_7_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9625 == GlobalFiModInstNr[0]) || (9625 == GlobalFiModInstNr[1]) || (9625 == GlobalFiModInstNr[2]) || (9625 == GlobalFiModInstNr[3]))));
	Tile mesh_7_31(
		.clock(clock),
		.io_in_a_0(r_255_0),
		.io_in_b_0(b_999_0),
		.io_in_d_0(b_2023_0),
		.io_in_control_0_dataflow(mesh_7_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3047_0),
		.io_in_last_0(r_4071_0),
		.io_in_valid_0(r_2023_0),
		.io_out_a_0(_mesh_7_31_io_out_a_0),
		.io_out_c_0(_mesh_7_31_io_out_c_0),
		.io_out_b_0(_mesh_7_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_31_io_out_id_0),
		.io_out_last_0(_mesh_7_31_io_out_last_0),
		.io_out_valid_0(_mesh_7_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9626 == GlobalFiModInstNr[0]) || (9626 == GlobalFiModInstNr[1]) || (9626 == GlobalFiModInstNr[2]) || (9626 == GlobalFiModInstNr[3]))));
	Tile mesh_8_0(
		.clock(clock),
		.io_in_a_0(r_256_0),
		.io_in_b_0(b_8_0),
		.io_in_d_0(b_1032_0),
		.io_in_control_0_dataflow(mesh_8_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2056_0),
		.io_in_last_0(r_3080_0),
		.io_in_valid_0(r_1032_0),
		.io_out_a_0(_mesh_8_0_io_out_a_0),
		.io_out_c_0(_mesh_8_0_io_out_c_0),
		.io_out_b_0(_mesh_8_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_0_io_out_id_0),
		.io_out_last_0(_mesh_8_0_io_out_last_0),
		.io_out_valid_0(_mesh_8_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9627 == GlobalFiModInstNr[0]) || (9627 == GlobalFiModInstNr[1]) || (9627 == GlobalFiModInstNr[2]) || (9627 == GlobalFiModInstNr[3]))));
	Tile mesh_8_1(
		.clock(clock),
		.io_in_a_0(r_257_0),
		.io_in_b_0(b_40_0),
		.io_in_d_0(b_1064_0),
		.io_in_control_0_dataflow(mesh_8_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2088_0),
		.io_in_last_0(r_3112_0),
		.io_in_valid_0(r_1064_0),
		.io_out_a_0(_mesh_8_1_io_out_a_0),
		.io_out_c_0(_mesh_8_1_io_out_c_0),
		.io_out_b_0(_mesh_8_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_1_io_out_id_0),
		.io_out_last_0(_mesh_8_1_io_out_last_0),
		.io_out_valid_0(_mesh_8_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9628 == GlobalFiModInstNr[0]) || (9628 == GlobalFiModInstNr[1]) || (9628 == GlobalFiModInstNr[2]) || (9628 == GlobalFiModInstNr[3]))));
	Tile mesh_8_2(
		.clock(clock),
		.io_in_a_0(r_258_0),
		.io_in_b_0(b_72_0),
		.io_in_d_0(b_1096_0),
		.io_in_control_0_dataflow(mesh_8_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2120_0),
		.io_in_last_0(r_3144_0),
		.io_in_valid_0(r_1096_0),
		.io_out_a_0(_mesh_8_2_io_out_a_0),
		.io_out_c_0(_mesh_8_2_io_out_c_0),
		.io_out_b_0(_mesh_8_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_2_io_out_id_0),
		.io_out_last_0(_mesh_8_2_io_out_last_0),
		.io_out_valid_0(_mesh_8_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9629 == GlobalFiModInstNr[0]) || (9629 == GlobalFiModInstNr[1]) || (9629 == GlobalFiModInstNr[2]) || (9629 == GlobalFiModInstNr[3]))));
	Tile mesh_8_3(
		.clock(clock),
		.io_in_a_0(r_259_0),
		.io_in_b_0(b_104_0),
		.io_in_d_0(b_1128_0),
		.io_in_control_0_dataflow(mesh_8_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2152_0),
		.io_in_last_0(r_3176_0),
		.io_in_valid_0(r_1128_0),
		.io_out_a_0(_mesh_8_3_io_out_a_0),
		.io_out_c_0(_mesh_8_3_io_out_c_0),
		.io_out_b_0(_mesh_8_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_3_io_out_id_0),
		.io_out_last_0(_mesh_8_3_io_out_last_0),
		.io_out_valid_0(_mesh_8_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9630 == GlobalFiModInstNr[0]) || (9630 == GlobalFiModInstNr[1]) || (9630 == GlobalFiModInstNr[2]) || (9630 == GlobalFiModInstNr[3]))));
	Tile mesh_8_4(
		.clock(clock),
		.io_in_a_0(r_260_0),
		.io_in_b_0(b_136_0),
		.io_in_d_0(b_1160_0),
		.io_in_control_0_dataflow(mesh_8_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2184_0),
		.io_in_last_0(r_3208_0),
		.io_in_valid_0(r_1160_0),
		.io_out_a_0(_mesh_8_4_io_out_a_0),
		.io_out_c_0(_mesh_8_4_io_out_c_0),
		.io_out_b_0(_mesh_8_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_4_io_out_id_0),
		.io_out_last_0(_mesh_8_4_io_out_last_0),
		.io_out_valid_0(_mesh_8_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9631 == GlobalFiModInstNr[0]) || (9631 == GlobalFiModInstNr[1]) || (9631 == GlobalFiModInstNr[2]) || (9631 == GlobalFiModInstNr[3]))));
	Tile mesh_8_5(
		.clock(clock),
		.io_in_a_0(r_261_0),
		.io_in_b_0(b_168_0),
		.io_in_d_0(b_1192_0),
		.io_in_control_0_dataflow(mesh_8_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2216_0),
		.io_in_last_0(r_3240_0),
		.io_in_valid_0(r_1192_0),
		.io_out_a_0(_mesh_8_5_io_out_a_0),
		.io_out_c_0(_mesh_8_5_io_out_c_0),
		.io_out_b_0(_mesh_8_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_5_io_out_id_0),
		.io_out_last_0(_mesh_8_5_io_out_last_0),
		.io_out_valid_0(_mesh_8_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9632 == GlobalFiModInstNr[0]) || (9632 == GlobalFiModInstNr[1]) || (9632 == GlobalFiModInstNr[2]) || (9632 == GlobalFiModInstNr[3]))));
	Tile mesh_8_6(
		.clock(clock),
		.io_in_a_0(r_262_0),
		.io_in_b_0(b_200_0),
		.io_in_d_0(b_1224_0),
		.io_in_control_0_dataflow(mesh_8_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2248_0),
		.io_in_last_0(r_3272_0),
		.io_in_valid_0(r_1224_0),
		.io_out_a_0(_mesh_8_6_io_out_a_0),
		.io_out_c_0(_mesh_8_6_io_out_c_0),
		.io_out_b_0(_mesh_8_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_6_io_out_id_0),
		.io_out_last_0(_mesh_8_6_io_out_last_0),
		.io_out_valid_0(_mesh_8_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9633 == GlobalFiModInstNr[0]) || (9633 == GlobalFiModInstNr[1]) || (9633 == GlobalFiModInstNr[2]) || (9633 == GlobalFiModInstNr[3]))));
	Tile mesh_8_7(
		.clock(clock),
		.io_in_a_0(r_263_0),
		.io_in_b_0(b_232_0),
		.io_in_d_0(b_1256_0),
		.io_in_control_0_dataflow(mesh_8_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2280_0),
		.io_in_last_0(r_3304_0),
		.io_in_valid_0(r_1256_0),
		.io_out_a_0(_mesh_8_7_io_out_a_0),
		.io_out_c_0(_mesh_8_7_io_out_c_0),
		.io_out_b_0(_mesh_8_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_7_io_out_id_0),
		.io_out_last_0(_mesh_8_7_io_out_last_0),
		.io_out_valid_0(_mesh_8_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9634 == GlobalFiModInstNr[0]) || (9634 == GlobalFiModInstNr[1]) || (9634 == GlobalFiModInstNr[2]) || (9634 == GlobalFiModInstNr[3]))));
	Tile mesh_8_8(
		.clock(clock),
		.io_in_a_0(r_264_0),
		.io_in_b_0(b_264_0),
		.io_in_d_0(b_1288_0),
		.io_in_control_0_dataflow(mesh_8_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2312_0),
		.io_in_last_0(r_3336_0),
		.io_in_valid_0(r_1288_0),
		.io_out_a_0(_mesh_8_8_io_out_a_0),
		.io_out_c_0(_mesh_8_8_io_out_c_0),
		.io_out_b_0(_mesh_8_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_8_io_out_id_0),
		.io_out_last_0(_mesh_8_8_io_out_last_0),
		.io_out_valid_0(_mesh_8_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9635 == GlobalFiModInstNr[0]) || (9635 == GlobalFiModInstNr[1]) || (9635 == GlobalFiModInstNr[2]) || (9635 == GlobalFiModInstNr[3]))));
	Tile mesh_8_9(
		.clock(clock),
		.io_in_a_0(r_265_0),
		.io_in_b_0(b_296_0),
		.io_in_d_0(b_1320_0),
		.io_in_control_0_dataflow(mesh_8_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2344_0),
		.io_in_last_0(r_3368_0),
		.io_in_valid_0(r_1320_0),
		.io_out_a_0(_mesh_8_9_io_out_a_0),
		.io_out_c_0(_mesh_8_9_io_out_c_0),
		.io_out_b_0(_mesh_8_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_9_io_out_id_0),
		.io_out_last_0(_mesh_8_9_io_out_last_0),
		.io_out_valid_0(_mesh_8_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9636 == GlobalFiModInstNr[0]) || (9636 == GlobalFiModInstNr[1]) || (9636 == GlobalFiModInstNr[2]) || (9636 == GlobalFiModInstNr[3]))));
	Tile mesh_8_10(
		.clock(clock),
		.io_in_a_0(r_266_0),
		.io_in_b_0(b_328_0),
		.io_in_d_0(b_1352_0),
		.io_in_control_0_dataflow(mesh_8_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2376_0),
		.io_in_last_0(r_3400_0),
		.io_in_valid_0(r_1352_0),
		.io_out_a_0(_mesh_8_10_io_out_a_0),
		.io_out_c_0(_mesh_8_10_io_out_c_0),
		.io_out_b_0(_mesh_8_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_10_io_out_id_0),
		.io_out_last_0(_mesh_8_10_io_out_last_0),
		.io_out_valid_0(_mesh_8_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9637 == GlobalFiModInstNr[0]) || (9637 == GlobalFiModInstNr[1]) || (9637 == GlobalFiModInstNr[2]) || (9637 == GlobalFiModInstNr[3]))));
	Tile mesh_8_11(
		.clock(clock),
		.io_in_a_0(r_267_0),
		.io_in_b_0(b_360_0),
		.io_in_d_0(b_1384_0),
		.io_in_control_0_dataflow(mesh_8_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2408_0),
		.io_in_last_0(r_3432_0),
		.io_in_valid_0(r_1384_0),
		.io_out_a_0(_mesh_8_11_io_out_a_0),
		.io_out_c_0(_mesh_8_11_io_out_c_0),
		.io_out_b_0(_mesh_8_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_11_io_out_id_0),
		.io_out_last_0(_mesh_8_11_io_out_last_0),
		.io_out_valid_0(_mesh_8_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9638 == GlobalFiModInstNr[0]) || (9638 == GlobalFiModInstNr[1]) || (9638 == GlobalFiModInstNr[2]) || (9638 == GlobalFiModInstNr[3]))));
	Tile mesh_8_12(
		.clock(clock),
		.io_in_a_0(r_268_0),
		.io_in_b_0(b_392_0),
		.io_in_d_0(b_1416_0),
		.io_in_control_0_dataflow(mesh_8_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2440_0),
		.io_in_last_0(r_3464_0),
		.io_in_valid_0(r_1416_0),
		.io_out_a_0(_mesh_8_12_io_out_a_0),
		.io_out_c_0(_mesh_8_12_io_out_c_0),
		.io_out_b_0(_mesh_8_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_12_io_out_id_0),
		.io_out_last_0(_mesh_8_12_io_out_last_0),
		.io_out_valid_0(_mesh_8_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9639 == GlobalFiModInstNr[0]) || (9639 == GlobalFiModInstNr[1]) || (9639 == GlobalFiModInstNr[2]) || (9639 == GlobalFiModInstNr[3]))));
	Tile mesh_8_13(
		.clock(clock),
		.io_in_a_0(r_269_0),
		.io_in_b_0(b_424_0),
		.io_in_d_0(b_1448_0),
		.io_in_control_0_dataflow(mesh_8_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2472_0),
		.io_in_last_0(r_3496_0),
		.io_in_valid_0(r_1448_0),
		.io_out_a_0(_mesh_8_13_io_out_a_0),
		.io_out_c_0(_mesh_8_13_io_out_c_0),
		.io_out_b_0(_mesh_8_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_13_io_out_id_0),
		.io_out_last_0(_mesh_8_13_io_out_last_0),
		.io_out_valid_0(_mesh_8_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9640 == GlobalFiModInstNr[0]) || (9640 == GlobalFiModInstNr[1]) || (9640 == GlobalFiModInstNr[2]) || (9640 == GlobalFiModInstNr[3]))));
	Tile mesh_8_14(
		.clock(clock),
		.io_in_a_0(r_270_0),
		.io_in_b_0(b_456_0),
		.io_in_d_0(b_1480_0),
		.io_in_control_0_dataflow(mesh_8_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2504_0),
		.io_in_last_0(r_3528_0),
		.io_in_valid_0(r_1480_0),
		.io_out_a_0(_mesh_8_14_io_out_a_0),
		.io_out_c_0(_mesh_8_14_io_out_c_0),
		.io_out_b_0(_mesh_8_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_14_io_out_id_0),
		.io_out_last_0(_mesh_8_14_io_out_last_0),
		.io_out_valid_0(_mesh_8_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9641 == GlobalFiModInstNr[0]) || (9641 == GlobalFiModInstNr[1]) || (9641 == GlobalFiModInstNr[2]) || (9641 == GlobalFiModInstNr[3]))));
	Tile mesh_8_15(
		.clock(clock),
		.io_in_a_0(r_271_0),
		.io_in_b_0(b_488_0),
		.io_in_d_0(b_1512_0),
		.io_in_control_0_dataflow(mesh_8_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2536_0),
		.io_in_last_0(r_3560_0),
		.io_in_valid_0(r_1512_0),
		.io_out_a_0(_mesh_8_15_io_out_a_0),
		.io_out_c_0(_mesh_8_15_io_out_c_0),
		.io_out_b_0(_mesh_8_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_15_io_out_id_0),
		.io_out_last_0(_mesh_8_15_io_out_last_0),
		.io_out_valid_0(_mesh_8_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9642 == GlobalFiModInstNr[0]) || (9642 == GlobalFiModInstNr[1]) || (9642 == GlobalFiModInstNr[2]) || (9642 == GlobalFiModInstNr[3]))));
	Tile mesh_8_16(
		.clock(clock),
		.io_in_a_0(r_272_0),
		.io_in_b_0(b_520_0),
		.io_in_d_0(b_1544_0),
		.io_in_control_0_dataflow(mesh_8_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2568_0),
		.io_in_last_0(r_3592_0),
		.io_in_valid_0(r_1544_0),
		.io_out_a_0(_mesh_8_16_io_out_a_0),
		.io_out_c_0(_mesh_8_16_io_out_c_0),
		.io_out_b_0(_mesh_8_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_16_io_out_id_0),
		.io_out_last_0(_mesh_8_16_io_out_last_0),
		.io_out_valid_0(_mesh_8_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9643 == GlobalFiModInstNr[0]) || (9643 == GlobalFiModInstNr[1]) || (9643 == GlobalFiModInstNr[2]) || (9643 == GlobalFiModInstNr[3]))));
	Tile mesh_8_17(
		.clock(clock),
		.io_in_a_0(r_273_0),
		.io_in_b_0(b_552_0),
		.io_in_d_0(b_1576_0),
		.io_in_control_0_dataflow(mesh_8_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2600_0),
		.io_in_last_0(r_3624_0),
		.io_in_valid_0(r_1576_0),
		.io_out_a_0(_mesh_8_17_io_out_a_0),
		.io_out_c_0(_mesh_8_17_io_out_c_0),
		.io_out_b_0(_mesh_8_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_17_io_out_id_0),
		.io_out_last_0(_mesh_8_17_io_out_last_0),
		.io_out_valid_0(_mesh_8_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9644 == GlobalFiModInstNr[0]) || (9644 == GlobalFiModInstNr[1]) || (9644 == GlobalFiModInstNr[2]) || (9644 == GlobalFiModInstNr[3]))));
	Tile mesh_8_18(
		.clock(clock),
		.io_in_a_0(r_274_0),
		.io_in_b_0(b_584_0),
		.io_in_d_0(b_1608_0),
		.io_in_control_0_dataflow(mesh_8_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2632_0),
		.io_in_last_0(r_3656_0),
		.io_in_valid_0(r_1608_0),
		.io_out_a_0(_mesh_8_18_io_out_a_0),
		.io_out_c_0(_mesh_8_18_io_out_c_0),
		.io_out_b_0(_mesh_8_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_18_io_out_id_0),
		.io_out_last_0(_mesh_8_18_io_out_last_0),
		.io_out_valid_0(_mesh_8_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9645 == GlobalFiModInstNr[0]) || (9645 == GlobalFiModInstNr[1]) || (9645 == GlobalFiModInstNr[2]) || (9645 == GlobalFiModInstNr[3]))));
	Tile mesh_8_19(
		.clock(clock),
		.io_in_a_0(r_275_0),
		.io_in_b_0(b_616_0),
		.io_in_d_0(b_1640_0),
		.io_in_control_0_dataflow(mesh_8_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2664_0),
		.io_in_last_0(r_3688_0),
		.io_in_valid_0(r_1640_0),
		.io_out_a_0(_mesh_8_19_io_out_a_0),
		.io_out_c_0(_mesh_8_19_io_out_c_0),
		.io_out_b_0(_mesh_8_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_19_io_out_id_0),
		.io_out_last_0(_mesh_8_19_io_out_last_0),
		.io_out_valid_0(_mesh_8_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9646 == GlobalFiModInstNr[0]) || (9646 == GlobalFiModInstNr[1]) || (9646 == GlobalFiModInstNr[2]) || (9646 == GlobalFiModInstNr[3]))));
	Tile mesh_8_20(
		.clock(clock),
		.io_in_a_0(r_276_0),
		.io_in_b_0(b_648_0),
		.io_in_d_0(b_1672_0),
		.io_in_control_0_dataflow(mesh_8_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2696_0),
		.io_in_last_0(r_3720_0),
		.io_in_valid_0(r_1672_0),
		.io_out_a_0(_mesh_8_20_io_out_a_0),
		.io_out_c_0(_mesh_8_20_io_out_c_0),
		.io_out_b_0(_mesh_8_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_20_io_out_id_0),
		.io_out_last_0(_mesh_8_20_io_out_last_0),
		.io_out_valid_0(_mesh_8_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9647 == GlobalFiModInstNr[0]) || (9647 == GlobalFiModInstNr[1]) || (9647 == GlobalFiModInstNr[2]) || (9647 == GlobalFiModInstNr[3]))));
	Tile mesh_8_21(
		.clock(clock),
		.io_in_a_0(r_277_0),
		.io_in_b_0(b_680_0),
		.io_in_d_0(b_1704_0),
		.io_in_control_0_dataflow(mesh_8_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2728_0),
		.io_in_last_0(r_3752_0),
		.io_in_valid_0(r_1704_0),
		.io_out_a_0(_mesh_8_21_io_out_a_0),
		.io_out_c_0(_mesh_8_21_io_out_c_0),
		.io_out_b_0(_mesh_8_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_21_io_out_id_0),
		.io_out_last_0(_mesh_8_21_io_out_last_0),
		.io_out_valid_0(_mesh_8_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9648 == GlobalFiModInstNr[0]) || (9648 == GlobalFiModInstNr[1]) || (9648 == GlobalFiModInstNr[2]) || (9648 == GlobalFiModInstNr[3]))));
	Tile mesh_8_22(
		.clock(clock),
		.io_in_a_0(r_278_0),
		.io_in_b_0(b_712_0),
		.io_in_d_0(b_1736_0),
		.io_in_control_0_dataflow(mesh_8_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2760_0),
		.io_in_last_0(r_3784_0),
		.io_in_valid_0(r_1736_0),
		.io_out_a_0(_mesh_8_22_io_out_a_0),
		.io_out_c_0(_mesh_8_22_io_out_c_0),
		.io_out_b_0(_mesh_8_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_22_io_out_id_0),
		.io_out_last_0(_mesh_8_22_io_out_last_0),
		.io_out_valid_0(_mesh_8_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9649 == GlobalFiModInstNr[0]) || (9649 == GlobalFiModInstNr[1]) || (9649 == GlobalFiModInstNr[2]) || (9649 == GlobalFiModInstNr[3]))));
	Tile mesh_8_23(
		.clock(clock),
		.io_in_a_0(r_279_0),
		.io_in_b_0(b_744_0),
		.io_in_d_0(b_1768_0),
		.io_in_control_0_dataflow(mesh_8_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2792_0),
		.io_in_last_0(r_3816_0),
		.io_in_valid_0(r_1768_0),
		.io_out_a_0(_mesh_8_23_io_out_a_0),
		.io_out_c_0(_mesh_8_23_io_out_c_0),
		.io_out_b_0(_mesh_8_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_23_io_out_id_0),
		.io_out_last_0(_mesh_8_23_io_out_last_0),
		.io_out_valid_0(_mesh_8_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9650 == GlobalFiModInstNr[0]) || (9650 == GlobalFiModInstNr[1]) || (9650 == GlobalFiModInstNr[2]) || (9650 == GlobalFiModInstNr[3]))));
	Tile mesh_8_24(
		.clock(clock),
		.io_in_a_0(r_280_0),
		.io_in_b_0(b_776_0),
		.io_in_d_0(b_1800_0),
		.io_in_control_0_dataflow(mesh_8_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2824_0),
		.io_in_last_0(r_3848_0),
		.io_in_valid_0(r_1800_0),
		.io_out_a_0(_mesh_8_24_io_out_a_0),
		.io_out_c_0(_mesh_8_24_io_out_c_0),
		.io_out_b_0(_mesh_8_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_24_io_out_id_0),
		.io_out_last_0(_mesh_8_24_io_out_last_0),
		.io_out_valid_0(_mesh_8_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9651 == GlobalFiModInstNr[0]) || (9651 == GlobalFiModInstNr[1]) || (9651 == GlobalFiModInstNr[2]) || (9651 == GlobalFiModInstNr[3]))));
	Tile mesh_8_25(
		.clock(clock),
		.io_in_a_0(r_281_0),
		.io_in_b_0(b_808_0),
		.io_in_d_0(b_1832_0),
		.io_in_control_0_dataflow(mesh_8_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2856_0),
		.io_in_last_0(r_3880_0),
		.io_in_valid_0(r_1832_0),
		.io_out_a_0(_mesh_8_25_io_out_a_0),
		.io_out_c_0(_mesh_8_25_io_out_c_0),
		.io_out_b_0(_mesh_8_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_25_io_out_id_0),
		.io_out_last_0(_mesh_8_25_io_out_last_0),
		.io_out_valid_0(_mesh_8_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9652 == GlobalFiModInstNr[0]) || (9652 == GlobalFiModInstNr[1]) || (9652 == GlobalFiModInstNr[2]) || (9652 == GlobalFiModInstNr[3]))));
	Tile mesh_8_26(
		.clock(clock),
		.io_in_a_0(r_282_0),
		.io_in_b_0(b_840_0),
		.io_in_d_0(b_1864_0),
		.io_in_control_0_dataflow(mesh_8_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2888_0),
		.io_in_last_0(r_3912_0),
		.io_in_valid_0(r_1864_0),
		.io_out_a_0(_mesh_8_26_io_out_a_0),
		.io_out_c_0(_mesh_8_26_io_out_c_0),
		.io_out_b_0(_mesh_8_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_26_io_out_id_0),
		.io_out_last_0(_mesh_8_26_io_out_last_0),
		.io_out_valid_0(_mesh_8_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9653 == GlobalFiModInstNr[0]) || (9653 == GlobalFiModInstNr[1]) || (9653 == GlobalFiModInstNr[2]) || (9653 == GlobalFiModInstNr[3]))));
	Tile mesh_8_27(
		.clock(clock),
		.io_in_a_0(r_283_0),
		.io_in_b_0(b_872_0),
		.io_in_d_0(b_1896_0),
		.io_in_control_0_dataflow(mesh_8_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2920_0),
		.io_in_last_0(r_3944_0),
		.io_in_valid_0(r_1896_0),
		.io_out_a_0(_mesh_8_27_io_out_a_0),
		.io_out_c_0(_mesh_8_27_io_out_c_0),
		.io_out_b_0(_mesh_8_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_27_io_out_id_0),
		.io_out_last_0(_mesh_8_27_io_out_last_0),
		.io_out_valid_0(_mesh_8_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9654 == GlobalFiModInstNr[0]) || (9654 == GlobalFiModInstNr[1]) || (9654 == GlobalFiModInstNr[2]) || (9654 == GlobalFiModInstNr[3]))));
	Tile mesh_8_28(
		.clock(clock),
		.io_in_a_0(r_284_0),
		.io_in_b_0(b_904_0),
		.io_in_d_0(b_1928_0),
		.io_in_control_0_dataflow(mesh_8_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2952_0),
		.io_in_last_0(r_3976_0),
		.io_in_valid_0(r_1928_0),
		.io_out_a_0(_mesh_8_28_io_out_a_0),
		.io_out_c_0(_mesh_8_28_io_out_c_0),
		.io_out_b_0(_mesh_8_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_28_io_out_id_0),
		.io_out_last_0(_mesh_8_28_io_out_last_0),
		.io_out_valid_0(_mesh_8_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9655 == GlobalFiModInstNr[0]) || (9655 == GlobalFiModInstNr[1]) || (9655 == GlobalFiModInstNr[2]) || (9655 == GlobalFiModInstNr[3]))));
	Tile mesh_8_29(
		.clock(clock),
		.io_in_a_0(r_285_0),
		.io_in_b_0(b_936_0),
		.io_in_d_0(b_1960_0),
		.io_in_control_0_dataflow(mesh_8_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2984_0),
		.io_in_last_0(r_4008_0),
		.io_in_valid_0(r_1960_0),
		.io_out_a_0(_mesh_8_29_io_out_a_0),
		.io_out_c_0(_mesh_8_29_io_out_c_0),
		.io_out_b_0(_mesh_8_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_29_io_out_id_0),
		.io_out_last_0(_mesh_8_29_io_out_last_0),
		.io_out_valid_0(_mesh_8_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9656 == GlobalFiModInstNr[0]) || (9656 == GlobalFiModInstNr[1]) || (9656 == GlobalFiModInstNr[2]) || (9656 == GlobalFiModInstNr[3]))));
	Tile mesh_8_30(
		.clock(clock),
		.io_in_a_0(r_286_0),
		.io_in_b_0(b_968_0),
		.io_in_d_0(b_1992_0),
		.io_in_control_0_dataflow(mesh_8_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3016_0),
		.io_in_last_0(r_4040_0),
		.io_in_valid_0(r_1992_0),
		.io_out_a_0(_mesh_8_30_io_out_a_0),
		.io_out_c_0(_mesh_8_30_io_out_c_0),
		.io_out_b_0(_mesh_8_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_30_io_out_id_0),
		.io_out_last_0(_mesh_8_30_io_out_last_0),
		.io_out_valid_0(_mesh_8_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9657 == GlobalFiModInstNr[0]) || (9657 == GlobalFiModInstNr[1]) || (9657 == GlobalFiModInstNr[2]) || (9657 == GlobalFiModInstNr[3]))));
	Tile mesh_8_31(
		.clock(clock),
		.io_in_a_0(r_287_0),
		.io_in_b_0(b_1000_0),
		.io_in_d_0(b_2024_0),
		.io_in_control_0_dataflow(mesh_8_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_8_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_8_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3048_0),
		.io_in_last_0(r_4072_0),
		.io_in_valid_0(r_2024_0),
		.io_out_a_0(_mesh_8_31_io_out_a_0),
		.io_out_c_0(_mesh_8_31_io_out_c_0),
		.io_out_b_0(_mesh_8_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_8_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_8_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_8_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_8_31_io_out_id_0),
		.io_out_last_0(_mesh_8_31_io_out_last_0),
		.io_out_valid_0(_mesh_8_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9658 == GlobalFiModInstNr[0]) || (9658 == GlobalFiModInstNr[1]) || (9658 == GlobalFiModInstNr[2]) || (9658 == GlobalFiModInstNr[3]))));
	Tile mesh_9_0(
		.clock(clock),
		.io_in_a_0(r_288_0),
		.io_in_b_0(b_9_0),
		.io_in_d_0(b_1033_0),
		.io_in_control_0_dataflow(mesh_9_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2057_0),
		.io_in_last_0(r_3081_0),
		.io_in_valid_0(r_1033_0),
		.io_out_a_0(_mesh_9_0_io_out_a_0),
		.io_out_c_0(_mesh_9_0_io_out_c_0),
		.io_out_b_0(_mesh_9_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_0_io_out_id_0),
		.io_out_last_0(_mesh_9_0_io_out_last_0),
		.io_out_valid_0(_mesh_9_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9659 == GlobalFiModInstNr[0]) || (9659 == GlobalFiModInstNr[1]) || (9659 == GlobalFiModInstNr[2]) || (9659 == GlobalFiModInstNr[3]))));
	Tile mesh_9_1(
		.clock(clock),
		.io_in_a_0(r_289_0),
		.io_in_b_0(b_41_0),
		.io_in_d_0(b_1065_0),
		.io_in_control_0_dataflow(mesh_9_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2089_0),
		.io_in_last_0(r_3113_0),
		.io_in_valid_0(r_1065_0),
		.io_out_a_0(_mesh_9_1_io_out_a_0),
		.io_out_c_0(_mesh_9_1_io_out_c_0),
		.io_out_b_0(_mesh_9_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_1_io_out_id_0),
		.io_out_last_0(_mesh_9_1_io_out_last_0),
		.io_out_valid_0(_mesh_9_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9660 == GlobalFiModInstNr[0]) || (9660 == GlobalFiModInstNr[1]) || (9660 == GlobalFiModInstNr[2]) || (9660 == GlobalFiModInstNr[3]))));
	Tile mesh_9_2(
		.clock(clock),
		.io_in_a_0(r_290_0),
		.io_in_b_0(b_73_0),
		.io_in_d_0(b_1097_0),
		.io_in_control_0_dataflow(mesh_9_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2121_0),
		.io_in_last_0(r_3145_0),
		.io_in_valid_0(r_1097_0),
		.io_out_a_0(_mesh_9_2_io_out_a_0),
		.io_out_c_0(_mesh_9_2_io_out_c_0),
		.io_out_b_0(_mesh_9_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_2_io_out_id_0),
		.io_out_last_0(_mesh_9_2_io_out_last_0),
		.io_out_valid_0(_mesh_9_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9661 == GlobalFiModInstNr[0]) || (9661 == GlobalFiModInstNr[1]) || (9661 == GlobalFiModInstNr[2]) || (9661 == GlobalFiModInstNr[3]))));
	Tile mesh_9_3(
		.clock(clock),
		.io_in_a_0(r_291_0),
		.io_in_b_0(b_105_0),
		.io_in_d_0(b_1129_0),
		.io_in_control_0_dataflow(mesh_9_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2153_0),
		.io_in_last_0(r_3177_0),
		.io_in_valid_0(r_1129_0),
		.io_out_a_0(_mesh_9_3_io_out_a_0),
		.io_out_c_0(_mesh_9_3_io_out_c_0),
		.io_out_b_0(_mesh_9_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_3_io_out_id_0),
		.io_out_last_0(_mesh_9_3_io_out_last_0),
		.io_out_valid_0(_mesh_9_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9662 == GlobalFiModInstNr[0]) || (9662 == GlobalFiModInstNr[1]) || (9662 == GlobalFiModInstNr[2]) || (9662 == GlobalFiModInstNr[3]))));
	Tile mesh_9_4(
		.clock(clock),
		.io_in_a_0(r_292_0),
		.io_in_b_0(b_137_0),
		.io_in_d_0(b_1161_0),
		.io_in_control_0_dataflow(mesh_9_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2185_0),
		.io_in_last_0(r_3209_0),
		.io_in_valid_0(r_1161_0),
		.io_out_a_0(_mesh_9_4_io_out_a_0),
		.io_out_c_0(_mesh_9_4_io_out_c_0),
		.io_out_b_0(_mesh_9_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_4_io_out_id_0),
		.io_out_last_0(_mesh_9_4_io_out_last_0),
		.io_out_valid_0(_mesh_9_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9663 == GlobalFiModInstNr[0]) || (9663 == GlobalFiModInstNr[1]) || (9663 == GlobalFiModInstNr[2]) || (9663 == GlobalFiModInstNr[3]))));
	Tile mesh_9_5(
		.clock(clock),
		.io_in_a_0(r_293_0),
		.io_in_b_0(b_169_0),
		.io_in_d_0(b_1193_0),
		.io_in_control_0_dataflow(mesh_9_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2217_0),
		.io_in_last_0(r_3241_0),
		.io_in_valid_0(r_1193_0),
		.io_out_a_0(_mesh_9_5_io_out_a_0),
		.io_out_c_0(_mesh_9_5_io_out_c_0),
		.io_out_b_0(_mesh_9_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_5_io_out_id_0),
		.io_out_last_0(_mesh_9_5_io_out_last_0),
		.io_out_valid_0(_mesh_9_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9664 == GlobalFiModInstNr[0]) || (9664 == GlobalFiModInstNr[1]) || (9664 == GlobalFiModInstNr[2]) || (9664 == GlobalFiModInstNr[3]))));
	Tile mesh_9_6(
		.clock(clock),
		.io_in_a_0(r_294_0),
		.io_in_b_0(b_201_0),
		.io_in_d_0(b_1225_0),
		.io_in_control_0_dataflow(mesh_9_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2249_0),
		.io_in_last_0(r_3273_0),
		.io_in_valid_0(r_1225_0),
		.io_out_a_0(_mesh_9_6_io_out_a_0),
		.io_out_c_0(_mesh_9_6_io_out_c_0),
		.io_out_b_0(_mesh_9_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_6_io_out_id_0),
		.io_out_last_0(_mesh_9_6_io_out_last_0),
		.io_out_valid_0(_mesh_9_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9665 == GlobalFiModInstNr[0]) || (9665 == GlobalFiModInstNr[1]) || (9665 == GlobalFiModInstNr[2]) || (9665 == GlobalFiModInstNr[3]))));
	Tile mesh_9_7(
		.clock(clock),
		.io_in_a_0(r_295_0),
		.io_in_b_0(b_233_0),
		.io_in_d_0(b_1257_0),
		.io_in_control_0_dataflow(mesh_9_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2281_0),
		.io_in_last_0(r_3305_0),
		.io_in_valid_0(r_1257_0),
		.io_out_a_0(_mesh_9_7_io_out_a_0),
		.io_out_c_0(_mesh_9_7_io_out_c_0),
		.io_out_b_0(_mesh_9_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_7_io_out_id_0),
		.io_out_last_0(_mesh_9_7_io_out_last_0),
		.io_out_valid_0(_mesh_9_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9666 == GlobalFiModInstNr[0]) || (9666 == GlobalFiModInstNr[1]) || (9666 == GlobalFiModInstNr[2]) || (9666 == GlobalFiModInstNr[3]))));
	Tile mesh_9_8(
		.clock(clock),
		.io_in_a_0(r_296_0),
		.io_in_b_0(b_265_0),
		.io_in_d_0(b_1289_0),
		.io_in_control_0_dataflow(mesh_9_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2313_0),
		.io_in_last_0(r_3337_0),
		.io_in_valid_0(r_1289_0),
		.io_out_a_0(_mesh_9_8_io_out_a_0),
		.io_out_c_0(_mesh_9_8_io_out_c_0),
		.io_out_b_0(_mesh_9_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_8_io_out_id_0),
		.io_out_last_0(_mesh_9_8_io_out_last_0),
		.io_out_valid_0(_mesh_9_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9667 == GlobalFiModInstNr[0]) || (9667 == GlobalFiModInstNr[1]) || (9667 == GlobalFiModInstNr[2]) || (9667 == GlobalFiModInstNr[3]))));
	Tile mesh_9_9(
		.clock(clock),
		.io_in_a_0(r_297_0),
		.io_in_b_0(b_297_0),
		.io_in_d_0(b_1321_0),
		.io_in_control_0_dataflow(mesh_9_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2345_0),
		.io_in_last_0(r_3369_0),
		.io_in_valid_0(r_1321_0),
		.io_out_a_0(_mesh_9_9_io_out_a_0),
		.io_out_c_0(_mesh_9_9_io_out_c_0),
		.io_out_b_0(_mesh_9_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_9_io_out_id_0),
		.io_out_last_0(_mesh_9_9_io_out_last_0),
		.io_out_valid_0(_mesh_9_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9668 == GlobalFiModInstNr[0]) || (9668 == GlobalFiModInstNr[1]) || (9668 == GlobalFiModInstNr[2]) || (9668 == GlobalFiModInstNr[3]))));
	Tile mesh_9_10(
		.clock(clock),
		.io_in_a_0(r_298_0),
		.io_in_b_0(b_329_0),
		.io_in_d_0(b_1353_0),
		.io_in_control_0_dataflow(mesh_9_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2377_0),
		.io_in_last_0(r_3401_0),
		.io_in_valid_0(r_1353_0),
		.io_out_a_0(_mesh_9_10_io_out_a_0),
		.io_out_c_0(_mesh_9_10_io_out_c_0),
		.io_out_b_0(_mesh_9_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_10_io_out_id_0),
		.io_out_last_0(_mesh_9_10_io_out_last_0),
		.io_out_valid_0(_mesh_9_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9669 == GlobalFiModInstNr[0]) || (9669 == GlobalFiModInstNr[1]) || (9669 == GlobalFiModInstNr[2]) || (9669 == GlobalFiModInstNr[3]))));
	Tile mesh_9_11(
		.clock(clock),
		.io_in_a_0(r_299_0),
		.io_in_b_0(b_361_0),
		.io_in_d_0(b_1385_0),
		.io_in_control_0_dataflow(mesh_9_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2409_0),
		.io_in_last_0(r_3433_0),
		.io_in_valid_0(r_1385_0),
		.io_out_a_0(_mesh_9_11_io_out_a_0),
		.io_out_c_0(_mesh_9_11_io_out_c_0),
		.io_out_b_0(_mesh_9_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_11_io_out_id_0),
		.io_out_last_0(_mesh_9_11_io_out_last_0),
		.io_out_valid_0(_mesh_9_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9670 == GlobalFiModInstNr[0]) || (9670 == GlobalFiModInstNr[1]) || (9670 == GlobalFiModInstNr[2]) || (9670 == GlobalFiModInstNr[3]))));
	Tile mesh_9_12(
		.clock(clock),
		.io_in_a_0(r_300_0),
		.io_in_b_0(b_393_0),
		.io_in_d_0(b_1417_0),
		.io_in_control_0_dataflow(mesh_9_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2441_0),
		.io_in_last_0(r_3465_0),
		.io_in_valid_0(r_1417_0),
		.io_out_a_0(_mesh_9_12_io_out_a_0),
		.io_out_c_0(_mesh_9_12_io_out_c_0),
		.io_out_b_0(_mesh_9_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_12_io_out_id_0),
		.io_out_last_0(_mesh_9_12_io_out_last_0),
		.io_out_valid_0(_mesh_9_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9671 == GlobalFiModInstNr[0]) || (9671 == GlobalFiModInstNr[1]) || (9671 == GlobalFiModInstNr[2]) || (9671 == GlobalFiModInstNr[3]))));
	Tile mesh_9_13(
		.clock(clock),
		.io_in_a_0(r_301_0),
		.io_in_b_0(b_425_0),
		.io_in_d_0(b_1449_0),
		.io_in_control_0_dataflow(mesh_9_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2473_0),
		.io_in_last_0(r_3497_0),
		.io_in_valid_0(r_1449_0),
		.io_out_a_0(_mesh_9_13_io_out_a_0),
		.io_out_c_0(_mesh_9_13_io_out_c_0),
		.io_out_b_0(_mesh_9_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_13_io_out_id_0),
		.io_out_last_0(_mesh_9_13_io_out_last_0),
		.io_out_valid_0(_mesh_9_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9672 == GlobalFiModInstNr[0]) || (9672 == GlobalFiModInstNr[1]) || (9672 == GlobalFiModInstNr[2]) || (9672 == GlobalFiModInstNr[3]))));
	Tile mesh_9_14(
		.clock(clock),
		.io_in_a_0(r_302_0),
		.io_in_b_0(b_457_0),
		.io_in_d_0(b_1481_0),
		.io_in_control_0_dataflow(mesh_9_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2505_0),
		.io_in_last_0(r_3529_0),
		.io_in_valid_0(r_1481_0),
		.io_out_a_0(_mesh_9_14_io_out_a_0),
		.io_out_c_0(_mesh_9_14_io_out_c_0),
		.io_out_b_0(_mesh_9_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_14_io_out_id_0),
		.io_out_last_0(_mesh_9_14_io_out_last_0),
		.io_out_valid_0(_mesh_9_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9673 == GlobalFiModInstNr[0]) || (9673 == GlobalFiModInstNr[1]) || (9673 == GlobalFiModInstNr[2]) || (9673 == GlobalFiModInstNr[3]))));
	Tile mesh_9_15(
		.clock(clock),
		.io_in_a_0(r_303_0),
		.io_in_b_0(b_489_0),
		.io_in_d_0(b_1513_0),
		.io_in_control_0_dataflow(mesh_9_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2537_0),
		.io_in_last_0(r_3561_0),
		.io_in_valid_0(r_1513_0),
		.io_out_a_0(_mesh_9_15_io_out_a_0),
		.io_out_c_0(_mesh_9_15_io_out_c_0),
		.io_out_b_0(_mesh_9_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_15_io_out_id_0),
		.io_out_last_0(_mesh_9_15_io_out_last_0),
		.io_out_valid_0(_mesh_9_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9674 == GlobalFiModInstNr[0]) || (9674 == GlobalFiModInstNr[1]) || (9674 == GlobalFiModInstNr[2]) || (9674 == GlobalFiModInstNr[3]))));
	Tile mesh_9_16(
		.clock(clock),
		.io_in_a_0(r_304_0),
		.io_in_b_0(b_521_0),
		.io_in_d_0(b_1545_0),
		.io_in_control_0_dataflow(mesh_9_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2569_0),
		.io_in_last_0(r_3593_0),
		.io_in_valid_0(r_1545_0),
		.io_out_a_0(_mesh_9_16_io_out_a_0),
		.io_out_c_0(_mesh_9_16_io_out_c_0),
		.io_out_b_0(_mesh_9_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_16_io_out_id_0),
		.io_out_last_0(_mesh_9_16_io_out_last_0),
		.io_out_valid_0(_mesh_9_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9675 == GlobalFiModInstNr[0]) || (9675 == GlobalFiModInstNr[1]) || (9675 == GlobalFiModInstNr[2]) || (9675 == GlobalFiModInstNr[3]))));
	Tile mesh_9_17(
		.clock(clock),
		.io_in_a_0(r_305_0),
		.io_in_b_0(b_553_0),
		.io_in_d_0(b_1577_0),
		.io_in_control_0_dataflow(mesh_9_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2601_0),
		.io_in_last_0(r_3625_0),
		.io_in_valid_0(r_1577_0),
		.io_out_a_0(_mesh_9_17_io_out_a_0),
		.io_out_c_0(_mesh_9_17_io_out_c_0),
		.io_out_b_0(_mesh_9_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_17_io_out_id_0),
		.io_out_last_0(_mesh_9_17_io_out_last_0),
		.io_out_valid_0(_mesh_9_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9676 == GlobalFiModInstNr[0]) || (9676 == GlobalFiModInstNr[1]) || (9676 == GlobalFiModInstNr[2]) || (9676 == GlobalFiModInstNr[3]))));
	Tile mesh_9_18(
		.clock(clock),
		.io_in_a_0(r_306_0),
		.io_in_b_0(b_585_0),
		.io_in_d_0(b_1609_0),
		.io_in_control_0_dataflow(mesh_9_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2633_0),
		.io_in_last_0(r_3657_0),
		.io_in_valid_0(r_1609_0),
		.io_out_a_0(_mesh_9_18_io_out_a_0),
		.io_out_c_0(_mesh_9_18_io_out_c_0),
		.io_out_b_0(_mesh_9_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_18_io_out_id_0),
		.io_out_last_0(_mesh_9_18_io_out_last_0),
		.io_out_valid_0(_mesh_9_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9677 == GlobalFiModInstNr[0]) || (9677 == GlobalFiModInstNr[1]) || (9677 == GlobalFiModInstNr[2]) || (9677 == GlobalFiModInstNr[3]))));
	Tile mesh_9_19(
		.clock(clock),
		.io_in_a_0(r_307_0),
		.io_in_b_0(b_617_0),
		.io_in_d_0(b_1641_0),
		.io_in_control_0_dataflow(mesh_9_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2665_0),
		.io_in_last_0(r_3689_0),
		.io_in_valid_0(r_1641_0),
		.io_out_a_0(_mesh_9_19_io_out_a_0),
		.io_out_c_0(_mesh_9_19_io_out_c_0),
		.io_out_b_0(_mesh_9_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_19_io_out_id_0),
		.io_out_last_0(_mesh_9_19_io_out_last_0),
		.io_out_valid_0(_mesh_9_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9678 == GlobalFiModInstNr[0]) || (9678 == GlobalFiModInstNr[1]) || (9678 == GlobalFiModInstNr[2]) || (9678 == GlobalFiModInstNr[3]))));
	Tile mesh_9_20(
		.clock(clock),
		.io_in_a_0(r_308_0),
		.io_in_b_0(b_649_0),
		.io_in_d_0(b_1673_0),
		.io_in_control_0_dataflow(mesh_9_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2697_0),
		.io_in_last_0(r_3721_0),
		.io_in_valid_0(r_1673_0),
		.io_out_a_0(_mesh_9_20_io_out_a_0),
		.io_out_c_0(_mesh_9_20_io_out_c_0),
		.io_out_b_0(_mesh_9_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_20_io_out_id_0),
		.io_out_last_0(_mesh_9_20_io_out_last_0),
		.io_out_valid_0(_mesh_9_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9679 == GlobalFiModInstNr[0]) || (9679 == GlobalFiModInstNr[1]) || (9679 == GlobalFiModInstNr[2]) || (9679 == GlobalFiModInstNr[3]))));
	Tile mesh_9_21(
		.clock(clock),
		.io_in_a_0(r_309_0),
		.io_in_b_0(b_681_0),
		.io_in_d_0(b_1705_0),
		.io_in_control_0_dataflow(mesh_9_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2729_0),
		.io_in_last_0(r_3753_0),
		.io_in_valid_0(r_1705_0),
		.io_out_a_0(_mesh_9_21_io_out_a_0),
		.io_out_c_0(_mesh_9_21_io_out_c_0),
		.io_out_b_0(_mesh_9_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_21_io_out_id_0),
		.io_out_last_0(_mesh_9_21_io_out_last_0),
		.io_out_valid_0(_mesh_9_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9680 == GlobalFiModInstNr[0]) || (9680 == GlobalFiModInstNr[1]) || (9680 == GlobalFiModInstNr[2]) || (9680 == GlobalFiModInstNr[3]))));
	Tile mesh_9_22(
		.clock(clock),
		.io_in_a_0(r_310_0),
		.io_in_b_0(b_713_0),
		.io_in_d_0(b_1737_0),
		.io_in_control_0_dataflow(mesh_9_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2761_0),
		.io_in_last_0(r_3785_0),
		.io_in_valid_0(r_1737_0),
		.io_out_a_0(_mesh_9_22_io_out_a_0),
		.io_out_c_0(_mesh_9_22_io_out_c_0),
		.io_out_b_0(_mesh_9_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_22_io_out_id_0),
		.io_out_last_0(_mesh_9_22_io_out_last_0),
		.io_out_valid_0(_mesh_9_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9681 == GlobalFiModInstNr[0]) || (9681 == GlobalFiModInstNr[1]) || (9681 == GlobalFiModInstNr[2]) || (9681 == GlobalFiModInstNr[3]))));
	Tile mesh_9_23(
		.clock(clock),
		.io_in_a_0(r_311_0),
		.io_in_b_0(b_745_0),
		.io_in_d_0(b_1769_0),
		.io_in_control_0_dataflow(mesh_9_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2793_0),
		.io_in_last_0(r_3817_0),
		.io_in_valid_0(r_1769_0),
		.io_out_a_0(_mesh_9_23_io_out_a_0),
		.io_out_c_0(_mesh_9_23_io_out_c_0),
		.io_out_b_0(_mesh_9_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_23_io_out_id_0),
		.io_out_last_0(_mesh_9_23_io_out_last_0),
		.io_out_valid_0(_mesh_9_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9682 == GlobalFiModInstNr[0]) || (9682 == GlobalFiModInstNr[1]) || (9682 == GlobalFiModInstNr[2]) || (9682 == GlobalFiModInstNr[3]))));
	Tile mesh_9_24(
		.clock(clock),
		.io_in_a_0(r_312_0),
		.io_in_b_0(b_777_0),
		.io_in_d_0(b_1801_0),
		.io_in_control_0_dataflow(mesh_9_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2825_0),
		.io_in_last_0(r_3849_0),
		.io_in_valid_0(r_1801_0),
		.io_out_a_0(_mesh_9_24_io_out_a_0),
		.io_out_c_0(_mesh_9_24_io_out_c_0),
		.io_out_b_0(_mesh_9_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_24_io_out_id_0),
		.io_out_last_0(_mesh_9_24_io_out_last_0),
		.io_out_valid_0(_mesh_9_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9683 == GlobalFiModInstNr[0]) || (9683 == GlobalFiModInstNr[1]) || (9683 == GlobalFiModInstNr[2]) || (9683 == GlobalFiModInstNr[3]))));
	Tile mesh_9_25(
		.clock(clock),
		.io_in_a_0(r_313_0),
		.io_in_b_0(b_809_0),
		.io_in_d_0(b_1833_0),
		.io_in_control_0_dataflow(mesh_9_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2857_0),
		.io_in_last_0(r_3881_0),
		.io_in_valid_0(r_1833_0),
		.io_out_a_0(_mesh_9_25_io_out_a_0),
		.io_out_c_0(_mesh_9_25_io_out_c_0),
		.io_out_b_0(_mesh_9_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_25_io_out_id_0),
		.io_out_last_0(_mesh_9_25_io_out_last_0),
		.io_out_valid_0(_mesh_9_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9684 == GlobalFiModInstNr[0]) || (9684 == GlobalFiModInstNr[1]) || (9684 == GlobalFiModInstNr[2]) || (9684 == GlobalFiModInstNr[3]))));
	Tile mesh_9_26(
		.clock(clock),
		.io_in_a_0(r_314_0),
		.io_in_b_0(b_841_0),
		.io_in_d_0(b_1865_0),
		.io_in_control_0_dataflow(mesh_9_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2889_0),
		.io_in_last_0(r_3913_0),
		.io_in_valid_0(r_1865_0),
		.io_out_a_0(_mesh_9_26_io_out_a_0),
		.io_out_c_0(_mesh_9_26_io_out_c_0),
		.io_out_b_0(_mesh_9_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_26_io_out_id_0),
		.io_out_last_0(_mesh_9_26_io_out_last_0),
		.io_out_valid_0(_mesh_9_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9685 == GlobalFiModInstNr[0]) || (9685 == GlobalFiModInstNr[1]) || (9685 == GlobalFiModInstNr[2]) || (9685 == GlobalFiModInstNr[3]))));
	Tile mesh_9_27(
		.clock(clock),
		.io_in_a_0(r_315_0),
		.io_in_b_0(b_873_0),
		.io_in_d_0(b_1897_0),
		.io_in_control_0_dataflow(mesh_9_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2921_0),
		.io_in_last_0(r_3945_0),
		.io_in_valid_0(r_1897_0),
		.io_out_a_0(_mesh_9_27_io_out_a_0),
		.io_out_c_0(_mesh_9_27_io_out_c_0),
		.io_out_b_0(_mesh_9_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_27_io_out_id_0),
		.io_out_last_0(_mesh_9_27_io_out_last_0),
		.io_out_valid_0(_mesh_9_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9686 == GlobalFiModInstNr[0]) || (9686 == GlobalFiModInstNr[1]) || (9686 == GlobalFiModInstNr[2]) || (9686 == GlobalFiModInstNr[3]))));
	Tile mesh_9_28(
		.clock(clock),
		.io_in_a_0(r_316_0),
		.io_in_b_0(b_905_0),
		.io_in_d_0(b_1929_0),
		.io_in_control_0_dataflow(mesh_9_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2953_0),
		.io_in_last_0(r_3977_0),
		.io_in_valid_0(r_1929_0),
		.io_out_a_0(_mesh_9_28_io_out_a_0),
		.io_out_c_0(_mesh_9_28_io_out_c_0),
		.io_out_b_0(_mesh_9_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_28_io_out_id_0),
		.io_out_last_0(_mesh_9_28_io_out_last_0),
		.io_out_valid_0(_mesh_9_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9687 == GlobalFiModInstNr[0]) || (9687 == GlobalFiModInstNr[1]) || (9687 == GlobalFiModInstNr[2]) || (9687 == GlobalFiModInstNr[3]))));
	Tile mesh_9_29(
		.clock(clock),
		.io_in_a_0(r_317_0),
		.io_in_b_0(b_937_0),
		.io_in_d_0(b_1961_0),
		.io_in_control_0_dataflow(mesh_9_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2985_0),
		.io_in_last_0(r_4009_0),
		.io_in_valid_0(r_1961_0),
		.io_out_a_0(_mesh_9_29_io_out_a_0),
		.io_out_c_0(_mesh_9_29_io_out_c_0),
		.io_out_b_0(_mesh_9_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_29_io_out_id_0),
		.io_out_last_0(_mesh_9_29_io_out_last_0),
		.io_out_valid_0(_mesh_9_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9688 == GlobalFiModInstNr[0]) || (9688 == GlobalFiModInstNr[1]) || (9688 == GlobalFiModInstNr[2]) || (9688 == GlobalFiModInstNr[3]))));
	Tile mesh_9_30(
		.clock(clock),
		.io_in_a_0(r_318_0),
		.io_in_b_0(b_969_0),
		.io_in_d_0(b_1993_0),
		.io_in_control_0_dataflow(mesh_9_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3017_0),
		.io_in_last_0(r_4041_0),
		.io_in_valid_0(r_1993_0),
		.io_out_a_0(_mesh_9_30_io_out_a_0),
		.io_out_c_0(_mesh_9_30_io_out_c_0),
		.io_out_b_0(_mesh_9_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_30_io_out_id_0),
		.io_out_last_0(_mesh_9_30_io_out_last_0),
		.io_out_valid_0(_mesh_9_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9689 == GlobalFiModInstNr[0]) || (9689 == GlobalFiModInstNr[1]) || (9689 == GlobalFiModInstNr[2]) || (9689 == GlobalFiModInstNr[3]))));
	Tile mesh_9_31(
		.clock(clock),
		.io_in_a_0(r_319_0),
		.io_in_b_0(b_1001_0),
		.io_in_d_0(b_2025_0),
		.io_in_control_0_dataflow(mesh_9_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_9_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_9_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3049_0),
		.io_in_last_0(r_4073_0),
		.io_in_valid_0(r_2025_0),
		.io_out_a_0(_mesh_9_31_io_out_a_0),
		.io_out_c_0(_mesh_9_31_io_out_c_0),
		.io_out_b_0(_mesh_9_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_9_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_9_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_9_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_9_31_io_out_id_0),
		.io_out_last_0(_mesh_9_31_io_out_last_0),
		.io_out_valid_0(_mesh_9_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9690 == GlobalFiModInstNr[0]) || (9690 == GlobalFiModInstNr[1]) || (9690 == GlobalFiModInstNr[2]) || (9690 == GlobalFiModInstNr[3]))));
	Tile mesh_10_0(
		.clock(clock),
		.io_in_a_0(r_320_0),
		.io_in_b_0(b_10_0),
		.io_in_d_0(b_1034_0),
		.io_in_control_0_dataflow(mesh_10_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2058_0),
		.io_in_last_0(r_3082_0),
		.io_in_valid_0(r_1034_0),
		.io_out_a_0(_mesh_10_0_io_out_a_0),
		.io_out_c_0(_mesh_10_0_io_out_c_0),
		.io_out_b_0(_mesh_10_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_0_io_out_id_0),
		.io_out_last_0(_mesh_10_0_io_out_last_0),
		.io_out_valid_0(_mesh_10_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9691 == GlobalFiModInstNr[0]) || (9691 == GlobalFiModInstNr[1]) || (9691 == GlobalFiModInstNr[2]) || (9691 == GlobalFiModInstNr[3]))));
	Tile mesh_10_1(
		.clock(clock),
		.io_in_a_0(r_321_0),
		.io_in_b_0(b_42_0),
		.io_in_d_0(b_1066_0),
		.io_in_control_0_dataflow(mesh_10_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2090_0),
		.io_in_last_0(r_3114_0),
		.io_in_valid_0(r_1066_0),
		.io_out_a_0(_mesh_10_1_io_out_a_0),
		.io_out_c_0(_mesh_10_1_io_out_c_0),
		.io_out_b_0(_mesh_10_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_1_io_out_id_0),
		.io_out_last_0(_mesh_10_1_io_out_last_0),
		.io_out_valid_0(_mesh_10_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9692 == GlobalFiModInstNr[0]) || (9692 == GlobalFiModInstNr[1]) || (9692 == GlobalFiModInstNr[2]) || (9692 == GlobalFiModInstNr[3]))));
	Tile mesh_10_2(
		.clock(clock),
		.io_in_a_0(r_322_0),
		.io_in_b_0(b_74_0),
		.io_in_d_0(b_1098_0),
		.io_in_control_0_dataflow(mesh_10_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2122_0),
		.io_in_last_0(r_3146_0),
		.io_in_valid_0(r_1098_0),
		.io_out_a_0(_mesh_10_2_io_out_a_0),
		.io_out_c_0(_mesh_10_2_io_out_c_0),
		.io_out_b_0(_mesh_10_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_2_io_out_id_0),
		.io_out_last_0(_mesh_10_2_io_out_last_0),
		.io_out_valid_0(_mesh_10_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9693 == GlobalFiModInstNr[0]) || (9693 == GlobalFiModInstNr[1]) || (9693 == GlobalFiModInstNr[2]) || (9693 == GlobalFiModInstNr[3]))));
	Tile mesh_10_3(
		.clock(clock),
		.io_in_a_0(r_323_0),
		.io_in_b_0(b_106_0),
		.io_in_d_0(b_1130_0),
		.io_in_control_0_dataflow(mesh_10_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2154_0),
		.io_in_last_0(r_3178_0),
		.io_in_valid_0(r_1130_0),
		.io_out_a_0(_mesh_10_3_io_out_a_0),
		.io_out_c_0(_mesh_10_3_io_out_c_0),
		.io_out_b_0(_mesh_10_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_3_io_out_id_0),
		.io_out_last_0(_mesh_10_3_io_out_last_0),
		.io_out_valid_0(_mesh_10_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9694 == GlobalFiModInstNr[0]) || (9694 == GlobalFiModInstNr[1]) || (9694 == GlobalFiModInstNr[2]) || (9694 == GlobalFiModInstNr[3]))));
	Tile mesh_10_4(
		.clock(clock),
		.io_in_a_0(r_324_0),
		.io_in_b_0(b_138_0),
		.io_in_d_0(b_1162_0),
		.io_in_control_0_dataflow(mesh_10_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2186_0),
		.io_in_last_0(r_3210_0),
		.io_in_valid_0(r_1162_0),
		.io_out_a_0(_mesh_10_4_io_out_a_0),
		.io_out_c_0(_mesh_10_4_io_out_c_0),
		.io_out_b_0(_mesh_10_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_4_io_out_id_0),
		.io_out_last_0(_mesh_10_4_io_out_last_0),
		.io_out_valid_0(_mesh_10_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9695 == GlobalFiModInstNr[0]) || (9695 == GlobalFiModInstNr[1]) || (9695 == GlobalFiModInstNr[2]) || (9695 == GlobalFiModInstNr[3]))));
	Tile mesh_10_5(
		.clock(clock),
		.io_in_a_0(r_325_0),
		.io_in_b_0(b_170_0),
		.io_in_d_0(b_1194_0),
		.io_in_control_0_dataflow(mesh_10_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2218_0),
		.io_in_last_0(r_3242_0),
		.io_in_valid_0(r_1194_0),
		.io_out_a_0(_mesh_10_5_io_out_a_0),
		.io_out_c_0(_mesh_10_5_io_out_c_0),
		.io_out_b_0(_mesh_10_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_5_io_out_id_0),
		.io_out_last_0(_mesh_10_5_io_out_last_0),
		.io_out_valid_0(_mesh_10_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9696 == GlobalFiModInstNr[0]) || (9696 == GlobalFiModInstNr[1]) || (9696 == GlobalFiModInstNr[2]) || (9696 == GlobalFiModInstNr[3]))));
	Tile mesh_10_6(
		.clock(clock),
		.io_in_a_0(r_326_0),
		.io_in_b_0(b_202_0),
		.io_in_d_0(b_1226_0),
		.io_in_control_0_dataflow(mesh_10_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2250_0),
		.io_in_last_0(r_3274_0),
		.io_in_valid_0(r_1226_0),
		.io_out_a_0(_mesh_10_6_io_out_a_0),
		.io_out_c_0(_mesh_10_6_io_out_c_0),
		.io_out_b_0(_mesh_10_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_6_io_out_id_0),
		.io_out_last_0(_mesh_10_6_io_out_last_0),
		.io_out_valid_0(_mesh_10_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9697 == GlobalFiModInstNr[0]) || (9697 == GlobalFiModInstNr[1]) || (9697 == GlobalFiModInstNr[2]) || (9697 == GlobalFiModInstNr[3]))));
	Tile mesh_10_7(
		.clock(clock),
		.io_in_a_0(r_327_0),
		.io_in_b_0(b_234_0),
		.io_in_d_0(b_1258_0),
		.io_in_control_0_dataflow(mesh_10_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2282_0),
		.io_in_last_0(r_3306_0),
		.io_in_valid_0(r_1258_0),
		.io_out_a_0(_mesh_10_7_io_out_a_0),
		.io_out_c_0(_mesh_10_7_io_out_c_0),
		.io_out_b_0(_mesh_10_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_7_io_out_id_0),
		.io_out_last_0(_mesh_10_7_io_out_last_0),
		.io_out_valid_0(_mesh_10_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9698 == GlobalFiModInstNr[0]) || (9698 == GlobalFiModInstNr[1]) || (9698 == GlobalFiModInstNr[2]) || (9698 == GlobalFiModInstNr[3]))));
	Tile mesh_10_8(
		.clock(clock),
		.io_in_a_0(r_328_0),
		.io_in_b_0(b_266_0),
		.io_in_d_0(b_1290_0),
		.io_in_control_0_dataflow(mesh_10_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2314_0),
		.io_in_last_0(r_3338_0),
		.io_in_valid_0(r_1290_0),
		.io_out_a_0(_mesh_10_8_io_out_a_0),
		.io_out_c_0(_mesh_10_8_io_out_c_0),
		.io_out_b_0(_mesh_10_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_8_io_out_id_0),
		.io_out_last_0(_mesh_10_8_io_out_last_0),
		.io_out_valid_0(_mesh_10_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9699 == GlobalFiModInstNr[0]) || (9699 == GlobalFiModInstNr[1]) || (9699 == GlobalFiModInstNr[2]) || (9699 == GlobalFiModInstNr[3]))));
	Tile mesh_10_9(
		.clock(clock),
		.io_in_a_0(r_329_0),
		.io_in_b_0(b_298_0),
		.io_in_d_0(b_1322_0),
		.io_in_control_0_dataflow(mesh_10_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2346_0),
		.io_in_last_0(r_3370_0),
		.io_in_valid_0(r_1322_0),
		.io_out_a_0(_mesh_10_9_io_out_a_0),
		.io_out_c_0(_mesh_10_9_io_out_c_0),
		.io_out_b_0(_mesh_10_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_9_io_out_id_0),
		.io_out_last_0(_mesh_10_9_io_out_last_0),
		.io_out_valid_0(_mesh_10_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9700 == GlobalFiModInstNr[0]) || (9700 == GlobalFiModInstNr[1]) || (9700 == GlobalFiModInstNr[2]) || (9700 == GlobalFiModInstNr[3]))));
	Tile mesh_10_10(
		.clock(clock),
		.io_in_a_0(r_330_0),
		.io_in_b_0(b_330_0),
		.io_in_d_0(b_1354_0),
		.io_in_control_0_dataflow(mesh_10_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2378_0),
		.io_in_last_0(r_3402_0),
		.io_in_valid_0(r_1354_0),
		.io_out_a_0(_mesh_10_10_io_out_a_0),
		.io_out_c_0(_mesh_10_10_io_out_c_0),
		.io_out_b_0(_mesh_10_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_10_io_out_id_0),
		.io_out_last_0(_mesh_10_10_io_out_last_0),
		.io_out_valid_0(_mesh_10_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9701 == GlobalFiModInstNr[0]) || (9701 == GlobalFiModInstNr[1]) || (9701 == GlobalFiModInstNr[2]) || (9701 == GlobalFiModInstNr[3]))));
	Tile mesh_10_11(
		.clock(clock),
		.io_in_a_0(r_331_0),
		.io_in_b_0(b_362_0),
		.io_in_d_0(b_1386_0),
		.io_in_control_0_dataflow(mesh_10_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2410_0),
		.io_in_last_0(r_3434_0),
		.io_in_valid_0(r_1386_0),
		.io_out_a_0(_mesh_10_11_io_out_a_0),
		.io_out_c_0(_mesh_10_11_io_out_c_0),
		.io_out_b_0(_mesh_10_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_11_io_out_id_0),
		.io_out_last_0(_mesh_10_11_io_out_last_0),
		.io_out_valid_0(_mesh_10_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9702 == GlobalFiModInstNr[0]) || (9702 == GlobalFiModInstNr[1]) || (9702 == GlobalFiModInstNr[2]) || (9702 == GlobalFiModInstNr[3]))));
	Tile mesh_10_12(
		.clock(clock),
		.io_in_a_0(r_332_0),
		.io_in_b_0(b_394_0),
		.io_in_d_0(b_1418_0),
		.io_in_control_0_dataflow(mesh_10_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2442_0),
		.io_in_last_0(r_3466_0),
		.io_in_valid_0(r_1418_0),
		.io_out_a_0(_mesh_10_12_io_out_a_0),
		.io_out_c_0(_mesh_10_12_io_out_c_0),
		.io_out_b_0(_mesh_10_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_12_io_out_id_0),
		.io_out_last_0(_mesh_10_12_io_out_last_0),
		.io_out_valid_0(_mesh_10_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9703 == GlobalFiModInstNr[0]) || (9703 == GlobalFiModInstNr[1]) || (9703 == GlobalFiModInstNr[2]) || (9703 == GlobalFiModInstNr[3]))));
	Tile mesh_10_13(
		.clock(clock),
		.io_in_a_0(r_333_0),
		.io_in_b_0(b_426_0),
		.io_in_d_0(b_1450_0),
		.io_in_control_0_dataflow(mesh_10_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2474_0),
		.io_in_last_0(r_3498_0),
		.io_in_valid_0(r_1450_0),
		.io_out_a_0(_mesh_10_13_io_out_a_0),
		.io_out_c_0(_mesh_10_13_io_out_c_0),
		.io_out_b_0(_mesh_10_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_13_io_out_id_0),
		.io_out_last_0(_mesh_10_13_io_out_last_0),
		.io_out_valid_0(_mesh_10_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9704 == GlobalFiModInstNr[0]) || (9704 == GlobalFiModInstNr[1]) || (9704 == GlobalFiModInstNr[2]) || (9704 == GlobalFiModInstNr[3]))));
	Tile mesh_10_14(
		.clock(clock),
		.io_in_a_0(r_334_0),
		.io_in_b_0(b_458_0),
		.io_in_d_0(b_1482_0),
		.io_in_control_0_dataflow(mesh_10_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2506_0),
		.io_in_last_0(r_3530_0),
		.io_in_valid_0(r_1482_0),
		.io_out_a_0(_mesh_10_14_io_out_a_0),
		.io_out_c_0(_mesh_10_14_io_out_c_0),
		.io_out_b_0(_mesh_10_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_14_io_out_id_0),
		.io_out_last_0(_mesh_10_14_io_out_last_0),
		.io_out_valid_0(_mesh_10_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9705 == GlobalFiModInstNr[0]) || (9705 == GlobalFiModInstNr[1]) || (9705 == GlobalFiModInstNr[2]) || (9705 == GlobalFiModInstNr[3]))));
	Tile mesh_10_15(
		.clock(clock),
		.io_in_a_0(r_335_0),
		.io_in_b_0(b_490_0),
		.io_in_d_0(b_1514_0),
		.io_in_control_0_dataflow(mesh_10_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2538_0),
		.io_in_last_0(r_3562_0),
		.io_in_valid_0(r_1514_0),
		.io_out_a_0(_mesh_10_15_io_out_a_0),
		.io_out_c_0(_mesh_10_15_io_out_c_0),
		.io_out_b_0(_mesh_10_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_15_io_out_id_0),
		.io_out_last_0(_mesh_10_15_io_out_last_0),
		.io_out_valid_0(_mesh_10_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9706 == GlobalFiModInstNr[0]) || (9706 == GlobalFiModInstNr[1]) || (9706 == GlobalFiModInstNr[2]) || (9706 == GlobalFiModInstNr[3]))));
	Tile mesh_10_16(
		.clock(clock),
		.io_in_a_0(r_336_0),
		.io_in_b_0(b_522_0),
		.io_in_d_0(b_1546_0),
		.io_in_control_0_dataflow(mesh_10_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2570_0),
		.io_in_last_0(r_3594_0),
		.io_in_valid_0(r_1546_0),
		.io_out_a_0(_mesh_10_16_io_out_a_0),
		.io_out_c_0(_mesh_10_16_io_out_c_0),
		.io_out_b_0(_mesh_10_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_16_io_out_id_0),
		.io_out_last_0(_mesh_10_16_io_out_last_0),
		.io_out_valid_0(_mesh_10_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9707 == GlobalFiModInstNr[0]) || (9707 == GlobalFiModInstNr[1]) || (9707 == GlobalFiModInstNr[2]) || (9707 == GlobalFiModInstNr[3]))));
	Tile mesh_10_17(
		.clock(clock),
		.io_in_a_0(r_337_0),
		.io_in_b_0(b_554_0),
		.io_in_d_0(b_1578_0),
		.io_in_control_0_dataflow(mesh_10_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2602_0),
		.io_in_last_0(r_3626_0),
		.io_in_valid_0(r_1578_0),
		.io_out_a_0(_mesh_10_17_io_out_a_0),
		.io_out_c_0(_mesh_10_17_io_out_c_0),
		.io_out_b_0(_mesh_10_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_17_io_out_id_0),
		.io_out_last_0(_mesh_10_17_io_out_last_0),
		.io_out_valid_0(_mesh_10_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9708 == GlobalFiModInstNr[0]) || (9708 == GlobalFiModInstNr[1]) || (9708 == GlobalFiModInstNr[2]) || (9708 == GlobalFiModInstNr[3]))));
	Tile mesh_10_18(
		.clock(clock),
		.io_in_a_0(r_338_0),
		.io_in_b_0(b_586_0),
		.io_in_d_0(b_1610_0),
		.io_in_control_0_dataflow(mesh_10_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2634_0),
		.io_in_last_0(r_3658_0),
		.io_in_valid_0(r_1610_0),
		.io_out_a_0(_mesh_10_18_io_out_a_0),
		.io_out_c_0(_mesh_10_18_io_out_c_0),
		.io_out_b_0(_mesh_10_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_18_io_out_id_0),
		.io_out_last_0(_mesh_10_18_io_out_last_0),
		.io_out_valid_0(_mesh_10_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9709 == GlobalFiModInstNr[0]) || (9709 == GlobalFiModInstNr[1]) || (9709 == GlobalFiModInstNr[2]) || (9709 == GlobalFiModInstNr[3]))));
	Tile mesh_10_19(
		.clock(clock),
		.io_in_a_0(r_339_0),
		.io_in_b_0(b_618_0),
		.io_in_d_0(b_1642_0),
		.io_in_control_0_dataflow(mesh_10_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2666_0),
		.io_in_last_0(r_3690_0),
		.io_in_valid_0(r_1642_0),
		.io_out_a_0(_mesh_10_19_io_out_a_0),
		.io_out_c_0(_mesh_10_19_io_out_c_0),
		.io_out_b_0(_mesh_10_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_19_io_out_id_0),
		.io_out_last_0(_mesh_10_19_io_out_last_0),
		.io_out_valid_0(_mesh_10_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9710 == GlobalFiModInstNr[0]) || (9710 == GlobalFiModInstNr[1]) || (9710 == GlobalFiModInstNr[2]) || (9710 == GlobalFiModInstNr[3]))));
	Tile mesh_10_20(
		.clock(clock),
		.io_in_a_0(r_340_0),
		.io_in_b_0(b_650_0),
		.io_in_d_0(b_1674_0),
		.io_in_control_0_dataflow(mesh_10_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2698_0),
		.io_in_last_0(r_3722_0),
		.io_in_valid_0(r_1674_0),
		.io_out_a_0(_mesh_10_20_io_out_a_0),
		.io_out_c_0(_mesh_10_20_io_out_c_0),
		.io_out_b_0(_mesh_10_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_20_io_out_id_0),
		.io_out_last_0(_mesh_10_20_io_out_last_0),
		.io_out_valid_0(_mesh_10_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9711 == GlobalFiModInstNr[0]) || (9711 == GlobalFiModInstNr[1]) || (9711 == GlobalFiModInstNr[2]) || (9711 == GlobalFiModInstNr[3]))));
	Tile mesh_10_21(
		.clock(clock),
		.io_in_a_0(r_341_0),
		.io_in_b_0(b_682_0),
		.io_in_d_0(b_1706_0),
		.io_in_control_0_dataflow(mesh_10_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2730_0),
		.io_in_last_0(r_3754_0),
		.io_in_valid_0(r_1706_0),
		.io_out_a_0(_mesh_10_21_io_out_a_0),
		.io_out_c_0(_mesh_10_21_io_out_c_0),
		.io_out_b_0(_mesh_10_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_21_io_out_id_0),
		.io_out_last_0(_mesh_10_21_io_out_last_0),
		.io_out_valid_0(_mesh_10_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9712 == GlobalFiModInstNr[0]) || (9712 == GlobalFiModInstNr[1]) || (9712 == GlobalFiModInstNr[2]) || (9712 == GlobalFiModInstNr[3]))));
	Tile mesh_10_22(
		.clock(clock),
		.io_in_a_0(r_342_0),
		.io_in_b_0(b_714_0),
		.io_in_d_0(b_1738_0),
		.io_in_control_0_dataflow(mesh_10_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2762_0),
		.io_in_last_0(r_3786_0),
		.io_in_valid_0(r_1738_0),
		.io_out_a_0(_mesh_10_22_io_out_a_0),
		.io_out_c_0(_mesh_10_22_io_out_c_0),
		.io_out_b_0(_mesh_10_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_22_io_out_id_0),
		.io_out_last_0(_mesh_10_22_io_out_last_0),
		.io_out_valid_0(_mesh_10_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9713 == GlobalFiModInstNr[0]) || (9713 == GlobalFiModInstNr[1]) || (9713 == GlobalFiModInstNr[2]) || (9713 == GlobalFiModInstNr[3]))));
	Tile mesh_10_23(
		.clock(clock),
		.io_in_a_0(r_343_0),
		.io_in_b_0(b_746_0),
		.io_in_d_0(b_1770_0),
		.io_in_control_0_dataflow(mesh_10_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2794_0),
		.io_in_last_0(r_3818_0),
		.io_in_valid_0(r_1770_0),
		.io_out_a_0(_mesh_10_23_io_out_a_0),
		.io_out_c_0(_mesh_10_23_io_out_c_0),
		.io_out_b_0(_mesh_10_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_23_io_out_id_0),
		.io_out_last_0(_mesh_10_23_io_out_last_0),
		.io_out_valid_0(_mesh_10_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9714 == GlobalFiModInstNr[0]) || (9714 == GlobalFiModInstNr[1]) || (9714 == GlobalFiModInstNr[2]) || (9714 == GlobalFiModInstNr[3]))));
	Tile mesh_10_24(
		.clock(clock),
		.io_in_a_0(r_344_0),
		.io_in_b_0(b_778_0),
		.io_in_d_0(b_1802_0),
		.io_in_control_0_dataflow(mesh_10_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2826_0),
		.io_in_last_0(r_3850_0),
		.io_in_valid_0(r_1802_0),
		.io_out_a_0(_mesh_10_24_io_out_a_0),
		.io_out_c_0(_mesh_10_24_io_out_c_0),
		.io_out_b_0(_mesh_10_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_24_io_out_id_0),
		.io_out_last_0(_mesh_10_24_io_out_last_0),
		.io_out_valid_0(_mesh_10_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9715 == GlobalFiModInstNr[0]) || (9715 == GlobalFiModInstNr[1]) || (9715 == GlobalFiModInstNr[2]) || (9715 == GlobalFiModInstNr[3]))));
	Tile mesh_10_25(
		.clock(clock),
		.io_in_a_0(r_345_0),
		.io_in_b_0(b_810_0),
		.io_in_d_0(b_1834_0),
		.io_in_control_0_dataflow(mesh_10_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2858_0),
		.io_in_last_0(r_3882_0),
		.io_in_valid_0(r_1834_0),
		.io_out_a_0(_mesh_10_25_io_out_a_0),
		.io_out_c_0(_mesh_10_25_io_out_c_0),
		.io_out_b_0(_mesh_10_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_25_io_out_id_0),
		.io_out_last_0(_mesh_10_25_io_out_last_0),
		.io_out_valid_0(_mesh_10_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9716 == GlobalFiModInstNr[0]) || (9716 == GlobalFiModInstNr[1]) || (9716 == GlobalFiModInstNr[2]) || (9716 == GlobalFiModInstNr[3]))));
	Tile mesh_10_26(
		.clock(clock),
		.io_in_a_0(r_346_0),
		.io_in_b_0(b_842_0),
		.io_in_d_0(b_1866_0),
		.io_in_control_0_dataflow(mesh_10_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2890_0),
		.io_in_last_0(r_3914_0),
		.io_in_valid_0(r_1866_0),
		.io_out_a_0(_mesh_10_26_io_out_a_0),
		.io_out_c_0(_mesh_10_26_io_out_c_0),
		.io_out_b_0(_mesh_10_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_26_io_out_id_0),
		.io_out_last_0(_mesh_10_26_io_out_last_0),
		.io_out_valid_0(_mesh_10_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9717 == GlobalFiModInstNr[0]) || (9717 == GlobalFiModInstNr[1]) || (9717 == GlobalFiModInstNr[2]) || (9717 == GlobalFiModInstNr[3]))));
	Tile mesh_10_27(
		.clock(clock),
		.io_in_a_0(r_347_0),
		.io_in_b_0(b_874_0),
		.io_in_d_0(b_1898_0),
		.io_in_control_0_dataflow(mesh_10_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2922_0),
		.io_in_last_0(r_3946_0),
		.io_in_valid_0(r_1898_0),
		.io_out_a_0(_mesh_10_27_io_out_a_0),
		.io_out_c_0(_mesh_10_27_io_out_c_0),
		.io_out_b_0(_mesh_10_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_27_io_out_id_0),
		.io_out_last_0(_mesh_10_27_io_out_last_0),
		.io_out_valid_0(_mesh_10_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9718 == GlobalFiModInstNr[0]) || (9718 == GlobalFiModInstNr[1]) || (9718 == GlobalFiModInstNr[2]) || (9718 == GlobalFiModInstNr[3]))));
	Tile mesh_10_28(
		.clock(clock),
		.io_in_a_0(r_348_0),
		.io_in_b_0(b_906_0),
		.io_in_d_0(b_1930_0),
		.io_in_control_0_dataflow(mesh_10_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2954_0),
		.io_in_last_0(r_3978_0),
		.io_in_valid_0(r_1930_0),
		.io_out_a_0(_mesh_10_28_io_out_a_0),
		.io_out_c_0(_mesh_10_28_io_out_c_0),
		.io_out_b_0(_mesh_10_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_28_io_out_id_0),
		.io_out_last_0(_mesh_10_28_io_out_last_0),
		.io_out_valid_0(_mesh_10_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9719 == GlobalFiModInstNr[0]) || (9719 == GlobalFiModInstNr[1]) || (9719 == GlobalFiModInstNr[2]) || (9719 == GlobalFiModInstNr[3]))));
	Tile mesh_10_29(
		.clock(clock),
		.io_in_a_0(r_349_0),
		.io_in_b_0(b_938_0),
		.io_in_d_0(b_1962_0),
		.io_in_control_0_dataflow(mesh_10_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2986_0),
		.io_in_last_0(r_4010_0),
		.io_in_valid_0(r_1962_0),
		.io_out_a_0(_mesh_10_29_io_out_a_0),
		.io_out_c_0(_mesh_10_29_io_out_c_0),
		.io_out_b_0(_mesh_10_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_29_io_out_id_0),
		.io_out_last_0(_mesh_10_29_io_out_last_0),
		.io_out_valid_0(_mesh_10_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9720 == GlobalFiModInstNr[0]) || (9720 == GlobalFiModInstNr[1]) || (9720 == GlobalFiModInstNr[2]) || (9720 == GlobalFiModInstNr[3]))));
	Tile mesh_10_30(
		.clock(clock),
		.io_in_a_0(r_350_0),
		.io_in_b_0(b_970_0),
		.io_in_d_0(b_1994_0),
		.io_in_control_0_dataflow(mesh_10_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3018_0),
		.io_in_last_0(r_4042_0),
		.io_in_valid_0(r_1994_0),
		.io_out_a_0(_mesh_10_30_io_out_a_0),
		.io_out_c_0(_mesh_10_30_io_out_c_0),
		.io_out_b_0(_mesh_10_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_30_io_out_id_0),
		.io_out_last_0(_mesh_10_30_io_out_last_0),
		.io_out_valid_0(_mesh_10_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9721 == GlobalFiModInstNr[0]) || (9721 == GlobalFiModInstNr[1]) || (9721 == GlobalFiModInstNr[2]) || (9721 == GlobalFiModInstNr[3]))));
	Tile mesh_10_31(
		.clock(clock),
		.io_in_a_0(r_351_0),
		.io_in_b_0(b_1002_0),
		.io_in_d_0(b_2026_0),
		.io_in_control_0_dataflow(mesh_10_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_10_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_10_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3050_0),
		.io_in_last_0(r_4074_0),
		.io_in_valid_0(r_2026_0),
		.io_out_a_0(_mesh_10_31_io_out_a_0),
		.io_out_c_0(_mesh_10_31_io_out_c_0),
		.io_out_b_0(_mesh_10_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_10_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_10_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_10_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_10_31_io_out_id_0),
		.io_out_last_0(_mesh_10_31_io_out_last_0),
		.io_out_valid_0(_mesh_10_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9722 == GlobalFiModInstNr[0]) || (9722 == GlobalFiModInstNr[1]) || (9722 == GlobalFiModInstNr[2]) || (9722 == GlobalFiModInstNr[3]))));
	Tile mesh_11_0(
		.clock(clock),
		.io_in_a_0(r_352_0),
		.io_in_b_0(b_11_0),
		.io_in_d_0(b_1035_0),
		.io_in_control_0_dataflow(mesh_11_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2059_0),
		.io_in_last_0(r_3083_0),
		.io_in_valid_0(r_1035_0),
		.io_out_a_0(_mesh_11_0_io_out_a_0),
		.io_out_c_0(_mesh_11_0_io_out_c_0),
		.io_out_b_0(_mesh_11_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_0_io_out_id_0),
		.io_out_last_0(_mesh_11_0_io_out_last_0),
		.io_out_valid_0(_mesh_11_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9723 == GlobalFiModInstNr[0]) || (9723 == GlobalFiModInstNr[1]) || (9723 == GlobalFiModInstNr[2]) || (9723 == GlobalFiModInstNr[3]))));
	Tile mesh_11_1(
		.clock(clock),
		.io_in_a_0(r_353_0),
		.io_in_b_0(b_43_0),
		.io_in_d_0(b_1067_0),
		.io_in_control_0_dataflow(mesh_11_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2091_0),
		.io_in_last_0(r_3115_0),
		.io_in_valid_0(r_1067_0),
		.io_out_a_0(_mesh_11_1_io_out_a_0),
		.io_out_c_0(_mesh_11_1_io_out_c_0),
		.io_out_b_0(_mesh_11_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_1_io_out_id_0),
		.io_out_last_0(_mesh_11_1_io_out_last_0),
		.io_out_valid_0(_mesh_11_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9724 == GlobalFiModInstNr[0]) || (9724 == GlobalFiModInstNr[1]) || (9724 == GlobalFiModInstNr[2]) || (9724 == GlobalFiModInstNr[3]))));
	Tile mesh_11_2(
		.clock(clock),
		.io_in_a_0(r_354_0),
		.io_in_b_0(b_75_0),
		.io_in_d_0(b_1099_0),
		.io_in_control_0_dataflow(mesh_11_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2123_0),
		.io_in_last_0(r_3147_0),
		.io_in_valid_0(r_1099_0),
		.io_out_a_0(_mesh_11_2_io_out_a_0),
		.io_out_c_0(_mesh_11_2_io_out_c_0),
		.io_out_b_0(_mesh_11_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_2_io_out_id_0),
		.io_out_last_0(_mesh_11_2_io_out_last_0),
		.io_out_valid_0(_mesh_11_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9725 == GlobalFiModInstNr[0]) || (9725 == GlobalFiModInstNr[1]) || (9725 == GlobalFiModInstNr[2]) || (9725 == GlobalFiModInstNr[3]))));
	Tile mesh_11_3(
		.clock(clock),
		.io_in_a_0(r_355_0),
		.io_in_b_0(b_107_0),
		.io_in_d_0(b_1131_0),
		.io_in_control_0_dataflow(mesh_11_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2155_0),
		.io_in_last_0(r_3179_0),
		.io_in_valid_0(r_1131_0),
		.io_out_a_0(_mesh_11_3_io_out_a_0),
		.io_out_c_0(_mesh_11_3_io_out_c_0),
		.io_out_b_0(_mesh_11_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_3_io_out_id_0),
		.io_out_last_0(_mesh_11_3_io_out_last_0),
		.io_out_valid_0(_mesh_11_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9726 == GlobalFiModInstNr[0]) || (9726 == GlobalFiModInstNr[1]) || (9726 == GlobalFiModInstNr[2]) || (9726 == GlobalFiModInstNr[3]))));
	Tile mesh_11_4(
		.clock(clock),
		.io_in_a_0(r_356_0),
		.io_in_b_0(b_139_0),
		.io_in_d_0(b_1163_0),
		.io_in_control_0_dataflow(mesh_11_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2187_0),
		.io_in_last_0(r_3211_0),
		.io_in_valid_0(r_1163_0),
		.io_out_a_0(_mesh_11_4_io_out_a_0),
		.io_out_c_0(_mesh_11_4_io_out_c_0),
		.io_out_b_0(_mesh_11_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_4_io_out_id_0),
		.io_out_last_0(_mesh_11_4_io_out_last_0),
		.io_out_valid_0(_mesh_11_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9727 == GlobalFiModInstNr[0]) || (9727 == GlobalFiModInstNr[1]) || (9727 == GlobalFiModInstNr[2]) || (9727 == GlobalFiModInstNr[3]))));
	Tile mesh_11_5(
		.clock(clock),
		.io_in_a_0(r_357_0),
		.io_in_b_0(b_171_0),
		.io_in_d_0(b_1195_0),
		.io_in_control_0_dataflow(mesh_11_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2219_0),
		.io_in_last_0(r_3243_0),
		.io_in_valid_0(r_1195_0),
		.io_out_a_0(_mesh_11_5_io_out_a_0),
		.io_out_c_0(_mesh_11_5_io_out_c_0),
		.io_out_b_0(_mesh_11_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_5_io_out_id_0),
		.io_out_last_0(_mesh_11_5_io_out_last_0),
		.io_out_valid_0(_mesh_11_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9728 == GlobalFiModInstNr[0]) || (9728 == GlobalFiModInstNr[1]) || (9728 == GlobalFiModInstNr[2]) || (9728 == GlobalFiModInstNr[3]))));
	Tile mesh_11_6(
		.clock(clock),
		.io_in_a_0(r_358_0),
		.io_in_b_0(b_203_0),
		.io_in_d_0(b_1227_0),
		.io_in_control_0_dataflow(mesh_11_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2251_0),
		.io_in_last_0(r_3275_0),
		.io_in_valid_0(r_1227_0),
		.io_out_a_0(_mesh_11_6_io_out_a_0),
		.io_out_c_0(_mesh_11_6_io_out_c_0),
		.io_out_b_0(_mesh_11_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_6_io_out_id_0),
		.io_out_last_0(_mesh_11_6_io_out_last_0),
		.io_out_valid_0(_mesh_11_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9729 == GlobalFiModInstNr[0]) || (9729 == GlobalFiModInstNr[1]) || (9729 == GlobalFiModInstNr[2]) || (9729 == GlobalFiModInstNr[3]))));
	Tile mesh_11_7(
		.clock(clock),
		.io_in_a_0(r_359_0),
		.io_in_b_0(b_235_0),
		.io_in_d_0(b_1259_0),
		.io_in_control_0_dataflow(mesh_11_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2283_0),
		.io_in_last_0(r_3307_0),
		.io_in_valid_0(r_1259_0),
		.io_out_a_0(_mesh_11_7_io_out_a_0),
		.io_out_c_0(_mesh_11_7_io_out_c_0),
		.io_out_b_0(_mesh_11_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_7_io_out_id_0),
		.io_out_last_0(_mesh_11_7_io_out_last_0),
		.io_out_valid_0(_mesh_11_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9730 == GlobalFiModInstNr[0]) || (9730 == GlobalFiModInstNr[1]) || (9730 == GlobalFiModInstNr[2]) || (9730 == GlobalFiModInstNr[3]))));
	Tile mesh_11_8(
		.clock(clock),
		.io_in_a_0(r_360_0),
		.io_in_b_0(b_267_0),
		.io_in_d_0(b_1291_0),
		.io_in_control_0_dataflow(mesh_11_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2315_0),
		.io_in_last_0(r_3339_0),
		.io_in_valid_0(r_1291_0),
		.io_out_a_0(_mesh_11_8_io_out_a_0),
		.io_out_c_0(_mesh_11_8_io_out_c_0),
		.io_out_b_0(_mesh_11_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_8_io_out_id_0),
		.io_out_last_0(_mesh_11_8_io_out_last_0),
		.io_out_valid_0(_mesh_11_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9731 == GlobalFiModInstNr[0]) || (9731 == GlobalFiModInstNr[1]) || (9731 == GlobalFiModInstNr[2]) || (9731 == GlobalFiModInstNr[3]))));
	Tile mesh_11_9(
		.clock(clock),
		.io_in_a_0(r_361_0),
		.io_in_b_0(b_299_0),
		.io_in_d_0(b_1323_0),
		.io_in_control_0_dataflow(mesh_11_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2347_0),
		.io_in_last_0(r_3371_0),
		.io_in_valid_0(r_1323_0),
		.io_out_a_0(_mesh_11_9_io_out_a_0),
		.io_out_c_0(_mesh_11_9_io_out_c_0),
		.io_out_b_0(_mesh_11_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_9_io_out_id_0),
		.io_out_last_0(_mesh_11_9_io_out_last_0),
		.io_out_valid_0(_mesh_11_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9732 == GlobalFiModInstNr[0]) || (9732 == GlobalFiModInstNr[1]) || (9732 == GlobalFiModInstNr[2]) || (9732 == GlobalFiModInstNr[3]))));
	Tile mesh_11_10(
		.clock(clock),
		.io_in_a_0(r_362_0),
		.io_in_b_0(b_331_0),
		.io_in_d_0(b_1355_0),
		.io_in_control_0_dataflow(mesh_11_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2379_0),
		.io_in_last_0(r_3403_0),
		.io_in_valid_0(r_1355_0),
		.io_out_a_0(_mesh_11_10_io_out_a_0),
		.io_out_c_0(_mesh_11_10_io_out_c_0),
		.io_out_b_0(_mesh_11_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_10_io_out_id_0),
		.io_out_last_0(_mesh_11_10_io_out_last_0),
		.io_out_valid_0(_mesh_11_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9733 == GlobalFiModInstNr[0]) || (9733 == GlobalFiModInstNr[1]) || (9733 == GlobalFiModInstNr[2]) || (9733 == GlobalFiModInstNr[3]))));
	Tile mesh_11_11(
		.clock(clock),
		.io_in_a_0(r_363_0),
		.io_in_b_0(b_363_0),
		.io_in_d_0(b_1387_0),
		.io_in_control_0_dataflow(mesh_11_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2411_0),
		.io_in_last_0(r_3435_0),
		.io_in_valid_0(r_1387_0),
		.io_out_a_0(_mesh_11_11_io_out_a_0),
		.io_out_c_0(_mesh_11_11_io_out_c_0),
		.io_out_b_0(_mesh_11_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_11_io_out_id_0),
		.io_out_last_0(_mesh_11_11_io_out_last_0),
		.io_out_valid_0(_mesh_11_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9734 == GlobalFiModInstNr[0]) || (9734 == GlobalFiModInstNr[1]) || (9734 == GlobalFiModInstNr[2]) || (9734 == GlobalFiModInstNr[3]))));
	Tile mesh_11_12(
		.clock(clock),
		.io_in_a_0(r_364_0),
		.io_in_b_0(b_395_0),
		.io_in_d_0(b_1419_0),
		.io_in_control_0_dataflow(mesh_11_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2443_0),
		.io_in_last_0(r_3467_0),
		.io_in_valid_0(r_1419_0),
		.io_out_a_0(_mesh_11_12_io_out_a_0),
		.io_out_c_0(_mesh_11_12_io_out_c_0),
		.io_out_b_0(_mesh_11_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_12_io_out_id_0),
		.io_out_last_0(_mesh_11_12_io_out_last_0),
		.io_out_valid_0(_mesh_11_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9735 == GlobalFiModInstNr[0]) || (9735 == GlobalFiModInstNr[1]) || (9735 == GlobalFiModInstNr[2]) || (9735 == GlobalFiModInstNr[3]))));
	Tile mesh_11_13(
		.clock(clock),
		.io_in_a_0(r_365_0),
		.io_in_b_0(b_427_0),
		.io_in_d_0(b_1451_0),
		.io_in_control_0_dataflow(mesh_11_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2475_0),
		.io_in_last_0(r_3499_0),
		.io_in_valid_0(r_1451_0),
		.io_out_a_0(_mesh_11_13_io_out_a_0),
		.io_out_c_0(_mesh_11_13_io_out_c_0),
		.io_out_b_0(_mesh_11_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_13_io_out_id_0),
		.io_out_last_0(_mesh_11_13_io_out_last_0),
		.io_out_valid_0(_mesh_11_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9736 == GlobalFiModInstNr[0]) || (9736 == GlobalFiModInstNr[1]) || (9736 == GlobalFiModInstNr[2]) || (9736 == GlobalFiModInstNr[3]))));
	Tile mesh_11_14(
		.clock(clock),
		.io_in_a_0(r_366_0),
		.io_in_b_0(b_459_0),
		.io_in_d_0(b_1483_0),
		.io_in_control_0_dataflow(mesh_11_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2507_0),
		.io_in_last_0(r_3531_0),
		.io_in_valid_0(r_1483_0),
		.io_out_a_0(_mesh_11_14_io_out_a_0),
		.io_out_c_0(_mesh_11_14_io_out_c_0),
		.io_out_b_0(_mesh_11_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_14_io_out_id_0),
		.io_out_last_0(_mesh_11_14_io_out_last_0),
		.io_out_valid_0(_mesh_11_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9737 == GlobalFiModInstNr[0]) || (9737 == GlobalFiModInstNr[1]) || (9737 == GlobalFiModInstNr[2]) || (9737 == GlobalFiModInstNr[3]))));
	Tile mesh_11_15(
		.clock(clock),
		.io_in_a_0(r_367_0),
		.io_in_b_0(b_491_0),
		.io_in_d_0(b_1515_0),
		.io_in_control_0_dataflow(mesh_11_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2539_0),
		.io_in_last_0(r_3563_0),
		.io_in_valid_0(r_1515_0),
		.io_out_a_0(_mesh_11_15_io_out_a_0),
		.io_out_c_0(_mesh_11_15_io_out_c_0),
		.io_out_b_0(_mesh_11_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_15_io_out_id_0),
		.io_out_last_0(_mesh_11_15_io_out_last_0),
		.io_out_valid_0(_mesh_11_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9738 == GlobalFiModInstNr[0]) || (9738 == GlobalFiModInstNr[1]) || (9738 == GlobalFiModInstNr[2]) || (9738 == GlobalFiModInstNr[3]))));
	Tile mesh_11_16(
		.clock(clock),
		.io_in_a_0(r_368_0),
		.io_in_b_0(b_523_0),
		.io_in_d_0(b_1547_0),
		.io_in_control_0_dataflow(mesh_11_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2571_0),
		.io_in_last_0(r_3595_0),
		.io_in_valid_0(r_1547_0),
		.io_out_a_0(_mesh_11_16_io_out_a_0),
		.io_out_c_0(_mesh_11_16_io_out_c_0),
		.io_out_b_0(_mesh_11_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_16_io_out_id_0),
		.io_out_last_0(_mesh_11_16_io_out_last_0),
		.io_out_valid_0(_mesh_11_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9739 == GlobalFiModInstNr[0]) || (9739 == GlobalFiModInstNr[1]) || (9739 == GlobalFiModInstNr[2]) || (9739 == GlobalFiModInstNr[3]))));
	Tile mesh_11_17(
		.clock(clock),
		.io_in_a_0(r_369_0),
		.io_in_b_0(b_555_0),
		.io_in_d_0(b_1579_0),
		.io_in_control_0_dataflow(mesh_11_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2603_0),
		.io_in_last_0(r_3627_0),
		.io_in_valid_0(r_1579_0),
		.io_out_a_0(_mesh_11_17_io_out_a_0),
		.io_out_c_0(_mesh_11_17_io_out_c_0),
		.io_out_b_0(_mesh_11_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_17_io_out_id_0),
		.io_out_last_0(_mesh_11_17_io_out_last_0),
		.io_out_valid_0(_mesh_11_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9740 == GlobalFiModInstNr[0]) || (9740 == GlobalFiModInstNr[1]) || (9740 == GlobalFiModInstNr[2]) || (9740 == GlobalFiModInstNr[3]))));
	Tile mesh_11_18(
		.clock(clock),
		.io_in_a_0(r_370_0),
		.io_in_b_0(b_587_0),
		.io_in_d_0(b_1611_0),
		.io_in_control_0_dataflow(mesh_11_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2635_0),
		.io_in_last_0(r_3659_0),
		.io_in_valid_0(r_1611_0),
		.io_out_a_0(_mesh_11_18_io_out_a_0),
		.io_out_c_0(_mesh_11_18_io_out_c_0),
		.io_out_b_0(_mesh_11_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_18_io_out_id_0),
		.io_out_last_0(_mesh_11_18_io_out_last_0),
		.io_out_valid_0(_mesh_11_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9741 == GlobalFiModInstNr[0]) || (9741 == GlobalFiModInstNr[1]) || (9741 == GlobalFiModInstNr[2]) || (9741 == GlobalFiModInstNr[3]))));
	Tile mesh_11_19(
		.clock(clock),
		.io_in_a_0(r_371_0),
		.io_in_b_0(b_619_0),
		.io_in_d_0(b_1643_0),
		.io_in_control_0_dataflow(mesh_11_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2667_0),
		.io_in_last_0(r_3691_0),
		.io_in_valid_0(r_1643_0),
		.io_out_a_0(_mesh_11_19_io_out_a_0),
		.io_out_c_0(_mesh_11_19_io_out_c_0),
		.io_out_b_0(_mesh_11_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_19_io_out_id_0),
		.io_out_last_0(_mesh_11_19_io_out_last_0),
		.io_out_valid_0(_mesh_11_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9742 == GlobalFiModInstNr[0]) || (9742 == GlobalFiModInstNr[1]) || (9742 == GlobalFiModInstNr[2]) || (9742 == GlobalFiModInstNr[3]))));
	Tile mesh_11_20(
		.clock(clock),
		.io_in_a_0(r_372_0),
		.io_in_b_0(b_651_0),
		.io_in_d_0(b_1675_0),
		.io_in_control_0_dataflow(mesh_11_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2699_0),
		.io_in_last_0(r_3723_0),
		.io_in_valid_0(r_1675_0),
		.io_out_a_0(_mesh_11_20_io_out_a_0),
		.io_out_c_0(_mesh_11_20_io_out_c_0),
		.io_out_b_0(_mesh_11_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_20_io_out_id_0),
		.io_out_last_0(_mesh_11_20_io_out_last_0),
		.io_out_valid_0(_mesh_11_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9743 == GlobalFiModInstNr[0]) || (9743 == GlobalFiModInstNr[1]) || (9743 == GlobalFiModInstNr[2]) || (9743 == GlobalFiModInstNr[3]))));
	Tile mesh_11_21(
		.clock(clock),
		.io_in_a_0(r_373_0),
		.io_in_b_0(b_683_0),
		.io_in_d_0(b_1707_0),
		.io_in_control_0_dataflow(mesh_11_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2731_0),
		.io_in_last_0(r_3755_0),
		.io_in_valid_0(r_1707_0),
		.io_out_a_0(_mesh_11_21_io_out_a_0),
		.io_out_c_0(_mesh_11_21_io_out_c_0),
		.io_out_b_0(_mesh_11_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_21_io_out_id_0),
		.io_out_last_0(_mesh_11_21_io_out_last_0),
		.io_out_valid_0(_mesh_11_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9744 == GlobalFiModInstNr[0]) || (9744 == GlobalFiModInstNr[1]) || (9744 == GlobalFiModInstNr[2]) || (9744 == GlobalFiModInstNr[3]))));
	Tile mesh_11_22(
		.clock(clock),
		.io_in_a_0(r_374_0),
		.io_in_b_0(b_715_0),
		.io_in_d_0(b_1739_0),
		.io_in_control_0_dataflow(mesh_11_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2763_0),
		.io_in_last_0(r_3787_0),
		.io_in_valid_0(r_1739_0),
		.io_out_a_0(_mesh_11_22_io_out_a_0),
		.io_out_c_0(_mesh_11_22_io_out_c_0),
		.io_out_b_0(_mesh_11_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_22_io_out_id_0),
		.io_out_last_0(_mesh_11_22_io_out_last_0),
		.io_out_valid_0(_mesh_11_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9745 == GlobalFiModInstNr[0]) || (9745 == GlobalFiModInstNr[1]) || (9745 == GlobalFiModInstNr[2]) || (9745 == GlobalFiModInstNr[3]))));
	Tile mesh_11_23(
		.clock(clock),
		.io_in_a_0(r_375_0),
		.io_in_b_0(b_747_0),
		.io_in_d_0(b_1771_0),
		.io_in_control_0_dataflow(mesh_11_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2795_0),
		.io_in_last_0(r_3819_0),
		.io_in_valid_0(r_1771_0),
		.io_out_a_0(_mesh_11_23_io_out_a_0),
		.io_out_c_0(_mesh_11_23_io_out_c_0),
		.io_out_b_0(_mesh_11_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_23_io_out_id_0),
		.io_out_last_0(_mesh_11_23_io_out_last_0),
		.io_out_valid_0(_mesh_11_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9746 == GlobalFiModInstNr[0]) || (9746 == GlobalFiModInstNr[1]) || (9746 == GlobalFiModInstNr[2]) || (9746 == GlobalFiModInstNr[3]))));
	Tile mesh_11_24(
		.clock(clock),
		.io_in_a_0(r_376_0),
		.io_in_b_0(b_779_0),
		.io_in_d_0(b_1803_0),
		.io_in_control_0_dataflow(mesh_11_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2827_0),
		.io_in_last_0(r_3851_0),
		.io_in_valid_0(r_1803_0),
		.io_out_a_0(_mesh_11_24_io_out_a_0),
		.io_out_c_0(_mesh_11_24_io_out_c_0),
		.io_out_b_0(_mesh_11_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_24_io_out_id_0),
		.io_out_last_0(_mesh_11_24_io_out_last_0),
		.io_out_valid_0(_mesh_11_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9747 == GlobalFiModInstNr[0]) || (9747 == GlobalFiModInstNr[1]) || (9747 == GlobalFiModInstNr[2]) || (9747 == GlobalFiModInstNr[3]))));
	Tile mesh_11_25(
		.clock(clock),
		.io_in_a_0(r_377_0),
		.io_in_b_0(b_811_0),
		.io_in_d_0(b_1835_0),
		.io_in_control_0_dataflow(mesh_11_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2859_0),
		.io_in_last_0(r_3883_0),
		.io_in_valid_0(r_1835_0),
		.io_out_a_0(_mesh_11_25_io_out_a_0),
		.io_out_c_0(_mesh_11_25_io_out_c_0),
		.io_out_b_0(_mesh_11_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_25_io_out_id_0),
		.io_out_last_0(_mesh_11_25_io_out_last_0),
		.io_out_valid_0(_mesh_11_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9748 == GlobalFiModInstNr[0]) || (9748 == GlobalFiModInstNr[1]) || (9748 == GlobalFiModInstNr[2]) || (9748 == GlobalFiModInstNr[3]))));
	Tile mesh_11_26(
		.clock(clock),
		.io_in_a_0(r_378_0),
		.io_in_b_0(b_843_0),
		.io_in_d_0(b_1867_0),
		.io_in_control_0_dataflow(mesh_11_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2891_0),
		.io_in_last_0(r_3915_0),
		.io_in_valid_0(r_1867_0),
		.io_out_a_0(_mesh_11_26_io_out_a_0),
		.io_out_c_0(_mesh_11_26_io_out_c_0),
		.io_out_b_0(_mesh_11_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_26_io_out_id_0),
		.io_out_last_0(_mesh_11_26_io_out_last_0),
		.io_out_valid_0(_mesh_11_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9749 == GlobalFiModInstNr[0]) || (9749 == GlobalFiModInstNr[1]) || (9749 == GlobalFiModInstNr[2]) || (9749 == GlobalFiModInstNr[3]))));
	Tile mesh_11_27(
		.clock(clock),
		.io_in_a_0(r_379_0),
		.io_in_b_0(b_875_0),
		.io_in_d_0(b_1899_0),
		.io_in_control_0_dataflow(mesh_11_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2923_0),
		.io_in_last_0(r_3947_0),
		.io_in_valid_0(r_1899_0),
		.io_out_a_0(_mesh_11_27_io_out_a_0),
		.io_out_c_0(_mesh_11_27_io_out_c_0),
		.io_out_b_0(_mesh_11_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_27_io_out_id_0),
		.io_out_last_0(_mesh_11_27_io_out_last_0),
		.io_out_valid_0(_mesh_11_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9750 == GlobalFiModInstNr[0]) || (9750 == GlobalFiModInstNr[1]) || (9750 == GlobalFiModInstNr[2]) || (9750 == GlobalFiModInstNr[3]))));
	Tile mesh_11_28(
		.clock(clock),
		.io_in_a_0(r_380_0),
		.io_in_b_0(b_907_0),
		.io_in_d_0(b_1931_0),
		.io_in_control_0_dataflow(mesh_11_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2955_0),
		.io_in_last_0(r_3979_0),
		.io_in_valid_0(r_1931_0),
		.io_out_a_0(_mesh_11_28_io_out_a_0),
		.io_out_c_0(_mesh_11_28_io_out_c_0),
		.io_out_b_0(_mesh_11_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_28_io_out_id_0),
		.io_out_last_0(_mesh_11_28_io_out_last_0),
		.io_out_valid_0(_mesh_11_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9751 == GlobalFiModInstNr[0]) || (9751 == GlobalFiModInstNr[1]) || (9751 == GlobalFiModInstNr[2]) || (9751 == GlobalFiModInstNr[3]))));
	Tile mesh_11_29(
		.clock(clock),
		.io_in_a_0(r_381_0),
		.io_in_b_0(b_939_0),
		.io_in_d_0(b_1963_0),
		.io_in_control_0_dataflow(mesh_11_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2987_0),
		.io_in_last_0(r_4011_0),
		.io_in_valid_0(r_1963_0),
		.io_out_a_0(_mesh_11_29_io_out_a_0),
		.io_out_c_0(_mesh_11_29_io_out_c_0),
		.io_out_b_0(_mesh_11_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_29_io_out_id_0),
		.io_out_last_0(_mesh_11_29_io_out_last_0),
		.io_out_valid_0(_mesh_11_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9752 == GlobalFiModInstNr[0]) || (9752 == GlobalFiModInstNr[1]) || (9752 == GlobalFiModInstNr[2]) || (9752 == GlobalFiModInstNr[3]))));
	Tile mesh_11_30(
		.clock(clock),
		.io_in_a_0(r_382_0),
		.io_in_b_0(b_971_0),
		.io_in_d_0(b_1995_0),
		.io_in_control_0_dataflow(mesh_11_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3019_0),
		.io_in_last_0(r_4043_0),
		.io_in_valid_0(r_1995_0),
		.io_out_a_0(_mesh_11_30_io_out_a_0),
		.io_out_c_0(_mesh_11_30_io_out_c_0),
		.io_out_b_0(_mesh_11_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_30_io_out_id_0),
		.io_out_last_0(_mesh_11_30_io_out_last_0),
		.io_out_valid_0(_mesh_11_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9753 == GlobalFiModInstNr[0]) || (9753 == GlobalFiModInstNr[1]) || (9753 == GlobalFiModInstNr[2]) || (9753 == GlobalFiModInstNr[3]))));
	Tile mesh_11_31(
		.clock(clock),
		.io_in_a_0(r_383_0),
		.io_in_b_0(b_1003_0),
		.io_in_d_0(b_2027_0),
		.io_in_control_0_dataflow(mesh_11_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_11_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_11_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3051_0),
		.io_in_last_0(r_4075_0),
		.io_in_valid_0(r_2027_0),
		.io_out_a_0(_mesh_11_31_io_out_a_0),
		.io_out_c_0(_mesh_11_31_io_out_c_0),
		.io_out_b_0(_mesh_11_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_11_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_11_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_11_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_11_31_io_out_id_0),
		.io_out_last_0(_mesh_11_31_io_out_last_0),
		.io_out_valid_0(_mesh_11_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9754 == GlobalFiModInstNr[0]) || (9754 == GlobalFiModInstNr[1]) || (9754 == GlobalFiModInstNr[2]) || (9754 == GlobalFiModInstNr[3]))));
	Tile mesh_12_0(
		.clock(clock),
		.io_in_a_0(r_384_0),
		.io_in_b_0(b_12_0),
		.io_in_d_0(b_1036_0),
		.io_in_control_0_dataflow(mesh_12_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2060_0),
		.io_in_last_0(r_3084_0),
		.io_in_valid_0(r_1036_0),
		.io_out_a_0(_mesh_12_0_io_out_a_0),
		.io_out_c_0(_mesh_12_0_io_out_c_0),
		.io_out_b_0(_mesh_12_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_0_io_out_id_0),
		.io_out_last_0(_mesh_12_0_io_out_last_0),
		.io_out_valid_0(_mesh_12_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9755 == GlobalFiModInstNr[0]) || (9755 == GlobalFiModInstNr[1]) || (9755 == GlobalFiModInstNr[2]) || (9755 == GlobalFiModInstNr[3]))));
	Tile mesh_12_1(
		.clock(clock),
		.io_in_a_0(r_385_0),
		.io_in_b_0(b_44_0),
		.io_in_d_0(b_1068_0),
		.io_in_control_0_dataflow(mesh_12_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2092_0),
		.io_in_last_0(r_3116_0),
		.io_in_valid_0(r_1068_0),
		.io_out_a_0(_mesh_12_1_io_out_a_0),
		.io_out_c_0(_mesh_12_1_io_out_c_0),
		.io_out_b_0(_mesh_12_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_1_io_out_id_0),
		.io_out_last_0(_mesh_12_1_io_out_last_0),
		.io_out_valid_0(_mesh_12_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9756 == GlobalFiModInstNr[0]) || (9756 == GlobalFiModInstNr[1]) || (9756 == GlobalFiModInstNr[2]) || (9756 == GlobalFiModInstNr[3]))));
	Tile mesh_12_2(
		.clock(clock),
		.io_in_a_0(r_386_0),
		.io_in_b_0(b_76_0),
		.io_in_d_0(b_1100_0),
		.io_in_control_0_dataflow(mesh_12_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2124_0),
		.io_in_last_0(r_3148_0),
		.io_in_valid_0(r_1100_0),
		.io_out_a_0(_mesh_12_2_io_out_a_0),
		.io_out_c_0(_mesh_12_2_io_out_c_0),
		.io_out_b_0(_mesh_12_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_2_io_out_id_0),
		.io_out_last_0(_mesh_12_2_io_out_last_0),
		.io_out_valid_0(_mesh_12_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9757 == GlobalFiModInstNr[0]) || (9757 == GlobalFiModInstNr[1]) || (9757 == GlobalFiModInstNr[2]) || (9757 == GlobalFiModInstNr[3]))));
	Tile mesh_12_3(
		.clock(clock),
		.io_in_a_0(r_387_0),
		.io_in_b_0(b_108_0),
		.io_in_d_0(b_1132_0),
		.io_in_control_0_dataflow(mesh_12_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2156_0),
		.io_in_last_0(r_3180_0),
		.io_in_valid_0(r_1132_0),
		.io_out_a_0(_mesh_12_3_io_out_a_0),
		.io_out_c_0(_mesh_12_3_io_out_c_0),
		.io_out_b_0(_mesh_12_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_3_io_out_id_0),
		.io_out_last_0(_mesh_12_3_io_out_last_0),
		.io_out_valid_0(_mesh_12_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9758 == GlobalFiModInstNr[0]) || (9758 == GlobalFiModInstNr[1]) || (9758 == GlobalFiModInstNr[2]) || (9758 == GlobalFiModInstNr[3]))));
	Tile mesh_12_4(
		.clock(clock),
		.io_in_a_0(r_388_0),
		.io_in_b_0(b_140_0),
		.io_in_d_0(b_1164_0),
		.io_in_control_0_dataflow(mesh_12_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2188_0),
		.io_in_last_0(r_3212_0),
		.io_in_valid_0(r_1164_0),
		.io_out_a_0(_mesh_12_4_io_out_a_0),
		.io_out_c_0(_mesh_12_4_io_out_c_0),
		.io_out_b_0(_mesh_12_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_4_io_out_id_0),
		.io_out_last_0(_mesh_12_4_io_out_last_0),
		.io_out_valid_0(_mesh_12_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9759 == GlobalFiModInstNr[0]) || (9759 == GlobalFiModInstNr[1]) || (9759 == GlobalFiModInstNr[2]) || (9759 == GlobalFiModInstNr[3]))));
	Tile mesh_12_5(
		.clock(clock),
		.io_in_a_0(r_389_0),
		.io_in_b_0(b_172_0),
		.io_in_d_0(b_1196_0),
		.io_in_control_0_dataflow(mesh_12_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2220_0),
		.io_in_last_0(r_3244_0),
		.io_in_valid_0(r_1196_0),
		.io_out_a_0(_mesh_12_5_io_out_a_0),
		.io_out_c_0(_mesh_12_5_io_out_c_0),
		.io_out_b_0(_mesh_12_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_5_io_out_id_0),
		.io_out_last_0(_mesh_12_5_io_out_last_0),
		.io_out_valid_0(_mesh_12_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9760 == GlobalFiModInstNr[0]) || (9760 == GlobalFiModInstNr[1]) || (9760 == GlobalFiModInstNr[2]) || (9760 == GlobalFiModInstNr[3]))));
	Tile mesh_12_6(
		.clock(clock),
		.io_in_a_0(r_390_0),
		.io_in_b_0(b_204_0),
		.io_in_d_0(b_1228_0),
		.io_in_control_0_dataflow(mesh_12_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2252_0),
		.io_in_last_0(r_3276_0),
		.io_in_valid_0(r_1228_0),
		.io_out_a_0(_mesh_12_6_io_out_a_0),
		.io_out_c_0(_mesh_12_6_io_out_c_0),
		.io_out_b_0(_mesh_12_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_6_io_out_id_0),
		.io_out_last_0(_mesh_12_6_io_out_last_0),
		.io_out_valid_0(_mesh_12_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9761 == GlobalFiModInstNr[0]) || (9761 == GlobalFiModInstNr[1]) || (9761 == GlobalFiModInstNr[2]) || (9761 == GlobalFiModInstNr[3]))));
	Tile mesh_12_7(
		.clock(clock),
		.io_in_a_0(r_391_0),
		.io_in_b_0(b_236_0),
		.io_in_d_0(b_1260_0),
		.io_in_control_0_dataflow(mesh_12_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2284_0),
		.io_in_last_0(r_3308_0),
		.io_in_valid_0(r_1260_0),
		.io_out_a_0(_mesh_12_7_io_out_a_0),
		.io_out_c_0(_mesh_12_7_io_out_c_0),
		.io_out_b_0(_mesh_12_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_7_io_out_id_0),
		.io_out_last_0(_mesh_12_7_io_out_last_0),
		.io_out_valid_0(_mesh_12_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9762 == GlobalFiModInstNr[0]) || (9762 == GlobalFiModInstNr[1]) || (9762 == GlobalFiModInstNr[2]) || (9762 == GlobalFiModInstNr[3]))));
	Tile mesh_12_8(
		.clock(clock),
		.io_in_a_0(r_392_0),
		.io_in_b_0(b_268_0),
		.io_in_d_0(b_1292_0),
		.io_in_control_0_dataflow(mesh_12_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2316_0),
		.io_in_last_0(r_3340_0),
		.io_in_valid_0(r_1292_0),
		.io_out_a_0(_mesh_12_8_io_out_a_0),
		.io_out_c_0(_mesh_12_8_io_out_c_0),
		.io_out_b_0(_mesh_12_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_8_io_out_id_0),
		.io_out_last_0(_mesh_12_8_io_out_last_0),
		.io_out_valid_0(_mesh_12_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9763 == GlobalFiModInstNr[0]) || (9763 == GlobalFiModInstNr[1]) || (9763 == GlobalFiModInstNr[2]) || (9763 == GlobalFiModInstNr[3]))));
	Tile mesh_12_9(
		.clock(clock),
		.io_in_a_0(r_393_0),
		.io_in_b_0(b_300_0),
		.io_in_d_0(b_1324_0),
		.io_in_control_0_dataflow(mesh_12_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2348_0),
		.io_in_last_0(r_3372_0),
		.io_in_valid_0(r_1324_0),
		.io_out_a_0(_mesh_12_9_io_out_a_0),
		.io_out_c_0(_mesh_12_9_io_out_c_0),
		.io_out_b_0(_mesh_12_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_9_io_out_id_0),
		.io_out_last_0(_mesh_12_9_io_out_last_0),
		.io_out_valid_0(_mesh_12_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9764 == GlobalFiModInstNr[0]) || (9764 == GlobalFiModInstNr[1]) || (9764 == GlobalFiModInstNr[2]) || (9764 == GlobalFiModInstNr[3]))));
	Tile mesh_12_10(
		.clock(clock),
		.io_in_a_0(r_394_0),
		.io_in_b_0(b_332_0),
		.io_in_d_0(b_1356_0),
		.io_in_control_0_dataflow(mesh_12_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2380_0),
		.io_in_last_0(r_3404_0),
		.io_in_valid_0(r_1356_0),
		.io_out_a_0(_mesh_12_10_io_out_a_0),
		.io_out_c_0(_mesh_12_10_io_out_c_0),
		.io_out_b_0(_mesh_12_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_10_io_out_id_0),
		.io_out_last_0(_mesh_12_10_io_out_last_0),
		.io_out_valid_0(_mesh_12_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9765 == GlobalFiModInstNr[0]) || (9765 == GlobalFiModInstNr[1]) || (9765 == GlobalFiModInstNr[2]) || (9765 == GlobalFiModInstNr[3]))));
	Tile mesh_12_11(
		.clock(clock),
		.io_in_a_0(r_395_0),
		.io_in_b_0(b_364_0),
		.io_in_d_0(b_1388_0),
		.io_in_control_0_dataflow(mesh_12_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2412_0),
		.io_in_last_0(r_3436_0),
		.io_in_valid_0(r_1388_0),
		.io_out_a_0(_mesh_12_11_io_out_a_0),
		.io_out_c_0(_mesh_12_11_io_out_c_0),
		.io_out_b_0(_mesh_12_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_11_io_out_id_0),
		.io_out_last_0(_mesh_12_11_io_out_last_0),
		.io_out_valid_0(_mesh_12_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9766 == GlobalFiModInstNr[0]) || (9766 == GlobalFiModInstNr[1]) || (9766 == GlobalFiModInstNr[2]) || (9766 == GlobalFiModInstNr[3]))));
	Tile mesh_12_12(
		.clock(clock),
		.io_in_a_0(r_396_0),
		.io_in_b_0(b_396_0),
		.io_in_d_0(b_1420_0),
		.io_in_control_0_dataflow(mesh_12_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2444_0),
		.io_in_last_0(r_3468_0),
		.io_in_valid_0(r_1420_0),
		.io_out_a_0(_mesh_12_12_io_out_a_0),
		.io_out_c_0(_mesh_12_12_io_out_c_0),
		.io_out_b_0(_mesh_12_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_12_io_out_id_0),
		.io_out_last_0(_mesh_12_12_io_out_last_0),
		.io_out_valid_0(_mesh_12_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9767 == GlobalFiModInstNr[0]) || (9767 == GlobalFiModInstNr[1]) || (9767 == GlobalFiModInstNr[2]) || (9767 == GlobalFiModInstNr[3]))));
	Tile mesh_12_13(
		.clock(clock),
		.io_in_a_0(r_397_0),
		.io_in_b_0(b_428_0),
		.io_in_d_0(b_1452_0),
		.io_in_control_0_dataflow(mesh_12_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2476_0),
		.io_in_last_0(r_3500_0),
		.io_in_valid_0(r_1452_0),
		.io_out_a_0(_mesh_12_13_io_out_a_0),
		.io_out_c_0(_mesh_12_13_io_out_c_0),
		.io_out_b_0(_mesh_12_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_13_io_out_id_0),
		.io_out_last_0(_mesh_12_13_io_out_last_0),
		.io_out_valid_0(_mesh_12_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9768 == GlobalFiModInstNr[0]) || (9768 == GlobalFiModInstNr[1]) || (9768 == GlobalFiModInstNr[2]) || (9768 == GlobalFiModInstNr[3]))));
	Tile mesh_12_14(
		.clock(clock),
		.io_in_a_0(r_398_0),
		.io_in_b_0(b_460_0),
		.io_in_d_0(b_1484_0),
		.io_in_control_0_dataflow(mesh_12_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2508_0),
		.io_in_last_0(r_3532_0),
		.io_in_valid_0(r_1484_0),
		.io_out_a_0(_mesh_12_14_io_out_a_0),
		.io_out_c_0(_mesh_12_14_io_out_c_0),
		.io_out_b_0(_mesh_12_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_14_io_out_id_0),
		.io_out_last_0(_mesh_12_14_io_out_last_0),
		.io_out_valid_0(_mesh_12_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9769 == GlobalFiModInstNr[0]) || (9769 == GlobalFiModInstNr[1]) || (9769 == GlobalFiModInstNr[2]) || (9769 == GlobalFiModInstNr[3]))));
	Tile mesh_12_15(
		.clock(clock),
		.io_in_a_0(r_399_0),
		.io_in_b_0(b_492_0),
		.io_in_d_0(b_1516_0),
		.io_in_control_0_dataflow(mesh_12_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2540_0),
		.io_in_last_0(r_3564_0),
		.io_in_valid_0(r_1516_0),
		.io_out_a_0(_mesh_12_15_io_out_a_0),
		.io_out_c_0(_mesh_12_15_io_out_c_0),
		.io_out_b_0(_mesh_12_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_15_io_out_id_0),
		.io_out_last_0(_mesh_12_15_io_out_last_0),
		.io_out_valid_0(_mesh_12_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9770 == GlobalFiModInstNr[0]) || (9770 == GlobalFiModInstNr[1]) || (9770 == GlobalFiModInstNr[2]) || (9770 == GlobalFiModInstNr[3]))));
	Tile mesh_12_16(
		.clock(clock),
		.io_in_a_0(r_400_0),
		.io_in_b_0(b_524_0),
		.io_in_d_0(b_1548_0),
		.io_in_control_0_dataflow(mesh_12_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2572_0),
		.io_in_last_0(r_3596_0),
		.io_in_valid_0(r_1548_0),
		.io_out_a_0(_mesh_12_16_io_out_a_0),
		.io_out_c_0(_mesh_12_16_io_out_c_0),
		.io_out_b_0(_mesh_12_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_16_io_out_id_0),
		.io_out_last_0(_mesh_12_16_io_out_last_0),
		.io_out_valid_0(_mesh_12_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9771 == GlobalFiModInstNr[0]) || (9771 == GlobalFiModInstNr[1]) || (9771 == GlobalFiModInstNr[2]) || (9771 == GlobalFiModInstNr[3]))));
	Tile mesh_12_17(
		.clock(clock),
		.io_in_a_0(r_401_0),
		.io_in_b_0(b_556_0),
		.io_in_d_0(b_1580_0),
		.io_in_control_0_dataflow(mesh_12_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2604_0),
		.io_in_last_0(r_3628_0),
		.io_in_valid_0(r_1580_0),
		.io_out_a_0(_mesh_12_17_io_out_a_0),
		.io_out_c_0(_mesh_12_17_io_out_c_0),
		.io_out_b_0(_mesh_12_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_17_io_out_id_0),
		.io_out_last_0(_mesh_12_17_io_out_last_0),
		.io_out_valid_0(_mesh_12_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9772 == GlobalFiModInstNr[0]) || (9772 == GlobalFiModInstNr[1]) || (9772 == GlobalFiModInstNr[2]) || (9772 == GlobalFiModInstNr[3]))));
	Tile mesh_12_18(
		.clock(clock),
		.io_in_a_0(r_402_0),
		.io_in_b_0(b_588_0),
		.io_in_d_0(b_1612_0),
		.io_in_control_0_dataflow(mesh_12_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2636_0),
		.io_in_last_0(r_3660_0),
		.io_in_valid_0(r_1612_0),
		.io_out_a_0(_mesh_12_18_io_out_a_0),
		.io_out_c_0(_mesh_12_18_io_out_c_0),
		.io_out_b_0(_mesh_12_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_18_io_out_id_0),
		.io_out_last_0(_mesh_12_18_io_out_last_0),
		.io_out_valid_0(_mesh_12_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9773 == GlobalFiModInstNr[0]) || (9773 == GlobalFiModInstNr[1]) || (9773 == GlobalFiModInstNr[2]) || (9773 == GlobalFiModInstNr[3]))));
	Tile mesh_12_19(
		.clock(clock),
		.io_in_a_0(r_403_0),
		.io_in_b_0(b_620_0),
		.io_in_d_0(b_1644_0),
		.io_in_control_0_dataflow(mesh_12_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2668_0),
		.io_in_last_0(r_3692_0),
		.io_in_valid_0(r_1644_0),
		.io_out_a_0(_mesh_12_19_io_out_a_0),
		.io_out_c_0(_mesh_12_19_io_out_c_0),
		.io_out_b_0(_mesh_12_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_19_io_out_id_0),
		.io_out_last_0(_mesh_12_19_io_out_last_0),
		.io_out_valid_0(_mesh_12_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9774 == GlobalFiModInstNr[0]) || (9774 == GlobalFiModInstNr[1]) || (9774 == GlobalFiModInstNr[2]) || (9774 == GlobalFiModInstNr[3]))));
	Tile mesh_12_20(
		.clock(clock),
		.io_in_a_0(r_404_0),
		.io_in_b_0(b_652_0),
		.io_in_d_0(b_1676_0),
		.io_in_control_0_dataflow(mesh_12_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2700_0),
		.io_in_last_0(r_3724_0),
		.io_in_valid_0(r_1676_0),
		.io_out_a_0(_mesh_12_20_io_out_a_0),
		.io_out_c_0(_mesh_12_20_io_out_c_0),
		.io_out_b_0(_mesh_12_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_20_io_out_id_0),
		.io_out_last_0(_mesh_12_20_io_out_last_0),
		.io_out_valid_0(_mesh_12_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9775 == GlobalFiModInstNr[0]) || (9775 == GlobalFiModInstNr[1]) || (9775 == GlobalFiModInstNr[2]) || (9775 == GlobalFiModInstNr[3]))));
	Tile mesh_12_21(
		.clock(clock),
		.io_in_a_0(r_405_0),
		.io_in_b_0(b_684_0),
		.io_in_d_0(b_1708_0),
		.io_in_control_0_dataflow(mesh_12_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2732_0),
		.io_in_last_0(r_3756_0),
		.io_in_valid_0(r_1708_0),
		.io_out_a_0(_mesh_12_21_io_out_a_0),
		.io_out_c_0(_mesh_12_21_io_out_c_0),
		.io_out_b_0(_mesh_12_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_21_io_out_id_0),
		.io_out_last_0(_mesh_12_21_io_out_last_0),
		.io_out_valid_0(_mesh_12_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9776 == GlobalFiModInstNr[0]) || (9776 == GlobalFiModInstNr[1]) || (9776 == GlobalFiModInstNr[2]) || (9776 == GlobalFiModInstNr[3]))));
	Tile mesh_12_22(
		.clock(clock),
		.io_in_a_0(r_406_0),
		.io_in_b_0(b_716_0),
		.io_in_d_0(b_1740_0),
		.io_in_control_0_dataflow(mesh_12_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2764_0),
		.io_in_last_0(r_3788_0),
		.io_in_valid_0(r_1740_0),
		.io_out_a_0(_mesh_12_22_io_out_a_0),
		.io_out_c_0(_mesh_12_22_io_out_c_0),
		.io_out_b_0(_mesh_12_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_22_io_out_id_0),
		.io_out_last_0(_mesh_12_22_io_out_last_0),
		.io_out_valid_0(_mesh_12_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9777 == GlobalFiModInstNr[0]) || (9777 == GlobalFiModInstNr[1]) || (9777 == GlobalFiModInstNr[2]) || (9777 == GlobalFiModInstNr[3]))));
	Tile mesh_12_23(
		.clock(clock),
		.io_in_a_0(r_407_0),
		.io_in_b_0(b_748_0),
		.io_in_d_0(b_1772_0),
		.io_in_control_0_dataflow(mesh_12_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2796_0),
		.io_in_last_0(r_3820_0),
		.io_in_valid_0(r_1772_0),
		.io_out_a_0(_mesh_12_23_io_out_a_0),
		.io_out_c_0(_mesh_12_23_io_out_c_0),
		.io_out_b_0(_mesh_12_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_23_io_out_id_0),
		.io_out_last_0(_mesh_12_23_io_out_last_0),
		.io_out_valid_0(_mesh_12_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9778 == GlobalFiModInstNr[0]) || (9778 == GlobalFiModInstNr[1]) || (9778 == GlobalFiModInstNr[2]) || (9778 == GlobalFiModInstNr[3]))));
	Tile mesh_12_24(
		.clock(clock),
		.io_in_a_0(r_408_0),
		.io_in_b_0(b_780_0),
		.io_in_d_0(b_1804_0),
		.io_in_control_0_dataflow(mesh_12_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2828_0),
		.io_in_last_0(r_3852_0),
		.io_in_valid_0(r_1804_0),
		.io_out_a_0(_mesh_12_24_io_out_a_0),
		.io_out_c_0(_mesh_12_24_io_out_c_0),
		.io_out_b_0(_mesh_12_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_24_io_out_id_0),
		.io_out_last_0(_mesh_12_24_io_out_last_0),
		.io_out_valid_0(_mesh_12_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9779 == GlobalFiModInstNr[0]) || (9779 == GlobalFiModInstNr[1]) || (9779 == GlobalFiModInstNr[2]) || (9779 == GlobalFiModInstNr[3]))));
	Tile mesh_12_25(
		.clock(clock),
		.io_in_a_0(r_409_0),
		.io_in_b_0(b_812_0),
		.io_in_d_0(b_1836_0),
		.io_in_control_0_dataflow(mesh_12_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2860_0),
		.io_in_last_0(r_3884_0),
		.io_in_valid_0(r_1836_0),
		.io_out_a_0(_mesh_12_25_io_out_a_0),
		.io_out_c_0(_mesh_12_25_io_out_c_0),
		.io_out_b_0(_mesh_12_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_25_io_out_id_0),
		.io_out_last_0(_mesh_12_25_io_out_last_0),
		.io_out_valid_0(_mesh_12_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9780 == GlobalFiModInstNr[0]) || (9780 == GlobalFiModInstNr[1]) || (9780 == GlobalFiModInstNr[2]) || (9780 == GlobalFiModInstNr[3]))));
	Tile mesh_12_26(
		.clock(clock),
		.io_in_a_0(r_410_0),
		.io_in_b_0(b_844_0),
		.io_in_d_0(b_1868_0),
		.io_in_control_0_dataflow(mesh_12_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2892_0),
		.io_in_last_0(r_3916_0),
		.io_in_valid_0(r_1868_0),
		.io_out_a_0(_mesh_12_26_io_out_a_0),
		.io_out_c_0(_mesh_12_26_io_out_c_0),
		.io_out_b_0(_mesh_12_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_26_io_out_id_0),
		.io_out_last_0(_mesh_12_26_io_out_last_0),
		.io_out_valid_0(_mesh_12_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9781 == GlobalFiModInstNr[0]) || (9781 == GlobalFiModInstNr[1]) || (9781 == GlobalFiModInstNr[2]) || (9781 == GlobalFiModInstNr[3]))));
	Tile mesh_12_27(
		.clock(clock),
		.io_in_a_0(r_411_0),
		.io_in_b_0(b_876_0),
		.io_in_d_0(b_1900_0),
		.io_in_control_0_dataflow(mesh_12_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2924_0),
		.io_in_last_0(r_3948_0),
		.io_in_valid_0(r_1900_0),
		.io_out_a_0(_mesh_12_27_io_out_a_0),
		.io_out_c_0(_mesh_12_27_io_out_c_0),
		.io_out_b_0(_mesh_12_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_27_io_out_id_0),
		.io_out_last_0(_mesh_12_27_io_out_last_0),
		.io_out_valid_0(_mesh_12_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9782 == GlobalFiModInstNr[0]) || (9782 == GlobalFiModInstNr[1]) || (9782 == GlobalFiModInstNr[2]) || (9782 == GlobalFiModInstNr[3]))));
	Tile mesh_12_28(
		.clock(clock),
		.io_in_a_0(r_412_0),
		.io_in_b_0(b_908_0),
		.io_in_d_0(b_1932_0),
		.io_in_control_0_dataflow(mesh_12_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2956_0),
		.io_in_last_0(r_3980_0),
		.io_in_valid_0(r_1932_0),
		.io_out_a_0(_mesh_12_28_io_out_a_0),
		.io_out_c_0(_mesh_12_28_io_out_c_0),
		.io_out_b_0(_mesh_12_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_28_io_out_id_0),
		.io_out_last_0(_mesh_12_28_io_out_last_0),
		.io_out_valid_0(_mesh_12_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9783 == GlobalFiModInstNr[0]) || (9783 == GlobalFiModInstNr[1]) || (9783 == GlobalFiModInstNr[2]) || (9783 == GlobalFiModInstNr[3]))));
	Tile mesh_12_29(
		.clock(clock),
		.io_in_a_0(r_413_0),
		.io_in_b_0(b_940_0),
		.io_in_d_0(b_1964_0),
		.io_in_control_0_dataflow(mesh_12_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2988_0),
		.io_in_last_0(r_4012_0),
		.io_in_valid_0(r_1964_0),
		.io_out_a_0(_mesh_12_29_io_out_a_0),
		.io_out_c_0(_mesh_12_29_io_out_c_0),
		.io_out_b_0(_mesh_12_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_29_io_out_id_0),
		.io_out_last_0(_mesh_12_29_io_out_last_0),
		.io_out_valid_0(_mesh_12_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9784 == GlobalFiModInstNr[0]) || (9784 == GlobalFiModInstNr[1]) || (9784 == GlobalFiModInstNr[2]) || (9784 == GlobalFiModInstNr[3]))));
	Tile mesh_12_30(
		.clock(clock),
		.io_in_a_0(r_414_0),
		.io_in_b_0(b_972_0),
		.io_in_d_0(b_1996_0),
		.io_in_control_0_dataflow(mesh_12_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3020_0),
		.io_in_last_0(r_4044_0),
		.io_in_valid_0(r_1996_0),
		.io_out_a_0(_mesh_12_30_io_out_a_0),
		.io_out_c_0(_mesh_12_30_io_out_c_0),
		.io_out_b_0(_mesh_12_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_30_io_out_id_0),
		.io_out_last_0(_mesh_12_30_io_out_last_0),
		.io_out_valid_0(_mesh_12_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9785 == GlobalFiModInstNr[0]) || (9785 == GlobalFiModInstNr[1]) || (9785 == GlobalFiModInstNr[2]) || (9785 == GlobalFiModInstNr[3]))));
	Tile mesh_12_31(
		.clock(clock),
		.io_in_a_0(r_415_0),
		.io_in_b_0(b_1004_0),
		.io_in_d_0(b_2028_0),
		.io_in_control_0_dataflow(mesh_12_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_12_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_12_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3052_0),
		.io_in_last_0(r_4076_0),
		.io_in_valid_0(r_2028_0),
		.io_out_a_0(_mesh_12_31_io_out_a_0),
		.io_out_c_0(_mesh_12_31_io_out_c_0),
		.io_out_b_0(_mesh_12_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_12_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_12_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_12_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_12_31_io_out_id_0),
		.io_out_last_0(_mesh_12_31_io_out_last_0),
		.io_out_valid_0(_mesh_12_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9786 == GlobalFiModInstNr[0]) || (9786 == GlobalFiModInstNr[1]) || (9786 == GlobalFiModInstNr[2]) || (9786 == GlobalFiModInstNr[3]))));
	Tile mesh_13_0(
		.clock(clock),
		.io_in_a_0(r_416_0),
		.io_in_b_0(b_13_0),
		.io_in_d_0(b_1037_0),
		.io_in_control_0_dataflow(mesh_13_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2061_0),
		.io_in_last_0(r_3085_0),
		.io_in_valid_0(r_1037_0),
		.io_out_a_0(_mesh_13_0_io_out_a_0),
		.io_out_c_0(_mesh_13_0_io_out_c_0),
		.io_out_b_0(_mesh_13_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_0_io_out_id_0),
		.io_out_last_0(_mesh_13_0_io_out_last_0),
		.io_out_valid_0(_mesh_13_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9787 == GlobalFiModInstNr[0]) || (9787 == GlobalFiModInstNr[1]) || (9787 == GlobalFiModInstNr[2]) || (9787 == GlobalFiModInstNr[3]))));
	Tile mesh_13_1(
		.clock(clock),
		.io_in_a_0(r_417_0),
		.io_in_b_0(b_45_0),
		.io_in_d_0(b_1069_0),
		.io_in_control_0_dataflow(mesh_13_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2093_0),
		.io_in_last_0(r_3117_0),
		.io_in_valid_0(r_1069_0),
		.io_out_a_0(_mesh_13_1_io_out_a_0),
		.io_out_c_0(_mesh_13_1_io_out_c_0),
		.io_out_b_0(_mesh_13_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_1_io_out_id_0),
		.io_out_last_0(_mesh_13_1_io_out_last_0),
		.io_out_valid_0(_mesh_13_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9788 == GlobalFiModInstNr[0]) || (9788 == GlobalFiModInstNr[1]) || (9788 == GlobalFiModInstNr[2]) || (9788 == GlobalFiModInstNr[3]))));
	Tile mesh_13_2(
		.clock(clock),
		.io_in_a_0(r_418_0),
		.io_in_b_0(b_77_0),
		.io_in_d_0(b_1101_0),
		.io_in_control_0_dataflow(mesh_13_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2125_0),
		.io_in_last_0(r_3149_0),
		.io_in_valid_0(r_1101_0),
		.io_out_a_0(_mesh_13_2_io_out_a_0),
		.io_out_c_0(_mesh_13_2_io_out_c_0),
		.io_out_b_0(_mesh_13_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_2_io_out_id_0),
		.io_out_last_0(_mesh_13_2_io_out_last_0),
		.io_out_valid_0(_mesh_13_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9789 == GlobalFiModInstNr[0]) || (9789 == GlobalFiModInstNr[1]) || (9789 == GlobalFiModInstNr[2]) || (9789 == GlobalFiModInstNr[3]))));
	Tile mesh_13_3(
		.clock(clock),
		.io_in_a_0(r_419_0),
		.io_in_b_0(b_109_0),
		.io_in_d_0(b_1133_0),
		.io_in_control_0_dataflow(mesh_13_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2157_0),
		.io_in_last_0(r_3181_0),
		.io_in_valid_0(r_1133_0),
		.io_out_a_0(_mesh_13_3_io_out_a_0),
		.io_out_c_0(_mesh_13_3_io_out_c_0),
		.io_out_b_0(_mesh_13_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_3_io_out_id_0),
		.io_out_last_0(_mesh_13_3_io_out_last_0),
		.io_out_valid_0(_mesh_13_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9790 == GlobalFiModInstNr[0]) || (9790 == GlobalFiModInstNr[1]) || (9790 == GlobalFiModInstNr[2]) || (9790 == GlobalFiModInstNr[3]))));
	Tile mesh_13_4(
		.clock(clock),
		.io_in_a_0(r_420_0),
		.io_in_b_0(b_141_0),
		.io_in_d_0(b_1165_0),
		.io_in_control_0_dataflow(mesh_13_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2189_0),
		.io_in_last_0(r_3213_0),
		.io_in_valid_0(r_1165_0),
		.io_out_a_0(_mesh_13_4_io_out_a_0),
		.io_out_c_0(_mesh_13_4_io_out_c_0),
		.io_out_b_0(_mesh_13_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_4_io_out_id_0),
		.io_out_last_0(_mesh_13_4_io_out_last_0),
		.io_out_valid_0(_mesh_13_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9791 == GlobalFiModInstNr[0]) || (9791 == GlobalFiModInstNr[1]) || (9791 == GlobalFiModInstNr[2]) || (9791 == GlobalFiModInstNr[3]))));
	Tile mesh_13_5(
		.clock(clock),
		.io_in_a_0(r_421_0),
		.io_in_b_0(b_173_0),
		.io_in_d_0(b_1197_0),
		.io_in_control_0_dataflow(mesh_13_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2221_0),
		.io_in_last_0(r_3245_0),
		.io_in_valid_0(r_1197_0),
		.io_out_a_0(_mesh_13_5_io_out_a_0),
		.io_out_c_0(_mesh_13_5_io_out_c_0),
		.io_out_b_0(_mesh_13_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_5_io_out_id_0),
		.io_out_last_0(_mesh_13_5_io_out_last_0),
		.io_out_valid_0(_mesh_13_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9792 == GlobalFiModInstNr[0]) || (9792 == GlobalFiModInstNr[1]) || (9792 == GlobalFiModInstNr[2]) || (9792 == GlobalFiModInstNr[3]))));
	Tile mesh_13_6(
		.clock(clock),
		.io_in_a_0(r_422_0),
		.io_in_b_0(b_205_0),
		.io_in_d_0(b_1229_0),
		.io_in_control_0_dataflow(mesh_13_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2253_0),
		.io_in_last_0(r_3277_0),
		.io_in_valid_0(r_1229_0),
		.io_out_a_0(_mesh_13_6_io_out_a_0),
		.io_out_c_0(_mesh_13_6_io_out_c_0),
		.io_out_b_0(_mesh_13_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_6_io_out_id_0),
		.io_out_last_0(_mesh_13_6_io_out_last_0),
		.io_out_valid_0(_mesh_13_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9793 == GlobalFiModInstNr[0]) || (9793 == GlobalFiModInstNr[1]) || (9793 == GlobalFiModInstNr[2]) || (9793 == GlobalFiModInstNr[3]))));
	Tile mesh_13_7(
		.clock(clock),
		.io_in_a_0(r_423_0),
		.io_in_b_0(b_237_0),
		.io_in_d_0(b_1261_0),
		.io_in_control_0_dataflow(mesh_13_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2285_0),
		.io_in_last_0(r_3309_0),
		.io_in_valid_0(r_1261_0),
		.io_out_a_0(_mesh_13_7_io_out_a_0),
		.io_out_c_0(_mesh_13_7_io_out_c_0),
		.io_out_b_0(_mesh_13_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_7_io_out_id_0),
		.io_out_last_0(_mesh_13_7_io_out_last_0),
		.io_out_valid_0(_mesh_13_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9794 == GlobalFiModInstNr[0]) || (9794 == GlobalFiModInstNr[1]) || (9794 == GlobalFiModInstNr[2]) || (9794 == GlobalFiModInstNr[3]))));
	Tile mesh_13_8(
		.clock(clock),
		.io_in_a_0(r_424_0),
		.io_in_b_0(b_269_0),
		.io_in_d_0(b_1293_0),
		.io_in_control_0_dataflow(mesh_13_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2317_0),
		.io_in_last_0(r_3341_0),
		.io_in_valid_0(r_1293_0),
		.io_out_a_0(_mesh_13_8_io_out_a_0),
		.io_out_c_0(_mesh_13_8_io_out_c_0),
		.io_out_b_0(_mesh_13_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_8_io_out_id_0),
		.io_out_last_0(_mesh_13_8_io_out_last_0),
		.io_out_valid_0(_mesh_13_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9795 == GlobalFiModInstNr[0]) || (9795 == GlobalFiModInstNr[1]) || (9795 == GlobalFiModInstNr[2]) || (9795 == GlobalFiModInstNr[3]))));
	Tile mesh_13_9(
		.clock(clock),
		.io_in_a_0(r_425_0),
		.io_in_b_0(b_301_0),
		.io_in_d_0(b_1325_0),
		.io_in_control_0_dataflow(mesh_13_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2349_0),
		.io_in_last_0(r_3373_0),
		.io_in_valid_0(r_1325_0),
		.io_out_a_0(_mesh_13_9_io_out_a_0),
		.io_out_c_0(_mesh_13_9_io_out_c_0),
		.io_out_b_0(_mesh_13_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_9_io_out_id_0),
		.io_out_last_0(_mesh_13_9_io_out_last_0),
		.io_out_valid_0(_mesh_13_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9796 == GlobalFiModInstNr[0]) || (9796 == GlobalFiModInstNr[1]) || (9796 == GlobalFiModInstNr[2]) || (9796 == GlobalFiModInstNr[3]))));
	Tile mesh_13_10(
		.clock(clock),
		.io_in_a_0(r_426_0),
		.io_in_b_0(b_333_0),
		.io_in_d_0(b_1357_0),
		.io_in_control_0_dataflow(mesh_13_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2381_0),
		.io_in_last_0(r_3405_0),
		.io_in_valid_0(r_1357_0),
		.io_out_a_0(_mesh_13_10_io_out_a_0),
		.io_out_c_0(_mesh_13_10_io_out_c_0),
		.io_out_b_0(_mesh_13_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_10_io_out_id_0),
		.io_out_last_0(_mesh_13_10_io_out_last_0),
		.io_out_valid_0(_mesh_13_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9797 == GlobalFiModInstNr[0]) || (9797 == GlobalFiModInstNr[1]) || (9797 == GlobalFiModInstNr[2]) || (9797 == GlobalFiModInstNr[3]))));
	Tile mesh_13_11(
		.clock(clock),
		.io_in_a_0(r_427_0),
		.io_in_b_0(b_365_0),
		.io_in_d_0(b_1389_0),
		.io_in_control_0_dataflow(mesh_13_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2413_0),
		.io_in_last_0(r_3437_0),
		.io_in_valid_0(r_1389_0),
		.io_out_a_0(_mesh_13_11_io_out_a_0),
		.io_out_c_0(_mesh_13_11_io_out_c_0),
		.io_out_b_0(_mesh_13_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_11_io_out_id_0),
		.io_out_last_0(_mesh_13_11_io_out_last_0),
		.io_out_valid_0(_mesh_13_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9798 == GlobalFiModInstNr[0]) || (9798 == GlobalFiModInstNr[1]) || (9798 == GlobalFiModInstNr[2]) || (9798 == GlobalFiModInstNr[3]))));
	Tile mesh_13_12(
		.clock(clock),
		.io_in_a_0(r_428_0),
		.io_in_b_0(b_397_0),
		.io_in_d_0(b_1421_0),
		.io_in_control_0_dataflow(mesh_13_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2445_0),
		.io_in_last_0(r_3469_0),
		.io_in_valid_0(r_1421_0),
		.io_out_a_0(_mesh_13_12_io_out_a_0),
		.io_out_c_0(_mesh_13_12_io_out_c_0),
		.io_out_b_0(_mesh_13_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_12_io_out_id_0),
		.io_out_last_0(_mesh_13_12_io_out_last_0),
		.io_out_valid_0(_mesh_13_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9799 == GlobalFiModInstNr[0]) || (9799 == GlobalFiModInstNr[1]) || (9799 == GlobalFiModInstNr[2]) || (9799 == GlobalFiModInstNr[3]))));
	Tile mesh_13_13(
		.clock(clock),
		.io_in_a_0(r_429_0),
		.io_in_b_0(b_429_0),
		.io_in_d_0(b_1453_0),
		.io_in_control_0_dataflow(mesh_13_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2477_0),
		.io_in_last_0(r_3501_0),
		.io_in_valid_0(r_1453_0),
		.io_out_a_0(_mesh_13_13_io_out_a_0),
		.io_out_c_0(_mesh_13_13_io_out_c_0),
		.io_out_b_0(_mesh_13_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_13_io_out_id_0),
		.io_out_last_0(_mesh_13_13_io_out_last_0),
		.io_out_valid_0(_mesh_13_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9800 == GlobalFiModInstNr[0]) || (9800 == GlobalFiModInstNr[1]) || (9800 == GlobalFiModInstNr[2]) || (9800 == GlobalFiModInstNr[3]))));
	Tile mesh_13_14(
		.clock(clock),
		.io_in_a_0(r_430_0),
		.io_in_b_0(b_461_0),
		.io_in_d_0(b_1485_0),
		.io_in_control_0_dataflow(mesh_13_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2509_0),
		.io_in_last_0(r_3533_0),
		.io_in_valid_0(r_1485_0),
		.io_out_a_0(_mesh_13_14_io_out_a_0),
		.io_out_c_0(_mesh_13_14_io_out_c_0),
		.io_out_b_0(_mesh_13_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_14_io_out_id_0),
		.io_out_last_0(_mesh_13_14_io_out_last_0),
		.io_out_valid_0(_mesh_13_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9801 == GlobalFiModInstNr[0]) || (9801 == GlobalFiModInstNr[1]) || (9801 == GlobalFiModInstNr[2]) || (9801 == GlobalFiModInstNr[3]))));
	Tile mesh_13_15(
		.clock(clock),
		.io_in_a_0(r_431_0),
		.io_in_b_0(b_493_0),
		.io_in_d_0(b_1517_0),
		.io_in_control_0_dataflow(mesh_13_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2541_0),
		.io_in_last_0(r_3565_0),
		.io_in_valid_0(r_1517_0),
		.io_out_a_0(_mesh_13_15_io_out_a_0),
		.io_out_c_0(_mesh_13_15_io_out_c_0),
		.io_out_b_0(_mesh_13_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_15_io_out_id_0),
		.io_out_last_0(_mesh_13_15_io_out_last_0),
		.io_out_valid_0(_mesh_13_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9802 == GlobalFiModInstNr[0]) || (9802 == GlobalFiModInstNr[1]) || (9802 == GlobalFiModInstNr[2]) || (9802 == GlobalFiModInstNr[3]))));
	Tile mesh_13_16(
		.clock(clock),
		.io_in_a_0(r_432_0),
		.io_in_b_0(b_525_0),
		.io_in_d_0(b_1549_0),
		.io_in_control_0_dataflow(mesh_13_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2573_0),
		.io_in_last_0(r_3597_0),
		.io_in_valid_0(r_1549_0),
		.io_out_a_0(_mesh_13_16_io_out_a_0),
		.io_out_c_0(_mesh_13_16_io_out_c_0),
		.io_out_b_0(_mesh_13_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_16_io_out_id_0),
		.io_out_last_0(_mesh_13_16_io_out_last_0),
		.io_out_valid_0(_mesh_13_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9803 == GlobalFiModInstNr[0]) || (9803 == GlobalFiModInstNr[1]) || (9803 == GlobalFiModInstNr[2]) || (9803 == GlobalFiModInstNr[3]))));
	Tile mesh_13_17(
		.clock(clock),
		.io_in_a_0(r_433_0),
		.io_in_b_0(b_557_0),
		.io_in_d_0(b_1581_0),
		.io_in_control_0_dataflow(mesh_13_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2605_0),
		.io_in_last_0(r_3629_0),
		.io_in_valid_0(r_1581_0),
		.io_out_a_0(_mesh_13_17_io_out_a_0),
		.io_out_c_0(_mesh_13_17_io_out_c_0),
		.io_out_b_0(_mesh_13_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_17_io_out_id_0),
		.io_out_last_0(_mesh_13_17_io_out_last_0),
		.io_out_valid_0(_mesh_13_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9804 == GlobalFiModInstNr[0]) || (9804 == GlobalFiModInstNr[1]) || (9804 == GlobalFiModInstNr[2]) || (9804 == GlobalFiModInstNr[3]))));
	Tile mesh_13_18(
		.clock(clock),
		.io_in_a_0(r_434_0),
		.io_in_b_0(b_589_0),
		.io_in_d_0(b_1613_0),
		.io_in_control_0_dataflow(mesh_13_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2637_0),
		.io_in_last_0(r_3661_0),
		.io_in_valid_0(r_1613_0),
		.io_out_a_0(_mesh_13_18_io_out_a_0),
		.io_out_c_0(_mesh_13_18_io_out_c_0),
		.io_out_b_0(_mesh_13_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_18_io_out_id_0),
		.io_out_last_0(_mesh_13_18_io_out_last_0),
		.io_out_valid_0(_mesh_13_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9805 == GlobalFiModInstNr[0]) || (9805 == GlobalFiModInstNr[1]) || (9805 == GlobalFiModInstNr[2]) || (9805 == GlobalFiModInstNr[3]))));
	Tile mesh_13_19(
		.clock(clock),
		.io_in_a_0(r_435_0),
		.io_in_b_0(b_621_0),
		.io_in_d_0(b_1645_0),
		.io_in_control_0_dataflow(mesh_13_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2669_0),
		.io_in_last_0(r_3693_0),
		.io_in_valid_0(r_1645_0),
		.io_out_a_0(_mesh_13_19_io_out_a_0),
		.io_out_c_0(_mesh_13_19_io_out_c_0),
		.io_out_b_0(_mesh_13_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_19_io_out_id_0),
		.io_out_last_0(_mesh_13_19_io_out_last_0),
		.io_out_valid_0(_mesh_13_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9806 == GlobalFiModInstNr[0]) || (9806 == GlobalFiModInstNr[1]) || (9806 == GlobalFiModInstNr[2]) || (9806 == GlobalFiModInstNr[3]))));
	Tile mesh_13_20(
		.clock(clock),
		.io_in_a_0(r_436_0),
		.io_in_b_0(b_653_0),
		.io_in_d_0(b_1677_0),
		.io_in_control_0_dataflow(mesh_13_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2701_0),
		.io_in_last_0(r_3725_0),
		.io_in_valid_0(r_1677_0),
		.io_out_a_0(_mesh_13_20_io_out_a_0),
		.io_out_c_0(_mesh_13_20_io_out_c_0),
		.io_out_b_0(_mesh_13_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_20_io_out_id_0),
		.io_out_last_0(_mesh_13_20_io_out_last_0),
		.io_out_valid_0(_mesh_13_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9807 == GlobalFiModInstNr[0]) || (9807 == GlobalFiModInstNr[1]) || (9807 == GlobalFiModInstNr[2]) || (9807 == GlobalFiModInstNr[3]))));
	Tile mesh_13_21(
		.clock(clock),
		.io_in_a_0(r_437_0),
		.io_in_b_0(b_685_0),
		.io_in_d_0(b_1709_0),
		.io_in_control_0_dataflow(mesh_13_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2733_0),
		.io_in_last_0(r_3757_0),
		.io_in_valid_0(r_1709_0),
		.io_out_a_0(_mesh_13_21_io_out_a_0),
		.io_out_c_0(_mesh_13_21_io_out_c_0),
		.io_out_b_0(_mesh_13_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_21_io_out_id_0),
		.io_out_last_0(_mesh_13_21_io_out_last_0),
		.io_out_valid_0(_mesh_13_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9808 == GlobalFiModInstNr[0]) || (9808 == GlobalFiModInstNr[1]) || (9808 == GlobalFiModInstNr[2]) || (9808 == GlobalFiModInstNr[3]))));
	Tile mesh_13_22(
		.clock(clock),
		.io_in_a_0(r_438_0),
		.io_in_b_0(b_717_0),
		.io_in_d_0(b_1741_0),
		.io_in_control_0_dataflow(mesh_13_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2765_0),
		.io_in_last_0(r_3789_0),
		.io_in_valid_0(r_1741_0),
		.io_out_a_0(_mesh_13_22_io_out_a_0),
		.io_out_c_0(_mesh_13_22_io_out_c_0),
		.io_out_b_0(_mesh_13_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_22_io_out_id_0),
		.io_out_last_0(_mesh_13_22_io_out_last_0),
		.io_out_valid_0(_mesh_13_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9809 == GlobalFiModInstNr[0]) || (9809 == GlobalFiModInstNr[1]) || (9809 == GlobalFiModInstNr[2]) || (9809 == GlobalFiModInstNr[3]))));
	Tile mesh_13_23(
		.clock(clock),
		.io_in_a_0(r_439_0),
		.io_in_b_0(b_749_0),
		.io_in_d_0(b_1773_0),
		.io_in_control_0_dataflow(mesh_13_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2797_0),
		.io_in_last_0(r_3821_0),
		.io_in_valid_0(r_1773_0),
		.io_out_a_0(_mesh_13_23_io_out_a_0),
		.io_out_c_0(_mesh_13_23_io_out_c_0),
		.io_out_b_0(_mesh_13_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_23_io_out_id_0),
		.io_out_last_0(_mesh_13_23_io_out_last_0),
		.io_out_valid_0(_mesh_13_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9810 == GlobalFiModInstNr[0]) || (9810 == GlobalFiModInstNr[1]) || (9810 == GlobalFiModInstNr[2]) || (9810 == GlobalFiModInstNr[3]))));
	Tile mesh_13_24(
		.clock(clock),
		.io_in_a_0(r_440_0),
		.io_in_b_0(b_781_0),
		.io_in_d_0(b_1805_0),
		.io_in_control_0_dataflow(mesh_13_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2829_0),
		.io_in_last_0(r_3853_0),
		.io_in_valid_0(r_1805_0),
		.io_out_a_0(_mesh_13_24_io_out_a_0),
		.io_out_c_0(_mesh_13_24_io_out_c_0),
		.io_out_b_0(_mesh_13_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_24_io_out_id_0),
		.io_out_last_0(_mesh_13_24_io_out_last_0),
		.io_out_valid_0(_mesh_13_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9811 == GlobalFiModInstNr[0]) || (9811 == GlobalFiModInstNr[1]) || (9811 == GlobalFiModInstNr[2]) || (9811 == GlobalFiModInstNr[3]))));
	Tile mesh_13_25(
		.clock(clock),
		.io_in_a_0(r_441_0),
		.io_in_b_0(b_813_0),
		.io_in_d_0(b_1837_0),
		.io_in_control_0_dataflow(mesh_13_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2861_0),
		.io_in_last_0(r_3885_0),
		.io_in_valid_0(r_1837_0),
		.io_out_a_0(_mesh_13_25_io_out_a_0),
		.io_out_c_0(_mesh_13_25_io_out_c_0),
		.io_out_b_0(_mesh_13_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_25_io_out_id_0),
		.io_out_last_0(_mesh_13_25_io_out_last_0),
		.io_out_valid_0(_mesh_13_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9812 == GlobalFiModInstNr[0]) || (9812 == GlobalFiModInstNr[1]) || (9812 == GlobalFiModInstNr[2]) || (9812 == GlobalFiModInstNr[3]))));
	Tile mesh_13_26(
		.clock(clock),
		.io_in_a_0(r_442_0),
		.io_in_b_0(b_845_0),
		.io_in_d_0(b_1869_0),
		.io_in_control_0_dataflow(mesh_13_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2893_0),
		.io_in_last_0(r_3917_0),
		.io_in_valid_0(r_1869_0),
		.io_out_a_0(_mesh_13_26_io_out_a_0),
		.io_out_c_0(_mesh_13_26_io_out_c_0),
		.io_out_b_0(_mesh_13_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_26_io_out_id_0),
		.io_out_last_0(_mesh_13_26_io_out_last_0),
		.io_out_valid_0(_mesh_13_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9813 == GlobalFiModInstNr[0]) || (9813 == GlobalFiModInstNr[1]) || (9813 == GlobalFiModInstNr[2]) || (9813 == GlobalFiModInstNr[3]))));
	Tile mesh_13_27(
		.clock(clock),
		.io_in_a_0(r_443_0),
		.io_in_b_0(b_877_0),
		.io_in_d_0(b_1901_0),
		.io_in_control_0_dataflow(mesh_13_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2925_0),
		.io_in_last_0(r_3949_0),
		.io_in_valid_0(r_1901_0),
		.io_out_a_0(_mesh_13_27_io_out_a_0),
		.io_out_c_0(_mesh_13_27_io_out_c_0),
		.io_out_b_0(_mesh_13_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_27_io_out_id_0),
		.io_out_last_0(_mesh_13_27_io_out_last_0),
		.io_out_valid_0(_mesh_13_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9814 == GlobalFiModInstNr[0]) || (9814 == GlobalFiModInstNr[1]) || (9814 == GlobalFiModInstNr[2]) || (9814 == GlobalFiModInstNr[3]))));
	Tile mesh_13_28(
		.clock(clock),
		.io_in_a_0(r_444_0),
		.io_in_b_0(b_909_0),
		.io_in_d_0(b_1933_0),
		.io_in_control_0_dataflow(mesh_13_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2957_0),
		.io_in_last_0(r_3981_0),
		.io_in_valid_0(r_1933_0),
		.io_out_a_0(_mesh_13_28_io_out_a_0),
		.io_out_c_0(_mesh_13_28_io_out_c_0),
		.io_out_b_0(_mesh_13_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_28_io_out_id_0),
		.io_out_last_0(_mesh_13_28_io_out_last_0),
		.io_out_valid_0(_mesh_13_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9815 == GlobalFiModInstNr[0]) || (9815 == GlobalFiModInstNr[1]) || (9815 == GlobalFiModInstNr[2]) || (9815 == GlobalFiModInstNr[3]))));
	Tile mesh_13_29(
		.clock(clock),
		.io_in_a_0(r_445_0),
		.io_in_b_0(b_941_0),
		.io_in_d_0(b_1965_0),
		.io_in_control_0_dataflow(mesh_13_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2989_0),
		.io_in_last_0(r_4013_0),
		.io_in_valid_0(r_1965_0),
		.io_out_a_0(_mesh_13_29_io_out_a_0),
		.io_out_c_0(_mesh_13_29_io_out_c_0),
		.io_out_b_0(_mesh_13_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_29_io_out_id_0),
		.io_out_last_0(_mesh_13_29_io_out_last_0),
		.io_out_valid_0(_mesh_13_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9816 == GlobalFiModInstNr[0]) || (9816 == GlobalFiModInstNr[1]) || (9816 == GlobalFiModInstNr[2]) || (9816 == GlobalFiModInstNr[3]))));
	Tile mesh_13_30(
		.clock(clock),
		.io_in_a_0(r_446_0),
		.io_in_b_0(b_973_0),
		.io_in_d_0(b_1997_0),
		.io_in_control_0_dataflow(mesh_13_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3021_0),
		.io_in_last_0(r_4045_0),
		.io_in_valid_0(r_1997_0),
		.io_out_a_0(_mesh_13_30_io_out_a_0),
		.io_out_c_0(_mesh_13_30_io_out_c_0),
		.io_out_b_0(_mesh_13_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_30_io_out_id_0),
		.io_out_last_0(_mesh_13_30_io_out_last_0),
		.io_out_valid_0(_mesh_13_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9817 == GlobalFiModInstNr[0]) || (9817 == GlobalFiModInstNr[1]) || (9817 == GlobalFiModInstNr[2]) || (9817 == GlobalFiModInstNr[3]))));
	Tile mesh_13_31(
		.clock(clock),
		.io_in_a_0(r_447_0),
		.io_in_b_0(b_1005_0),
		.io_in_d_0(b_2029_0),
		.io_in_control_0_dataflow(mesh_13_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_13_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_13_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3053_0),
		.io_in_last_0(r_4077_0),
		.io_in_valid_0(r_2029_0),
		.io_out_a_0(_mesh_13_31_io_out_a_0),
		.io_out_c_0(_mesh_13_31_io_out_c_0),
		.io_out_b_0(_mesh_13_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_13_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_13_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_13_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_13_31_io_out_id_0),
		.io_out_last_0(_mesh_13_31_io_out_last_0),
		.io_out_valid_0(_mesh_13_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9818 == GlobalFiModInstNr[0]) || (9818 == GlobalFiModInstNr[1]) || (9818 == GlobalFiModInstNr[2]) || (9818 == GlobalFiModInstNr[3]))));
	Tile mesh_14_0(
		.clock(clock),
		.io_in_a_0(r_448_0),
		.io_in_b_0(b_14_0),
		.io_in_d_0(b_1038_0),
		.io_in_control_0_dataflow(mesh_14_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2062_0),
		.io_in_last_0(r_3086_0),
		.io_in_valid_0(r_1038_0),
		.io_out_a_0(_mesh_14_0_io_out_a_0),
		.io_out_c_0(_mesh_14_0_io_out_c_0),
		.io_out_b_0(_mesh_14_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_0_io_out_id_0),
		.io_out_last_0(_mesh_14_0_io_out_last_0),
		.io_out_valid_0(_mesh_14_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9819 == GlobalFiModInstNr[0]) || (9819 == GlobalFiModInstNr[1]) || (9819 == GlobalFiModInstNr[2]) || (9819 == GlobalFiModInstNr[3]))));
	Tile mesh_14_1(
		.clock(clock),
		.io_in_a_0(r_449_0),
		.io_in_b_0(b_46_0),
		.io_in_d_0(b_1070_0),
		.io_in_control_0_dataflow(mesh_14_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2094_0),
		.io_in_last_0(r_3118_0),
		.io_in_valid_0(r_1070_0),
		.io_out_a_0(_mesh_14_1_io_out_a_0),
		.io_out_c_0(_mesh_14_1_io_out_c_0),
		.io_out_b_0(_mesh_14_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_1_io_out_id_0),
		.io_out_last_0(_mesh_14_1_io_out_last_0),
		.io_out_valid_0(_mesh_14_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9820 == GlobalFiModInstNr[0]) || (9820 == GlobalFiModInstNr[1]) || (9820 == GlobalFiModInstNr[2]) || (9820 == GlobalFiModInstNr[3]))));
	Tile mesh_14_2(
		.clock(clock),
		.io_in_a_0(r_450_0),
		.io_in_b_0(b_78_0),
		.io_in_d_0(b_1102_0),
		.io_in_control_0_dataflow(mesh_14_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2126_0),
		.io_in_last_0(r_3150_0),
		.io_in_valid_0(r_1102_0),
		.io_out_a_0(_mesh_14_2_io_out_a_0),
		.io_out_c_0(_mesh_14_2_io_out_c_0),
		.io_out_b_0(_mesh_14_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_2_io_out_id_0),
		.io_out_last_0(_mesh_14_2_io_out_last_0),
		.io_out_valid_0(_mesh_14_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9821 == GlobalFiModInstNr[0]) || (9821 == GlobalFiModInstNr[1]) || (9821 == GlobalFiModInstNr[2]) || (9821 == GlobalFiModInstNr[3]))));
	Tile mesh_14_3(
		.clock(clock),
		.io_in_a_0(r_451_0),
		.io_in_b_0(b_110_0),
		.io_in_d_0(b_1134_0),
		.io_in_control_0_dataflow(mesh_14_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2158_0),
		.io_in_last_0(r_3182_0),
		.io_in_valid_0(r_1134_0),
		.io_out_a_0(_mesh_14_3_io_out_a_0),
		.io_out_c_0(_mesh_14_3_io_out_c_0),
		.io_out_b_0(_mesh_14_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_3_io_out_id_0),
		.io_out_last_0(_mesh_14_3_io_out_last_0),
		.io_out_valid_0(_mesh_14_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9822 == GlobalFiModInstNr[0]) || (9822 == GlobalFiModInstNr[1]) || (9822 == GlobalFiModInstNr[2]) || (9822 == GlobalFiModInstNr[3]))));
	Tile mesh_14_4(
		.clock(clock),
		.io_in_a_0(r_452_0),
		.io_in_b_0(b_142_0),
		.io_in_d_0(b_1166_0),
		.io_in_control_0_dataflow(mesh_14_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2190_0),
		.io_in_last_0(r_3214_0),
		.io_in_valid_0(r_1166_0),
		.io_out_a_0(_mesh_14_4_io_out_a_0),
		.io_out_c_0(_mesh_14_4_io_out_c_0),
		.io_out_b_0(_mesh_14_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_4_io_out_id_0),
		.io_out_last_0(_mesh_14_4_io_out_last_0),
		.io_out_valid_0(_mesh_14_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9823 == GlobalFiModInstNr[0]) || (9823 == GlobalFiModInstNr[1]) || (9823 == GlobalFiModInstNr[2]) || (9823 == GlobalFiModInstNr[3]))));
	Tile mesh_14_5(
		.clock(clock),
		.io_in_a_0(r_453_0),
		.io_in_b_0(b_174_0),
		.io_in_d_0(b_1198_0),
		.io_in_control_0_dataflow(mesh_14_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2222_0),
		.io_in_last_0(r_3246_0),
		.io_in_valid_0(r_1198_0),
		.io_out_a_0(_mesh_14_5_io_out_a_0),
		.io_out_c_0(_mesh_14_5_io_out_c_0),
		.io_out_b_0(_mesh_14_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_5_io_out_id_0),
		.io_out_last_0(_mesh_14_5_io_out_last_0),
		.io_out_valid_0(_mesh_14_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9824 == GlobalFiModInstNr[0]) || (9824 == GlobalFiModInstNr[1]) || (9824 == GlobalFiModInstNr[2]) || (9824 == GlobalFiModInstNr[3]))));
	Tile mesh_14_6(
		.clock(clock),
		.io_in_a_0(r_454_0),
		.io_in_b_0(b_206_0),
		.io_in_d_0(b_1230_0),
		.io_in_control_0_dataflow(mesh_14_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2254_0),
		.io_in_last_0(r_3278_0),
		.io_in_valid_0(r_1230_0),
		.io_out_a_0(_mesh_14_6_io_out_a_0),
		.io_out_c_0(_mesh_14_6_io_out_c_0),
		.io_out_b_0(_mesh_14_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_6_io_out_id_0),
		.io_out_last_0(_mesh_14_6_io_out_last_0),
		.io_out_valid_0(_mesh_14_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9825 == GlobalFiModInstNr[0]) || (9825 == GlobalFiModInstNr[1]) || (9825 == GlobalFiModInstNr[2]) || (9825 == GlobalFiModInstNr[3]))));
	Tile mesh_14_7(
		.clock(clock),
		.io_in_a_0(r_455_0),
		.io_in_b_0(b_238_0),
		.io_in_d_0(b_1262_0),
		.io_in_control_0_dataflow(mesh_14_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2286_0),
		.io_in_last_0(r_3310_0),
		.io_in_valid_0(r_1262_0),
		.io_out_a_0(_mesh_14_7_io_out_a_0),
		.io_out_c_0(_mesh_14_7_io_out_c_0),
		.io_out_b_0(_mesh_14_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_7_io_out_id_0),
		.io_out_last_0(_mesh_14_7_io_out_last_0),
		.io_out_valid_0(_mesh_14_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9826 == GlobalFiModInstNr[0]) || (9826 == GlobalFiModInstNr[1]) || (9826 == GlobalFiModInstNr[2]) || (9826 == GlobalFiModInstNr[3]))));
	Tile mesh_14_8(
		.clock(clock),
		.io_in_a_0(r_456_0),
		.io_in_b_0(b_270_0),
		.io_in_d_0(b_1294_0),
		.io_in_control_0_dataflow(mesh_14_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2318_0),
		.io_in_last_0(r_3342_0),
		.io_in_valid_0(r_1294_0),
		.io_out_a_0(_mesh_14_8_io_out_a_0),
		.io_out_c_0(_mesh_14_8_io_out_c_0),
		.io_out_b_0(_mesh_14_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_8_io_out_id_0),
		.io_out_last_0(_mesh_14_8_io_out_last_0),
		.io_out_valid_0(_mesh_14_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9827 == GlobalFiModInstNr[0]) || (9827 == GlobalFiModInstNr[1]) || (9827 == GlobalFiModInstNr[2]) || (9827 == GlobalFiModInstNr[3]))));
	Tile mesh_14_9(
		.clock(clock),
		.io_in_a_0(r_457_0),
		.io_in_b_0(b_302_0),
		.io_in_d_0(b_1326_0),
		.io_in_control_0_dataflow(mesh_14_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2350_0),
		.io_in_last_0(r_3374_0),
		.io_in_valid_0(r_1326_0),
		.io_out_a_0(_mesh_14_9_io_out_a_0),
		.io_out_c_0(_mesh_14_9_io_out_c_0),
		.io_out_b_0(_mesh_14_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_9_io_out_id_0),
		.io_out_last_0(_mesh_14_9_io_out_last_0),
		.io_out_valid_0(_mesh_14_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9828 == GlobalFiModInstNr[0]) || (9828 == GlobalFiModInstNr[1]) || (9828 == GlobalFiModInstNr[2]) || (9828 == GlobalFiModInstNr[3]))));
	Tile mesh_14_10(
		.clock(clock),
		.io_in_a_0(r_458_0),
		.io_in_b_0(b_334_0),
		.io_in_d_0(b_1358_0),
		.io_in_control_0_dataflow(mesh_14_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2382_0),
		.io_in_last_0(r_3406_0),
		.io_in_valid_0(r_1358_0),
		.io_out_a_0(_mesh_14_10_io_out_a_0),
		.io_out_c_0(_mesh_14_10_io_out_c_0),
		.io_out_b_0(_mesh_14_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_10_io_out_id_0),
		.io_out_last_0(_mesh_14_10_io_out_last_0),
		.io_out_valid_0(_mesh_14_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9829 == GlobalFiModInstNr[0]) || (9829 == GlobalFiModInstNr[1]) || (9829 == GlobalFiModInstNr[2]) || (9829 == GlobalFiModInstNr[3]))));
	Tile mesh_14_11(
		.clock(clock),
		.io_in_a_0(r_459_0),
		.io_in_b_0(b_366_0),
		.io_in_d_0(b_1390_0),
		.io_in_control_0_dataflow(mesh_14_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2414_0),
		.io_in_last_0(r_3438_0),
		.io_in_valid_0(r_1390_0),
		.io_out_a_0(_mesh_14_11_io_out_a_0),
		.io_out_c_0(_mesh_14_11_io_out_c_0),
		.io_out_b_0(_mesh_14_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_11_io_out_id_0),
		.io_out_last_0(_mesh_14_11_io_out_last_0),
		.io_out_valid_0(_mesh_14_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9830 == GlobalFiModInstNr[0]) || (9830 == GlobalFiModInstNr[1]) || (9830 == GlobalFiModInstNr[2]) || (9830 == GlobalFiModInstNr[3]))));
	Tile mesh_14_12(
		.clock(clock),
		.io_in_a_0(r_460_0),
		.io_in_b_0(b_398_0),
		.io_in_d_0(b_1422_0),
		.io_in_control_0_dataflow(mesh_14_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2446_0),
		.io_in_last_0(r_3470_0),
		.io_in_valid_0(r_1422_0),
		.io_out_a_0(_mesh_14_12_io_out_a_0),
		.io_out_c_0(_mesh_14_12_io_out_c_0),
		.io_out_b_0(_mesh_14_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_12_io_out_id_0),
		.io_out_last_0(_mesh_14_12_io_out_last_0),
		.io_out_valid_0(_mesh_14_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9831 == GlobalFiModInstNr[0]) || (9831 == GlobalFiModInstNr[1]) || (9831 == GlobalFiModInstNr[2]) || (9831 == GlobalFiModInstNr[3]))));
	Tile mesh_14_13(
		.clock(clock),
		.io_in_a_0(r_461_0),
		.io_in_b_0(b_430_0),
		.io_in_d_0(b_1454_0),
		.io_in_control_0_dataflow(mesh_14_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2478_0),
		.io_in_last_0(r_3502_0),
		.io_in_valid_0(r_1454_0),
		.io_out_a_0(_mesh_14_13_io_out_a_0),
		.io_out_c_0(_mesh_14_13_io_out_c_0),
		.io_out_b_0(_mesh_14_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_13_io_out_id_0),
		.io_out_last_0(_mesh_14_13_io_out_last_0),
		.io_out_valid_0(_mesh_14_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9832 == GlobalFiModInstNr[0]) || (9832 == GlobalFiModInstNr[1]) || (9832 == GlobalFiModInstNr[2]) || (9832 == GlobalFiModInstNr[3]))));
	Tile mesh_14_14(
		.clock(clock),
		.io_in_a_0(r_462_0),
		.io_in_b_0(b_462_0),
		.io_in_d_0(b_1486_0),
		.io_in_control_0_dataflow(mesh_14_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2510_0),
		.io_in_last_0(r_3534_0),
		.io_in_valid_0(r_1486_0),
		.io_out_a_0(_mesh_14_14_io_out_a_0),
		.io_out_c_0(_mesh_14_14_io_out_c_0),
		.io_out_b_0(_mesh_14_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_14_io_out_id_0),
		.io_out_last_0(_mesh_14_14_io_out_last_0),
		.io_out_valid_0(_mesh_14_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9833 == GlobalFiModInstNr[0]) || (9833 == GlobalFiModInstNr[1]) || (9833 == GlobalFiModInstNr[2]) || (9833 == GlobalFiModInstNr[3]))));
	Tile mesh_14_15(
		.clock(clock),
		.io_in_a_0(r_463_0),
		.io_in_b_0(b_494_0),
		.io_in_d_0(b_1518_0),
		.io_in_control_0_dataflow(mesh_14_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2542_0),
		.io_in_last_0(r_3566_0),
		.io_in_valid_0(r_1518_0),
		.io_out_a_0(_mesh_14_15_io_out_a_0),
		.io_out_c_0(_mesh_14_15_io_out_c_0),
		.io_out_b_0(_mesh_14_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_15_io_out_id_0),
		.io_out_last_0(_mesh_14_15_io_out_last_0),
		.io_out_valid_0(_mesh_14_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9834 == GlobalFiModInstNr[0]) || (9834 == GlobalFiModInstNr[1]) || (9834 == GlobalFiModInstNr[2]) || (9834 == GlobalFiModInstNr[3]))));
	Tile mesh_14_16(
		.clock(clock),
		.io_in_a_0(r_464_0),
		.io_in_b_0(b_526_0),
		.io_in_d_0(b_1550_0),
		.io_in_control_0_dataflow(mesh_14_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2574_0),
		.io_in_last_0(r_3598_0),
		.io_in_valid_0(r_1550_0),
		.io_out_a_0(_mesh_14_16_io_out_a_0),
		.io_out_c_0(_mesh_14_16_io_out_c_0),
		.io_out_b_0(_mesh_14_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_16_io_out_id_0),
		.io_out_last_0(_mesh_14_16_io_out_last_0),
		.io_out_valid_0(_mesh_14_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9835 == GlobalFiModInstNr[0]) || (9835 == GlobalFiModInstNr[1]) || (9835 == GlobalFiModInstNr[2]) || (9835 == GlobalFiModInstNr[3]))));
	Tile mesh_14_17(
		.clock(clock),
		.io_in_a_0(r_465_0),
		.io_in_b_0(b_558_0),
		.io_in_d_0(b_1582_0),
		.io_in_control_0_dataflow(mesh_14_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2606_0),
		.io_in_last_0(r_3630_0),
		.io_in_valid_0(r_1582_0),
		.io_out_a_0(_mesh_14_17_io_out_a_0),
		.io_out_c_0(_mesh_14_17_io_out_c_0),
		.io_out_b_0(_mesh_14_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_17_io_out_id_0),
		.io_out_last_0(_mesh_14_17_io_out_last_0),
		.io_out_valid_0(_mesh_14_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9836 == GlobalFiModInstNr[0]) || (9836 == GlobalFiModInstNr[1]) || (9836 == GlobalFiModInstNr[2]) || (9836 == GlobalFiModInstNr[3]))));
	Tile mesh_14_18(
		.clock(clock),
		.io_in_a_0(r_466_0),
		.io_in_b_0(b_590_0),
		.io_in_d_0(b_1614_0),
		.io_in_control_0_dataflow(mesh_14_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2638_0),
		.io_in_last_0(r_3662_0),
		.io_in_valid_0(r_1614_0),
		.io_out_a_0(_mesh_14_18_io_out_a_0),
		.io_out_c_0(_mesh_14_18_io_out_c_0),
		.io_out_b_0(_mesh_14_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_18_io_out_id_0),
		.io_out_last_0(_mesh_14_18_io_out_last_0),
		.io_out_valid_0(_mesh_14_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9837 == GlobalFiModInstNr[0]) || (9837 == GlobalFiModInstNr[1]) || (9837 == GlobalFiModInstNr[2]) || (9837 == GlobalFiModInstNr[3]))));
	Tile mesh_14_19(
		.clock(clock),
		.io_in_a_0(r_467_0),
		.io_in_b_0(b_622_0),
		.io_in_d_0(b_1646_0),
		.io_in_control_0_dataflow(mesh_14_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2670_0),
		.io_in_last_0(r_3694_0),
		.io_in_valid_0(r_1646_0),
		.io_out_a_0(_mesh_14_19_io_out_a_0),
		.io_out_c_0(_mesh_14_19_io_out_c_0),
		.io_out_b_0(_mesh_14_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_19_io_out_id_0),
		.io_out_last_0(_mesh_14_19_io_out_last_0),
		.io_out_valid_0(_mesh_14_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9838 == GlobalFiModInstNr[0]) || (9838 == GlobalFiModInstNr[1]) || (9838 == GlobalFiModInstNr[2]) || (9838 == GlobalFiModInstNr[3]))));
	Tile mesh_14_20(
		.clock(clock),
		.io_in_a_0(r_468_0),
		.io_in_b_0(b_654_0),
		.io_in_d_0(b_1678_0),
		.io_in_control_0_dataflow(mesh_14_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2702_0),
		.io_in_last_0(r_3726_0),
		.io_in_valid_0(r_1678_0),
		.io_out_a_0(_mesh_14_20_io_out_a_0),
		.io_out_c_0(_mesh_14_20_io_out_c_0),
		.io_out_b_0(_mesh_14_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_20_io_out_id_0),
		.io_out_last_0(_mesh_14_20_io_out_last_0),
		.io_out_valid_0(_mesh_14_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9839 == GlobalFiModInstNr[0]) || (9839 == GlobalFiModInstNr[1]) || (9839 == GlobalFiModInstNr[2]) || (9839 == GlobalFiModInstNr[3]))));
	Tile mesh_14_21(
		.clock(clock),
		.io_in_a_0(r_469_0),
		.io_in_b_0(b_686_0),
		.io_in_d_0(b_1710_0),
		.io_in_control_0_dataflow(mesh_14_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2734_0),
		.io_in_last_0(r_3758_0),
		.io_in_valid_0(r_1710_0),
		.io_out_a_0(_mesh_14_21_io_out_a_0),
		.io_out_c_0(_mesh_14_21_io_out_c_0),
		.io_out_b_0(_mesh_14_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_21_io_out_id_0),
		.io_out_last_0(_mesh_14_21_io_out_last_0),
		.io_out_valid_0(_mesh_14_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9840 == GlobalFiModInstNr[0]) || (9840 == GlobalFiModInstNr[1]) || (9840 == GlobalFiModInstNr[2]) || (9840 == GlobalFiModInstNr[3]))));
	Tile mesh_14_22(
		.clock(clock),
		.io_in_a_0(r_470_0),
		.io_in_b_0(b_718_0),
		.io_in_d_0(b_1742_0),
		.io_in_control_0_dataflow(mesh_14_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2766_0),
		.io_in_last_0(r_3790_0),
		.io_in_valid_0(r_1742_0),
		.io_out_a_0(_mesh_14_22_io_out_a_0),
		.io_out_c_0(_mesh_14_22_io_out_c_0),
		.io_out_b_0(_mesh_14_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_22_io_out_id_0),
		.io_out_last_0(_mesh_14_22_io_out_last_0),
		.io_out_valid_0(_mesh_14_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9841 == GlobalFiModInstNr[0]) || (9841 == GlobalFiModInstNr[1]) || (9841 == GlobalFiModInstNr[2]) || (9841 == GlobalFiModInstNr[3]))));
	Tile mesh_14_23(
		.clock(clock),
		.io_in_a_0(r_471_0),
		.io_in_b_0(b_750_0),
		.io_in_d_0(b_1774_0),
		.io_in_control_0_dataflow(mesh_14_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2798_0),
		.io_in_last_0(r_3822_0),
		.io_in_valid_0(r_1774_0),
		.io_out_a_0(_mesh_14_23_io_out_a_0),
		.io_out_c_0(_mesh_14_23_io_out_c_0),
		.io_out_b_0(_mesh_14_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_23_io_out_id_0),
		.io_out_last_0(_mesh_14_23_io_out_last_0),
		.io_out_valid_0(_mesh_14_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9842 == GlobalFiModInstNr[0]) || (9842 == GlobalFiModInstNr[1]) || (9842 == GlobalFiModInstNr[2]) || (9842 == GlobalFiModInstNr[3]))));
	Tile mesh_14_24(
		.clock(clock),
		.io_in_a_0(r_472_0),
		.io_in_b_0(b_782_0),
		.io_in_d_0(b_1806_0),
		.io_in_control_0_dataflow(mesh_14_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2830_0),
		.io_in_last_0(r_3854_0),
		.io_in_valid_0(r_1806_0),
		.io_out_a_0(_mesh_14_24_io_out_a_0),
		.io_out_c_0(_mesh_14_24_io_out_c_0),
		.io_out_b_0(_mesh_14_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_24_io_out_id_0),
		.io_out_last_0(_mesh_14_24_io_out_last_0),
		.io_out_valid_0(_mesh_14_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9843 == GlobalFiModInstNr[0]) || (9843 == GlobalFiModInstNr[1]) || (9843 == GlobalFiModInstNr[2]) || (9843 == GlobalFiModInstNr[3]))));
	Tile mesh_14_25(
		.clock(clock),
		.io_in_a_0(r_473_0),
		.io_in_b_0(b_814_0),
		.io_in_d_0(b_1838_0),
		.io_in_control_0_dataflow(mesh_14_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2862_0),
		.io_in_last_0(r_3886_0),
		.io_in_valid_0(r_1838_0),
		.io_out_a_0(_mesh_14_25_io_out_a_0),
		.io_out_c_0(_mesh_14_25_io_out_c_0),
		.io_out_b_0(_mesh_14_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_25_io_out_id_0),
		.io_out_last_0(_mesh_14_25_io_out_last_0),
		.io_out_valid_0(_mesh_14_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9844 == GlobalFiModInstNr[0]) || (9844 == GlobalFiModInstNr[1]) || (9844 == GlobalFiModInstNr[2]) || (9844 == GlobalFiModInstNr[3]))));
	Tile mesh_14_26(
		.clock(clock),
		.io_in_a_0(r_474_0),
		.io_in_b_0(b_846_0),
		.io_in_d_0(b_1870_0),
		.io_in_control_0_dataflow(mesh_14_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2894_0),
		.io_in_last_0(r_3918_0),
		.io_in_valid_0(r_1870_0),
		.io_out_a_0(_mesh_14_26_io_out_a_0),
		.io_out_c_0(_mesh_14_26_io_out_c_0),
		.io_out_b_0(_mesh_14_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_26_io_out_id_0),
		.io_out_last_0(_mesh_14_26_io_out_last_0),
		.io_out_valid_0(_mesh_14_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9845 == GlobalFiModInstNr[0]) || (9845 == GlobalFiModInstNr[1]) || (9845 == GlobalFiModInstNr[2]) || (9845 == GlobalFiModInstNr[3]))));
	Tile mesh_14_27(
		.clock(clock),
		.io_in_a_0(r_475_0),
		.io_in_b_0(b_878_0),
		.io_in_d_0(b_1902_0),
		.io_in_control_0_dataflow(mesh_14_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2926_0),
		.io_in_last_0(r_3950_0),
		.io_in_valid_0(r_1902_0),
		.io_out_a_0(_mesh_14_27_io_out_a_0),
		.io_out_c_0(_mesh_14_27_io_out_c_0),
		.io_out_b_0(_mesh_14_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_27_io_out_id_0),
		.io_out_last_0(_mesh_14_27_io_out_last_0),
		.io_out_valid_0(_mesh_14_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9846 == GlobalFiModInstNr[0]) || (9846 == GlobalFiModInstNr[1]) || (9846 == GlobalFiModInstNr[2]) || (9846 == GlobalFiModInstNr[3]))));
	Tile mesh_14_28(
		.clock(clock),
		.io_in_a_0(r_476_0),
		.io_in_b_0(b_910_0),
		.io_in_d_0(b_1934_0),
		.io_in_control_0_dataflow(mesh_14_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2958_0),
		.io_in_last_0(r_3982_0),
		.io_in_valid_0(r_1934_0),
		.io_out_a_0(_mesh_14_28_io_out_a_0),
		.io_out_c_0(_mesh_14_28_io_out_c_0),
		.io_out_b_0(_mesh_14_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_28_io_out_id_0),
		.io_out_last_0(_mesh_14_28_io_out_last_0),
		.io_out_valid_0(_mesh_14_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9847 == GlobalFiModInstNr[0]) || (9847 == GlobalFiModInstNr[1]) || (9847 == GlobalFiModInstNr[2]) || (9847 == GlobalFiModInstNr[3]))));
	Tile mesh_14_29(
		.clock(clock),
		.io_in_a_0(r_477_0),
		.io_in_b_0(b_942_0),
		.io_in_d_0(b_1966_0),
		.io_in_control_0_dataflow(mesh_14_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2990_0),
		.io_in_last_0(r_4014_0),
		.io_in_valid_0(r_1966_0),
		.io_out_a_0(_mesh_14_29_io_out_a_0),
		.io_out_c_0(_mesh_14_29_io_out_c_0),
		.io_out_b_0(_mesh_14_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_29_io_out_id_0),
		.io_out_last_0(_mesh_14_29_io_out_last_0),
		.io_out_valid_0(_mesh_14_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9848 == GlobalFiModInstNr[0]) || (9848 == GlobalFiModInstNr[1]) || (9848 == GlobalFiModInstNr[2]) || (9848 == GlobalFiModInstNr[3]))));
	Tile mesh_14_30(
		.clock(clock),
		.io_in_a_0(r_478_0),
		.io_in_b_0(b_974_0),
		.io_in_d_0(b_1998_0),
		.io_in_control_0_dataflow(mesh_14_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3022_0),
		.io_in_last_0(r_4046_0),
		.io_in_valid_0(r_1998_0),
		.io_out_a_0(_mesh_14_30_io_out_a_0),
		.io_out_c_0(_mesh_14_30_io_out_c_0),
		.io_out_b_0(_mesh_14_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_30_io_out_id_0),
		.io_out_last_0(_mesh_14_30_io_out_last_0),
		.io_out_valid_0(_mesh_14_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9849 == GlobalFiModInstNr[0]) || (9849 == GlobalFiModInstNr[1]) || (9849 == GlobalFiModInstNr[2]) || (9849 == GlobalFiModInstNr[3]))));
	Tile mesh_14_31(
		.clock(clock),
		.io_in_a_0(r_479_0),
		.io_in_b_0(b_1006_0),
		.io_in_d_0(b_2030_0),
		.io_in_control_0_dataflow(mesh_14_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_14_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_14_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3054_0),
		.io_in_last_0(r_4078_0),
		.io_in_valid_0(r_2030_0),
		.io_out_a_0(_mesh_14_31_io_out_a_0),
		.io_out_c_0(_mesh_14_31_io_out_c_0),
		.io_out_b_0(_mesh_14_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_14_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_14_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_14_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_14_31_io_out_id_0),
		.io_out_last_0(_mesh_14_31_io_out_last_0),
		.io_out_valid_0(_mesh_14_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9850 == GlobalFiModInstNr[0]) || (9850 == GlobalFiModInstNr[1]) || (9850 == GlobalFiModInstNr[2]) || (9850 == GlobalFiModInstNr[3]))));
	Tile mesh_15_0(
		.clock(clock),
		.io_in_a_0(r_480_0),
		.io_in_b_0(b_15_0),
		.io_in_d_0(b_1039_0),
		.io_in_control_0_dataflow(mesh_15_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2063_0),
		.io_in_last_0(r_3087_0),
		.io_in_valid_0(r_1039_0),
		.io_out_a_0(_mesh_15_0_io_out_a_0),
		.io_out_c_0(_mesh_15_0_io_out_c_0),
		.io_out_b_0(_mesh_15_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_0_io_out_id_0),
		.io_out_last_0(_mesh_15_0_io_out_last_0),
		.io_out_valid_0(_mesh_15_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9851 == GlobalFiModInstNr[0]) || (9851 == GlobalFiModInstNr[1]) || (9851 == GlobalFiModInstNr[2]) || (9851 == GlobalFiModInstNr[3]))));
	Tile mesh_15_1(
		.clock(clock),
		.io_in_a_0(r_481_0),
		.io_in_b_0(b_47_0),
		.io_in_d_0(b_1071_0),
		.io_in_control_0_dataflow(mesh_15_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2095_0),
		.io_in_last_0(r_3119_0),
		.io_in_valid_0(r_1071_0),
		.io_out_a_0(_mesh_15_1_io_out_a_0),
		.io_out_c_0(_mesh_15_1_io_out_c_0),
		.io_out_b_0(_mesh_15_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_1_io_out_id_0),
		.io_out_last_0(_mesh_15_1_io_out_last_0),
		.io_out_valid_0(_mesh_15_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9852 == GlobalFiModInstNr[0]) || (9852 == GlobalFiModInstNr[1]) || (9852 == GlobalFiModInstNr[2]) || (9852 == GlobalFiModInstNr[3]))));
	Tile mesh_15_2(
		.clock(clock),
		.io_in_a_0(r_482_0),
		.io_in_b_0(b_79_0),
		.io_in_d_0(b_1103_0),
		.io_in_control_0_dataflow(mesh_15_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2127_0),
		.io_in_last_0(r_3151_0),
		.io_in_valid_0(r_1103_0),
		.io_out_a_0(_mesh_15_2_io_out_a_0),
		.io_out_c_0(_mesh_15_2_io_out_c_0),
		.io_out_b_0(_mesh_15_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_2_io_out_id_0),
		.io_out_last_0(_mesh_15_2_io_out_last_0),
		.io_out_valid_0(_mesh_15_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9853 == GlobalFiModInstNr[0]) || (9853 == GlobalFiModInstNr[1]) || (9853 == GlobalFiModInstNr[2]) || (9853 == GlobalFiModInstNr[3]))));
	Tile mesh_15_3(
		.clock(clock),
		.io_in_a_0(r_483_0),
		.io_in_b_0(b_111_0),
		.io_in_d_0(b_1135_0),
		.io_in_control_0_dataflow(mesh_15_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2159_0),
		.io_in_last_0(r_3183_0),
		.io_in_valid_0(r_1135_0),
		.io_out_a_0(_mesh_15_3_io_out_a_0),
		.io_out_c_0(_mesh_15_3_io_out_c_0),
		.io_out_b_0(_mesh_15_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_3_io_out_id_0),
		.io_out_last_0(_mesh_15_3_io_out_last_0),
		.io_out_valid_0(_mesh_15_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9854 == GlobalFiModInstNr[0]) || (9854 == GlobalFiModInstNr[1]) || (9854 == GlobalFiModInstNr[2]) || (9854 == GlobalFiModInstNr[3]))));
	Tile mesh_15_4(
		.clock(clock),
		.io_in_a_0(r_484_0),
		.io_in_b_0(b_143_0),
		.io_in_d_0(b_1167_0),
		.io_in_control_0_dataflow(mesh_15_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2191_0),
		.io_in_last_0(r_3215_0),
		.io_in_valid_0(r_1167_0),
		.io_out_a_0(_mesh_15_4_io_out_a_0),
		.io_out_c_0(_mesh_15_4_io_out_c_0),
		.io_out_b_0(_mesh_15_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_4_io_out_id_0),
		.io_out_last_0(_mesh_15_4_io_out_last_0),
		.io_out_valid_0(_mesh_15_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9855 == GlobalFiModInstNr[0]) || (9855 == GlobalFiModInstNr[1]) || (9855 == GlobalFiModInstNr[2]) || (9855 == GlobalFiModInstNr[3]))));
	Tile mesh_15_5(
		.clock(clock),
		.io_in_a_0(r_485_0),
		.io_in_b_0(b_175_0),
		.io_in_d_0(b_1199_0),
		.io_in_control_0_dataflow(mesh_15_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2223_0),
		.io_in_last_0(r_3247_0),
		.io_in_valid_0(r_1199_0),
		.io_out_a_0(_mesh_15_5_io_out_a_0),
		.io_out_c_0(_mesh_15_5_io_out_c_0),
		.io_out_b_0(_mesh_15_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_5_io_out_id_0),
		.io_out_last_0(_mesh_15_5_io_out_last_0),
		.io_out_valid_0(_mesh_15_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9856 == GlobalFiModInstNr[0]) || (9856 == GlobalFiModInstNr[1]) || (9856 == GlobalFiModInstNr[2]) || (9856 == GlobalFiModInstNr[3]))));
	Tile mesh_15_6(
		.clock(clock),
		.io_in_a_0(r_486_0),
		.io_in_b_0(b_207_0),
		.io_in_d_0(b_1231_0),
		.io_in_control_0_dataflow(mesh_15_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2255_0),
		.io_in_last_0(r_3279_0),
		.io_in_valid_0(r_1231_0),
		.io_out_a_0(_mesh_15_6_io_out_a_0),
		.io_out_c_0(_mesh_15_6_io_out_c_0),
		.io_out_b_0(_mesh_15_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_6_io_out_id_0),
		.io_out_last_0(_mesh_15_6_io_out_last_0),
		.io_out_valid_0(_mesh_15_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9857 == GlobalFiModInstNr[0]) || (9857 == GlobalFiModInstNr[1]) || (9857 == GlobalFiModInstNr[2]) || (9857 == GlobalFiModInstNr[3]))));
	Tile mesh_15_7(
		.clock(clock),
		.io_in_a_0(r_487_0),
		.io_in_b_0(b_239_0),
		.io_in_d_0(b_1263_0),
		.io_in_control_0_dataflow(mesh_15_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2287_0),
		.io_in_last_0(r_3311_0),
		.io_in_valid_0(r_1263_0),
		.io_out_a_0(_mesh_15_7_io_out_a_0),
		.io_out_c_0(_mesh_15_7_io_out_c_0),
		.io_out_b_0(_mesh_15_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_7_io_out_id_0),
		.io_out_last_0(_mesh_15_7_io_out_last_0),
		.io_out_valid_0(_mesh_15_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9858 == GlobalFiModInstNr[0]) || (9858 == GlobalFiModInstNr[1]) || (9858 == GlobalFiModInstNr[2]) || (9858 == GlobalFiModInstNr[3]))));
	Tile mesh_15_8(
		.clock(clock),
		.io_in_a_0(r_488_0),
		.io_in_b_0(b_271_0),
		.io_in_d_0(b_1295_0),
		.io_in_control_0_dataflow(mesh_15_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2319_0),
		.io_in_last_0(r_3343_0),
		.io_in_valid_0(r_1295_0),
		.io_out_a_0(_mesh_15_8_io_out_a_0),
		.io_out_c_0(_mesh_15_8_io_out_c_0),
		.io_out_b_0(_mesh_15_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_8_io_out_id_0),
		.io_out_last_0(_mesh_15_8_io_out_last_0),
		.io_out_valid_0(_mesh_15_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9859 == GlobalFiModInstNr[0]) || (9859 == GlobalFiModInstNr[1]) || (9859 == GlobalFiModInstNr[2]) || (9859 == GlobalFiModInstNr[3]))));
	Tile mesh_15_9(
		.clock(clock),
		.io_in_a_0(r_489_0),
		.io_in_b_0(b_303_0),
		.io_in_d_0(b_1327_0),
		.io_in_control_0_dataflow(mesh_15_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2351_0),
		.io_in_last_0(r_3375_0),
		.io_in_valid_0(r_1327_0),
		.io_out_a_0(_mesh_15_9_io_out_a_0),
		.io_out_c_0(_mesh_15_9_io_out_c_0),
		.io_out_b_0(_mesh_15_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_9_io_out_id_0),
		.io_out_last_0(_mesh_15_9_io_out_last_0),
		.io_out_valid_0(_mesh_15_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9860 == GlobalFiModInstNr[0]) || (9860 == GlobalFiModInstNr[1]) || (9860 == GlobalFiModInstNr[2]) || (9860 == GlobalFiModInstNr[3]))));
	Tile mesh_15_10(
		.clock(clock),
		.io_in_a_0(r_490_0),
		.io_in_b_0(b_335_0),
		.io_in_d_0(b_1359_0),
		.io_in_control_0_dataflow(mesh_15_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2383_0),
		.io_in_last_0(r_3407_0),
		.io_in_valid_0(r_1359_0),
		.io_out_a_0(_mesh_15_10_io_out_a_0),
		.io_out_c_0(_mesh_15_10_io_out_c_0),
		.io_out_b_0(_mesh_15_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_10_io_out_id_0),
		.io_out_last_0(_mesh_15_10_io_out_last_0),
		.io_out_valid_0(_mesh_15_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9861 == GlobalFiModInstNr[0]) || (9861 == GlobalFiModInstNr[1]) || (9861 == GlobalFiModInstNr[2]) || (9861 == GlobalFiModInstNr[3]))));
	Tile mesh_15_11(
		.clock(clock),
		.io_in_a_0(r_491_0),
		.io_in_b_0(b_367_0),
		.io_in_d_0(b_1391_0),
		.io_in_control_0_dataflow(mesh_15_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2415_0),
		.io_in_last_0(r_3439_0),
		.io_in_valid_0(r_1391_0),
		.io_out_a_0(_mesh_15_11_io_out_a_0),
		.io_out_c_0(_mesh_15_11_io_out_c_0),
		.io_out_b_0(_mesh_15_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_11_io_out_id_0),
		.io_out_last_0(_mesh_15_11_io_out_last_0),
		.io_out_valid_0(_mesh_15_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9862 == GlobalFiModInstNr[0]) || (9862 == GlobalFiModInstNr[1]) || (9862 == GlobalFiModInstNr[2]) || (9862 == GlobalFiModInstNr[3]))));
	Tile mesh_15_12(
		.clock(clock),
		.io_in_a_0(r_492_0),
		.io_in_b_0(b_399_0),
		.io_in_d_0(b_1423_0),
		.io_in_control_0_dataflow(mesh_15_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2447_0),
		.io_in_last_0(r_3471_0),
		.io_in_valid_0(r_1423_0),
		.io_out_a_0(_mesh_15_12_io_out_a_0),
		.io_out_c_0(_mesh_15_12_io_out_c_0),
		.io_out_b_0(_mesh_15_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_12_io_out_id_0),
		.io_out_last_0(_mesh_15_12_io_out_last_0),
		.io_out_valid_0(_mesh_15_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9863 == GlobalFiModInstNr[0]) || (9863 == GlobalFiModInstNr[1]) || (9863 == GlobalFiModInstNr[2]) || (9863 == GlobalFiModInstNr[3]))));
	Tile mesh_15_13(
		.clock(clock),
		.io_in_a_0(r_493_0),
		.io_in_b_0(b_431_0),
		.io_in_d_0(b_1455_0),
		.io_in_control_0_dataflow(mesh_15_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2479_0),
		.io_in_last_0(r_3503_0),
		.io_in_valid_0(r_1455_0),
		.io_out_a_0(_mesh_15_13_io_out_a_0),
		.io_out_c_0(_mesh_15_13_io_out_c_0),
		.io_out_b_0(_mesh_15_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_13_io_out_id_0),
		.io_out_last_0(_mesh_15_13_io_out_last_0),
		.io_out_valid_0(_mesh_15_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9864 == GlobalFiModInstNr[0]) || (9864 == GlobalFiModInstNr[1]) || (9864 == GlobalFiModInstNr[2]) || (9864 == GlobalFiModInstNr[3]))));
	Tile mesh_15_14(
		.clock(clock),
		.io_in_a_0(r_494_0),
		.io_in_b_0(b_463_0),
		.io_in_d_0(b_1487_0),
		.io_in_control_0_dataflow(mesh_15_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2511_0),
		.io_in_last_0(r_3535_0),
		.io_in_valid_0(r_1487_0),
		.io_out_a_0(_mesh_15_14_io_out_a_0),
		.io_out_c_0(_mesh_15_14_io_out_c_0),
		.io_out_b_0(_mesh_15_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_14_io_out_id_0),
		.io_out_last_0(_mesh_15_14_io_out_last_0),
		.io_out_valid_0(_mesh_15_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9865 == GlobalFiModInstNr[0]) || (9865 == GlobalFiModInstNr[1]) || (9865 == GlobalFiModInstNr[2]) || (9865 == GlobalFiModInstNr[3]))));
	Tile mesh_15_15(
		.clock(clock),
		.io_in_a_0(r_495_0),
		.io_in_b_0(b_495_0),
		.io_in_d_0(b_1519_0),
		.io_in_control_0_dataflow(mesh_15_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2543_0),
		.io_in_last_0(r_3567_0),
		.io_in_valid_0(r_1519_0),
		.io_out_a_0(_mesh_15_15_io_out_a_0),
		.io_out_c_0(_mesh_15_15_io_out_c_0),
		.io_out_b_0(_mesh_15_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_15_io_out_id_0),
		.io_out_last_0(_mesh_15_15_io_out_last_0),
		.io_out_valid_0(_mesh_15_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9866 == GlobalFiModInstNr[0]) || (9866 == GlobalFiModInstNr[1]) || (9866 == GlobalFiModInstNr[2]) || (9866 == GlobalFiModInstNr[3]))));
	Tile mesh_15_16(
		.clock(clock),
		.io_in_a_0(r_496_0),
		.io_in_b_0(b_527_0),
		.io_in_d_0(b_1551_0),
		.io_in_control_0_dataflow(mesh_15_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2575_0),
		.io_in_last_0(r_3599_0),
		.io_in_valid_0(r_1551_0),
		.io_out_a_0(_mesh_15_16_io_out_a_0),
		.io_out_c_0(_mesh_15_16_io_out_c_0),
		.io_out_b_0(_mesh_15_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_16_io_out_id_0),
		.io_out_last_0(_mesh_15_16_io_out_last_0),
		.io_out_valid_0(_mesh_15_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9867 == GlobalFiModInstNr[0]) || (9867 == GlobalFiModInstNr[1]) || (9867 == GlobalFiModInstNr[2]) || (9867 == GlobalFiModInstNr[3]))));
	Tile mesh_15_17(
		.clock(clock),
		.io_in_a_0(r_497_0),
		.io_in_b_0(b_559_0),
		.io_in_d_0(b_1583_0),
		.io_in_control_0_dataflow(mesh_15_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2607_0),
		.io_in_last_0(r_3631_0),
		.io_in_valid_0(r_1583_0),
		.io_out_a_0(_mesh_15_17_io_out_a_0),
		.io_out_c_0(_mesh_15_17_io_out_c_0),
		.io_out_b_0(_mesh_15_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_17_io_out_id_0),
		.io_out_last_0(_mesh_15_17_io_out_last_0),
		.io_out_valid_0(_mesh_15_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9868 == GlobalFiModInstNr[0]) || (9868 == GlobalFiModInstNr[1]) || (9868 == GlobalFiModInstNr[2]) || (9868 == GlobalFiModInstNr[3]))));
	Tile mesh_15_18(
		.clock(clock),
		.io_in_a_0(r_498_0),
		.io_in_b_0(b_591_0),
		.io_in_d_0(b_1615_0),
		.io_in_control_0_dataflow(mesh_15_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2639_0),
		.io_in_last_0(r_3663_0),
		.io_in_valid_0(r_1615_0),
		.io_out_a_0(_mesh_15_18_io_out_a_0),
		.io_out_c_0(_mesh_15_18_io_out_c_0),
		.io_out_b_0(_mesh_15_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_18_io_out_id_0),
		.io_out_last_0(_mesh_15_18_io_out_last_0),
		.io_out_valid_0(_mesh_15_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9869 == GlobalFiModInstNr[0]) || (9869 == GlobalFiModInstNr[1]) || (9869 == GlobalFiModInstNr[2]) || (9869 == GlobalFiModInstNr[3]))));
	Tile mesh_15_19(
		.clock(clock),
		.io_in_a_0(r_499_0),
		.io_in_b_0(b_623_0),
		.io_in_d_0(b_1647_0),
		.io_in_control_0_dataflow(mesh_15_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2671_0),
		.io_in_last_0(r_3695_0),
		.io_in_valid_0(r_1647_0),
		.io_out_a_0(_mesh_15_19_io_out_a_0),
		.io_out_c_0(_mesh_15_19_io_out_c_0),
		.io_out_b_0(_mesh_15_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_19_io_out_id_0),
		.io_out_last_0(_mesh_15_19_io_out_last_0),
		.io_out_valid_0(_mesh_15_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9870 == GlobalFiModInstNr[0]) || (9870 == GlobalFiModInstNr[1]) || (9870 == GlobalFiModInstNr[2]) || (9870 == GlobalFiModInstNr[3]))));
	Tile mesh_15_20(
		.clock(clock),
		.io_in_a_0(r_500_0),
		.io_in_b_0(b_655_0),
		.io_in_d_0(b_1679_0),
		.io_in_control_0_dataflow(mesh_15_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2703_0),
		.io_in_last_0(r_3727_0),
		.io_in_valid_0(r_1679_0),
		.io_out_a_0(_mesh_15_20_io_out_a_0),
		.io_out_c_0(_mesh_15_20_io_out_c_0),
		.io_out_b_0(_mesh_15_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_20_io_out_id_0),
		.io_out_last_0(_mesh_15_20_io_out_last_0),
		.io_out_valid_0(_mesh_15_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9871 == GlobalFiModInstNr[0]) || (9871 == GlobalFiModInstNr[1]) || (9871 == GlobalFiModInstNr[2]) || (9871 == GlobalFiModInstNr[3]))));
	Tile mesh_15_21(
		.clock(clock),
		.io_in_a_0(r_501_0),
		.io_in_b_0(b_687_0),
		.io_in_d_0(b_1711_0),
		.io_in_control_0_dataflow(mesh_15_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2735_0),
		.io_in_last_0(r_3759_0),
		.io_in_valid_0(r_1711_0),
		.io_out_a_0(_mesh_15_21_io_out_a_0),
		.io_out_c_0(_mesh_15_21_io_out_c_0),
		.io_out_b_0(_mesh_15_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_21_io_out_id_0),
		.io_out_last_0(_mesh_15_21_io_out_last_0),
		.io_out_valid_0(_mesh_15_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9872 == GlobalFiModInstNr[0]) || (9872 == GlobalFiModInstNr[1]) || (9872 == GlobalFiModInstNr[2]) || (9872 == GlobalFiModInstNr[3]))));
	Tile mesh_15_22(
		.clock(clock),
		.io_in_a_0(r_502_0),
		.io_in_b_0(b_719_0),
		.io_in_d_0(b_1743_0),
		.io_in_control_0_dataflow(mesh_15_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2767_0),
		.io_in_last_0(r_3791_0),
		.io_in_valid_0(r_1743_0),
		.io_out_a_0(_mesh_15_22_io_out_a_0),
		.io_out_c_0(_mesh_15_22_io_out_c_0),
		.io_out_b_0(_mesh_15_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_22_io_out_id_0),
		.io_out_last_0(_mesh_15_22_io_out_last_0),
		.io_out_valid_0(_mesh_15_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9873 == GlobalFiModInstNr[0]) || (9873 == GlobalFiModInstNr[1]) || (9873 == GlobalFiModInstNr[2]) || (9873 == GlobalFiModInstNr[3]))));
	Tile mesh_15_23(
		.clock(clock),
		.io_in_a_0(r_503_0),
		.io_in_b_0(b_751_0),
		.io_in_d_0(b_1775_0),
		.io_in_control_0_dataflow(mesh_15_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2799_0),
		.io_in_last_0(r_3823_0),
		.io_in_valid_0(r_1775_0),
		.io_out_a_0(_mesh_15_23_io_out_a_0),
		.io_out_c_0(_mesh_15_23_io_out_c_0),
		.io_out_b_0(_mesh_15_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_23_io_out_id_0),
		.io_out_last_0(_mesh_15_23_io_out_last_0),
		.io_out_valid_0(_mesh_15_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9874 == GlobalFiModInstNr[0]) || (9874 == GlobalFiModInstNr[1]) || (9874 == GlobalFiModInstNr[2]) || (9874 == GlobalFiModInstNr[3]))));
	Tile mesh_15_24(
		.clock(clock),
		.io_in_a_0(r_504_0),
		.io_in_b_0(b_783_0),
		.io_in_d_0(b_1807_0),
		.io_in_control_0_dataflow(mesh_15_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2831_0),
		.io_in_last_0(r_3855_0),
		.io_in_valid_0(r_1807_0),
		.io_out_a_0(_mesh_15_24_io_out_a_0),
		.io_out_c_0(_mesh_15_24_io_out_c_0),
		.io_out_b_0(_mesh_15_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_24_io_out_id_0),
		.io_out_last_0(_mesh_15_24_io_out_last_0),
		.io_out_valid_0(_mesh_15_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9875 == GlobalFiModInstNr[0]) || (9875 == GlobalFiModInstNr[1]) || (9875 == GlobalFiModInstNr[2]) || (9875 == GlobalFiModInstNr[3]))));
	Tile mesh_15_25(
		.clock(clock),
		.io_in_a_0(r_505_0),
		.io_in_b_0(b_815_0),
		.io_in_d_0(b_1839_0),
		.io_in_control_0_dataflow(mesh_15_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2863_0),
		.io_in_last_0(r_3887_0),
		.io_in_valid_0(r_1839_0),
		.io_out_a_0(_mesh_15_25_io_out_a_0),
		.io_out_c_0(_mesh_15_25_io_out_c_0),
		.io_out_b_0(_mesh_15_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_25_io_out_id_0),
		.io_out_last_0(_mesh_15_25_io_out_last_0),
		.io_out_valid_0(_mesh_15_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9876 == GlobalFiModInstNr[0]) || (9876 == GlobalFiModInstNr[1]) || (9876 == GlobalFiModInstNr[2]) || (9876 == GlobalFiModInstNr[3]))));
	Tile mesh_15_26(
		.clock(clock),
		.io_in_a_0(r_506_0),
		.io_in_b_0(b_847_0),
		.io_in_d_0(b_1871_0),
		.io_in_control_0_dataflow(mesh_15_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2895_0),
		.io_in_last_0(r_3919_0),
		.io_in_valid_0(r_1871_0),
		.io_out_a_0(_mesh_15_26_io_out_a_0),
		.io_out_c_0(_mesh_15_26_io_out_c_0),
		.io_out_b_0(_mesh_15_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_26_io_out_id_0),
		.io_out_last_0(_mesh_15_26_io_out_last_0),
		.io_out_valid_0(_mesh_15_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9877 == GlobalFiModInstNr[0]) || (9877 == GlobalFiModInstNr[1]) || (9877 == GlobalFiModInstNr[2]) || (9877 == GlobalFiModInstNr[3]))));
	Tile mesh_15_27(
		.clock(clock),
		.io_in_a_0(r_507_0),
		.io_in_b_0(b_879_0),
		.io_in_d_0(b_1903_0),
		.io_in_control_0_dataflow(mesh_15_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2927_0),
		.io_in_last_0(r_3951_0),
		.io_in_valid_0(r_1903_0),
		.io_out_a_0(_mesh_15_27_io_out_a_0),
		.io_out_c_0(_mesh_15_27_io_out_c_0),
		.io_out_b_0(_mesh_15_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_27_io_out_id_0),
		.io_out_last_0(_mesh_15_27_io_out_last_0),
		.io_out_valid_0(_mesh_15_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9878 == GlobalFiModInstNr[0]) || (9878 == GlobalFiModInstNr[1]) || (9878 == GlobalFiModInstNr[2]) || (9878 == GlobalFiModInstNr[3]))));
	Tile mesh_15_28(
		.clock(clock),
		.io_in_a_0(r_508_0),
		.io_in_b_0(b_911_0),
		.io_in_d_0(b_1935_0),
		.io_in_control_0_dataflow(mesh_15_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2959_0),
		.io_in_last_0(r_3983_0),
		.io_in_valid_0(r_1935_0),
		.io_out_a_0(_mesh_15_28_io_out_a_0),
		.io_out_c_0(_mesh_15_28_io_out_c_0),
		.io_out_b_0(_mesh_15_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_28_io_out_id_0),
		.io_out_last_0(_mesh_15_28_io_out_last_0),
		.io_out_valid_0(_mesh_15_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9879 == GlobalFiModInstNr[0]) || (9879 == GlobalFiModInstNr[1]) || (9879 == GlobalFiModInstNr[2]) || (9879 == GlobalFiModInstNr[3]))));
	Tile mesh_15_29(
		.clock(clock),
		.io_in_a_0(r_509_0),
		.io_in_b_0(b_943_0),
		.io_in_d_0(b_1967_0),
		.io_in_control_0_dataflow(mesh_15_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2991_0),
		.io_in_last_0(r_4015_0),
		.io_in_valid_0(r_1967_0),
		.io_out_a_0(_mesh_15_29_io_out_a_0),
		.io_out_c_0(_mesh_15_29_io_out_c_0),
		.io_out_b_0(_mesh_15_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_29_io_out_id_0),
		.io_out_last_0(_mesh_15_29_io_out_last_0),
		.io_out_valid_0(_mesh_15_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9880 == GlobalFiModInstNr[0]) || (9880 == GlobalFiModInstNr[1]) || (9880 == GlobalFiModInstNr[2]) || (9880 == GlobalFiModInstNr[3]))));
	Tile mesh_15_30(
		.clock(clock),
		.io_in_a_0(r_510_0),
		.io_in_b_0(b_975_0),
		.io_in_d_0(b_1999_0),
		.io_in_control_0_dataflow(mesh_15_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3023_0),
		.io_in_last_0(r_4047_0),
		.io_in_valid_0(r_1999_0),
		.io_out_a_0(_mesh_15_30_io_out_a_0),
		.io_out_c_0(_mesh_15_30_io_out_c_0),
		.io_out_b_0(_mesh_15_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_30_io_out_id_0),
		.io_out_last_0(_mesh_15_30_io_out_last_0),
		.io_out_valid_0(_mesh_15_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9881 == GlobalFiModInstNr[0]) || (9881 == GlobalFiModInstNr[1]) || (9881 == GlobalFiModInstNr[2]) || (9881 == GlobalFiModInstNr[3]))));
	Tile mesh_15_31(
		.clock(clock),
		.io_in_a_0(r_511_0),
		.io_in_b_0(b_1007_0),
		.io_in_d_0(b_2031_0),
		.io_in_control_0_dataflow(mesh_15_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_15_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_15_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3055_0),
		.io_in_last_0(r_4079_0),
		.io_in_valid_0(r_2031_0),
		.io_out_a_0(_mesh_15_31_io_out_a_0),
		.io_out_c_0(_mesh_15_31_io_out_c_0),
		.io_out_b_0(_mesh_15_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_15_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_15_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_15_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_15_31_io_out_id_0),
		.io_out_last_0(_mesh_15_31_io_out_last_0),
		.io_out_valid_0(_mesh_15_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9882 == GlobalFiModInstNr[0]) || (9882 == GlobalFiModInstNr[1]) || (9882 == GlobalFiModInstNr[2]) || (9882 == GlobalFiModInstNr[3]))));
	Tile mesh_16_0(
		.clock(clock),
		.io_in_a_0(r_512_0),
		.io_in_b_0(b_16_0),
		.io_in_d_0(b_1040_0),
		.io_in_control_0_dataflow(mesh_16_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2064_0),
		.io_in_last_0(r_3088_0),
		.io_in_valid_0(r_1040_0),
		.io_out_a_0(_mesh_16_0_io_out_a_0),
		.io_out_c_0(_mesh_16_0_io_out_c_0),
		.io_out_b_0(_mesh_16_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_0_io_out_id_0),
		.io_out_last_0(_mesh_16_0_io_out_last_0),
		.io_out_valid_0(_mesh_16_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9883 == GlobalFiModInstNr[0]) || (9883 == GlobalFiModInstNr[1]) || (9883 == GlobalFiModInstNr[2]) || (9883 == GlobalFiModInstNr[3]))));
	Tile mesh_16_1(
		.clock(clock),
		.io_in_a_0(r_513_0),
		.io_in_b_0(b_48_0),
		.io_in_d_0(b_1072_0),
		.io_in_control_0_dataflow(mesh_16_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2096_0),
		.io_in_last_0(r_3120_0),
		.io_in_valid_0(r_1072_0),
		.io_out_a_0(_mesh_16_1_io_out_a_0),
		.io_out_c_0(_mesh_16_1_io_out_c_0),
		.io_out_b_0(_mesh_16_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_1_io_out_id_0),
		.io_out_last_0(_mesh_16_1_io_out_last_0),
		.io_out_valid_0(_mesh_16_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9884 == GlobalFiModInstNr[0]) || (9884 == GlobalFiModInstNr[1]) || (9884 == GlobalFiModInstNr[2]) || (9884 == GlobalFiModInstNr[3]))));
	Tile mesh_16_2(
		.clock(clock),
		.io_in_a_0(r_514_0),
		.io_in_b_0(b_80_0),
		.io_in_d_0(b_1104_0),
		.io_in_control_0_dataflow(mesh_16_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2128_0),
		.io_in_last_0(r_3152_0),
		.io_in_valid_0(r_1104_0),
		.io_out_a_0(_mesh_16_2_io_out_a_0),
		.io_out_c_0(_mesh_16_2_io_out_c_0),
		.io_out_b_0(_mesh_16_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_2_io_out_id_0),
		.io_out_last_0(_mesh_16_2_io_out_last_0),
		.io_out_valid_0(_mesh_16_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9885 == GlobalFiModInstNr[0]) || (9885 == GlobalFiModInstNr[1]) || (9885 == GlobalFiModInstNr[2]) || (9885 == GlobalFiModInstNr[3]))));
	Tile mesh_16_3(
		.clock(clock),
		.io_in_a_0(r_515_0),
		.io_in_b_0(b_112_0),
		.io_in_d_0(b_1136_0),
		.io_in_control_0_dataflow(mesh_16_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2160_0),
		.io_in_last_0(r_3184_0),
		.io_in_valid_0(r_1136_0),
		.io_out_a_0(_mesh_16_3_io_out_a_0),
		.io_out_c_0(_mesh_16_3_io_out_c_0),
		.io_out_b_0(_mesh_16_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_3_io_out_id_0),
		.io_out_last_0(_mesh_16_3_io_out_last_0),
		.io_out_valid_0(_mesh_16_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9886 == GlobalFiModInstNr[0]) || (9886 == GlobalFiModInstNr[1]) || (9886 == GlobalFiModInstNr[2]) || (9886 == GlobalFiModInstNr[3]))));
	Tile mesh_16_4(
		.clock(clock),
		.io_in_a_0(r_516_0),
		.io_in_b_0(b_144_0),
		.io_in_d_0(b_1168_0),
		.io_in_control_0_dataflow(mesh_16_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2192_0),
		.io_in_last_0(r_3216_0),
		.io_in_valid_0(r_1168_0),
		.io_out_a_0(_mesh_16_4_io_out_a_0),
		.io_out_c_0(_mesh_16_4_io_out_c_0),
		.io_out_b_0(_mesh_16_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_4_io_out_id_0),
		.io_out_last_0(_mesh_16_4_io_out_last_0),
		.io_out_valid_0(_mesh_16_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9887 == GlobalFiModInstNr[0]) || (9887 == GlobalFiModInstNr[1]) || (9887 == GlobalFiModInstNr[2]) || (9887 == GlobalFiModInstNr[3]))));
	Tile mesh_16_5(
		.clock(clock),
		.io_in_a_0(r_517_0),
		.io_in_b_0(b_176_0),
		.io_in_d_0(b_1200_0),
		.io_in_control_0_dataflow(mesh_16_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2224_0),
		.io_in_last_0(r_3248_0),
		.io_in_valid_0(r_1200_0),
		.io_out_a_0(_mesh_16_5_io_out_a_0),
		.io_out_c_0(_mesh_16_5_io_out_c_0),
		.io_out_b_0(_mesh_16_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_5_io_out_id_0),
		.io_out_last_0(_mesh_16_5_io_out_last_0),
		.io_out_valid_0(_mesh_16_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9888 == GlobalFiModInstNr[0]) || (9888 == GlobalFiModInstNr[1]) || (9888 == GlobalFiModInstNr[2]) || (9888 == GlobalFiModInstNr[3]))));
	Tile mesh_16_6(
		.clock(clock),
		.io_in_a_0(r_518_0),
		.io_in_b_0(b_208_0),
		.io_in_d_0(b_1232_0),
		.io_in_control_0_dataflow(mesh_16_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2256_0),
		.io_in_last_0(r_3280_0),
		.io_in_valid_0(r_1232_0),
		.io_out_a_0(_mesh_16_6_io_out_a_0),
		.io_out_c_0(_mesh_16_6_io_out_c_0),
		.io_out_b_0(_mesh_16_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_6_io_out_id_0),
		.io_out_last_0(_mesh_16_6_io_out_last_0),
		.io_out_valid_0(_mesh_16_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9889 == GlobalFiModInstNr[0]) || (9889 == GlobalFiModInstNr[1]) || (9889 == GlobalFiModInstNr[2]) || (9889 == GlobalFiModInstNr[3]))));
	Tile mesh_16_7(
		.clock(clock),
		.io_in_a_0(r_519_0),
		.io_in_b_0(b_240_0),
		.io_in_d_0(b_1264_0),
		.io_in_control_0_dataflow(mesh_16_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2288_0),
		.io_in_last_0(r_3312_0),
		.io_in_valid_0(r_1264_0),
		.io_out_a_0(_mesh_16_7_io_out_a_0),
		.io_out_c_0(_mesh_16_7_io_out_c_0),
		.io_out_b_0(_mesh_16_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_7_io_out_id_0),
		.io_out_last_0(_mesh_16_7_io_out_last_0),
		.io_out_valid_0(_mesh_16_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9890 == GlobalFiModInstNr[0]) || (9890 == GlobalFiModInstNr[1]) || (9890 == GlobalFiModInstNr[2]) || (9890 == GlobalFiModInstNr[3]))));
	Tile mesh_16_8(
		.clock(clock),
		.io_in_a_0(r_520_0),
		.io_in_b_0(b_272_0),
		.io_in_d_0(b_1296_0),
		.io_in_control_0_dataflow(mesh_16_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2320_0),
		.io_in_last_0(r_3344_0),
		.io_in_valid_0(r_1296_0),
		.io_out_a_0(_mesh_16_8_io_out_a_0),
		.io_out_c_0(_mesh_16_8_io_out_c_0),
		.io_out_b_0(_mesh_16_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_8_io_out_id_0),
		.io_out_last_0(_mesh_16_8_io_out_last_0),
		.io_out_valid_0(_mesh_16_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9891 == GlobalFiModInstNr[0]) || (9891 == GlobalFiModInstNr[1]) || (9891 == GlobalFiModInstNr[2]) || (9891 == GlobalFiModInstNr[3]))));
	Tile mesh_16_9(
		.clock(clock),
		.io_in_a_0(r_521_0),
		.io_in_b_0(b_304_0),
		.io_in_d_0(b_1328_0),
		.io_in_control_0_dataflow(mesh_16_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2352_0),
		.io_in_last_0(r_3376_0),
		.io_in_valid_0(r_1328_0),
		.io_out_a_0(_mesh_16_9_io_out_a_0),
		.io_out_c_0(_mesh_16_9_io_out_c_0),
		.io_out_b_0(_mesh_16_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_9_io_out_id_0),
		.io_out_last_0(_mesh_16_9_io_out_last_0),
		.io_out_valid_0(_mesh_16_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9892 == GlobalFiModInstNr[0]) || (9892 == GlobalFiModInstNr[1]) || (9892 == GlobalFiModInstNr[2]) || (9892 == GlobalFiModInstNr[3]))));
	Tile mesh_16_10(
		.clock(clock),
		.io_in_a_0(r_522_0),
		.io_in_b_0(b_336_0),
		.io_in_d_0(b_1360_0),
		.io_in_control_0_dataflow(mesh_16_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2384_0),
		.io_in_last_0(r_3408_0),
		.io_in_valid_0(r_1360_0),
		.io_out_a_0(_mesh_16_10_io_out_a_0),
		.io_out_c_0(_mesh_16_10_io_out_c_0),
		.io_out_b_0(_mesh_16_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_10_io_out_id_0),
		.io_out_last_0(_mesh_16_10_io_out_last_0),
		.io_out_valid_0(_mesh_16_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9893 == GlobalFiModInstNr[0]) || (9893 == GlobalFiModInstNr[1]) || (9893 == GlobalFiModInstNr[2]) || (9893 == GlobalFiModInstNr[3]))));
	Tile mesh_16_11(
		.clock(clock),
		.io_in_a_0(r_523_0),
		.io_in_b_0(b_368_0),
		.io_in_d_0(b_1392_0),
		.io_in_control_0_dataflow(mesh_16_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2416_0),
		.io_in_last_0(r_3440_0),
		.io_in_valid_0(r_1392_0),
		.io_out_a_0(_mesh_16_11_io_out_a_0),
		.io_out_c_0(_mesh_16_11_io_out_c_0),
		.io_out_b_0(_mesh_16_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_11_io_out_id_0),
		.io_out_last_0(_mesh_16_11_io_out_last_0),
		.io_out_valid_0(_mesh_16_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9894 == GlobalFiModInstNr[0]) || (9894 == GlobalFiModInstNr[1]) || (9894 == GlobalFiModInstNr[2]) || (9894 == GlobalFiModInstNr[3]))));
	Tile mesh_16_12(
		.clock(clock),
		.io_in_a_0(r_524_0),
		.io_in_b_0(b_400_0),
		.io_in_d_0(b_1424_0),
		.io_in_control_0_dataflow(mesh_16_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2448_0),
		.io_in_last_0(r_3472_0),
		.io_in_valid_0(r_1424_0),
		.io_out_a_0(_mesh_16_12_io_out_a_0),
		.io_out_c_0(_mesh_16_12_io_out_c_0),
		.io_out_b_0(_mesh_16_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_12_io_out_id_0),
		.io_out_last_0(_mesh_16_12_io_out_last_0),
		.io_out_valid_0(_mesh_16_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9895 == GlobalFiModInstNr[0]) || (9895 == GlobalFiModInstNr[1]) || (9895 == GlobalFiModInstNr[2]) || (9895 == GlobalFiModInstNr[3]))));
	Tile mesh_16_13(
		.clock(clock),
		.io_in_a_0(r_525_0),
		.io_in_b_0(b_432_0),
		.io_in_d_0(b_1456_0),
		.io_in_control_0_dataflow(mesh_16_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2480_0),
		.io_in_last_0(r_3504_0),
		.io_in_valid_0(r_1456_0),
		.io_out_a_0(_mesh_16_13_io_out_a_0),
		.io_out_c_0(_mesh_16_13_io_out_c_0),
		.io_out_b_0(_mesh_16_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_13_io_out_id_0),
		.io_out_last_0(_mesh_16_13_io_out_last_0),
		.io_out_valid_0(_mesh_16_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9896 == GlobalFiModInstNr[0]) || (9896 == GlobalFiModInstNr[1]) || (9896 == GlobalFiModInstNr[2]) || (9896 == GlobalFiModInstNr[3]))));
	Tile mesh_16_14(
		.clock(clock),
		.io_in_a_0(r_526_0),
		.io_in_b_0(b_464_0),
		.io_in_d_0(b_1488_0),
		.io_in_control_0_dataflow(mesh_16_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2512_0),
		.io_in_last_0(r_3536_0),
		.io_in_valid_0(r_1488_0),
		.io_out_a_0(_mesh_16_14_io_out_a_0),
		.io_out_c_0(_mesh_16_14_io_out_c_0),
		.io_out_b_0(_mesh_16_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_14_io_out_id_0),
		.io_out_last_0(_mesh_16_14_io_out_last_0),
		.io_out_valid_0(_mesh_16_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9897 == GlobalFiModInstNr[0]) || (9897 == GlobalFiModInstNr[1]) || (9897 == GlobalFiModInstNr[2]) || (9897 == GlobalFiModInstNr[3]))));
	Tile mesh_16_15(
		.clock(clock),
		.io_in_a_0(r_527_0),
		.io_in_b_0(b_496_0),
		.io_in_d_0(b_1520_0),
		.io_in_control_0_dataflow(mesh_16_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2544_0),
		.io_in_last_0(r_3568_0),
		.io_in_valid_0(r_1520_0),
		.io_out_a_0(_mesh_16_15_io_out_a_0),
		.io_out_c_0(_mesh_16_15_io_out_c_0),
		.io_out_b_0(_mesh_16_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_15_io_out_id_0),
		.io_out_last_0(_mesh_16_15_io_out_last_0),
		.io_out_valid_0(_mesh_16_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9898 == GlobalFiModInstNr[0]) || (9898 == GlobalFiModInstNr[1]) || (9898 == GlobalFiModInstNr[2]) || (9898 == GlobalFiModInstNr[3]))));
	Tile mesh_16_16(
		.clock(clock),
		.io_in_a_0(r_528_0),
		.io_in_b_0(b_528_0),
		.io_in_d_0(b_1552_0),
		.io_in_control_0_dataflow(mesh_16_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2576_0),
		.io_in_last_0(r_3600_0),
		.io_in_valid_0(r_1552_0),
		.io_out_a_0(_mesh_16_16_io_out_a_0),
		.io_out_c_0(_mesh_16_16_io_out_c_0),
		.io_out_b_0(_mesh_16_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_16_io_out_id_0),
		.io_out_last_0(_mesh_16_16_io_out_last_0),
		.io_out_valid_0(_mesh_16_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9899 == GlobalFiModInstNr[0]) || (9899 == GlobalFiModInstNr[1]) || (9899 == GlobalFiModInstNr[2]) || (9899 == GlobalFiModInstNr[3]))));
	Tile mesh_16_17(
		.clock(clock),
		.io_in_a_0(r_529_0),
		.io_in_b_0(b_560_0),
		.io_in_d_0(b_1584_0),
		.io_in_control_0_dataflow(mesh_16_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2608_0),
		.io_in_last_0(r_3632_0),
		.io_in_valid_0(r_1584_0),
		.io_out_a_0(_mesh_16_17_io_out_a_0),
		.io_out_c_0(_mesh_16_17_io_out_c_0),
		.io_out_b_0(_mesh_16_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_17_io_out_id_0),
		.io_out_last_0(_mesh_16_17_io_out_last_0),
		.io_out_valid_0(_mesh_16_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9900 == GlobalFiModInstNr[0]) || (9900 == GlobalFiModInstNr[1]) || (9900 == GlobalFiModInstNr[2]) || (9900 == GlobalFiModInstNr[3]))));
	Tile mesh_16_18(
		.clock(clock),
		.io_in_a_0(r_530_0),
		.io_in_b_0(b_592_0),
		.io_in_d_0(b_1616_0),
		.io_in_control_0_dataflow(mesh_16_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2640_0),
		.io_in_last_0(r_3664_0),
		.io_in_valid_0(r_1616_0),
		.io_out_a_0(_mesh_16_18_io_out_a_0),
		.io_out_c_0(_mesh_16_18_io_out_c_0),
		.io_out_b_0(_mesh_16_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_18_io_out_id_0),
		.io_out_last_0(_mesh_16_18_io_out_last_0),
		.io_out_valid_0(_mesh_16_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9901 == GlobalFiModInstNr[0]) || (9901 == GlobalFiModInstNr[1]) || (9901 == GlobalFiModInstNr[2]) || (9901 == GlobalFiModInstNr[3]))));
	Tile mesh_16_19(
		.clock(clock),
		.io_in_a_0(r_531_0),
		.io_in_b_0(b_624_0),
		.io_in_d_0(b_1648_0),
		.io_in_control_0_dataflow(mesh_16_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2672_0),
		.io_in_last_0(r_3696_0),
		.io_in_valid_0(r_1648_0),
		.io_out_a_0(_mesh_16_19_io_out_a_0),
		.io_out_c_0(_mesh_16_19_io_out_c_0),
		.io_out_b_0(_mesh_16_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_19_io_out_id_0),
		.io_out_last_0(_mesh_16_19_io_out_last_0),
		.io_out_valid_0(_mesh_16_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9902 == GlobalFiModInstNr[0]) || (9902 == GlobalFiModInstNr[1]) || (9902 == GlobalFiModInstNr[2]) || (9902 == GlobalFiModInstNr[3]))));
	Tile mesh_16_20(
		.clock(clock),
		.io_in_a_0(r_532_0),
		.io_in_b_0(b_656_0),
		.io_in_d_0(b_1680_0),
		.io_in_control_0_dataflow(mesh_16_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2704_0),
		.io_in_last_0(r_3728_0),
		.io_in_valid_0(r_1680_0),
		.io_out_a_0(_mesh_16_20_io_out_a_0),
		.io_out_c_0(_mesh_16_20_io_out_c_0),
		.io_out_b_0(_mesh_16_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_20_io_out_id_0),
		.io_out_last_0(_mesh_16_20_io_out_last_0),
		.io_out_valid_0(_mesh_16_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9903 == GlobalFiModInstNr[0]) || (9903 == GlobalFiModInstNr[1]) || (9903 == GlobalFiModInstNr[2]) || (9903 == GlobalFiModInstNr[3]))));
	Tile mesh_16_21(
		.clock(clock),
		.io_in_a_0(r_533_0),
		.io_in_b_0(b_688_0),
		.io_in_d_0(b_1712_0),
		.io_in_control_0_dataflow(mesh_16_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2736_0),
		.io_in_last_0(r_3760_0),
		.io_in_valid_0(r_1712_0),
		.io_out_a_0(_mesh_16_21_io_out_a_0),
		.io_out_c_0(_mesh_16_21_io_out_c_0),
		.io_out_b_0(_mesh_16_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_21_io_out_id_0),
		.io_out_last_0(_mesh_16_21_io_out_last_0),
		.io_out_valid_0(_mesh_16_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9904 == GlobalFiModInstNr[0]) || (9904 == GlobalFiModInstNr[1]) || (9904 == GlobalFiModInstNr[2]) || (9904 == GlobalFiModInstNr[3]))));
	Tile mesh_16_22(
		.clock(clock),
		.io_in_a_0(r_534_0),
		.io_in_b_0(b_720_0),
		.io_in_d_0(b_1744_0),
		.io_in_control_0_dataflow(mesh_16_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2768_0),
		.io_in_last_0(r_3792_0),
		.io_in_valid_0(r_1744_0),
		.io_out_a_0(_mesh_16_22_io_out_a_0),
		.io_out_c_0(_mesh_16_22_io_out_c_0),
		.io_out_b_0(_mesh_16_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_22_io_out_id_0),
		.io_out_last_0(_mesh_16_22_io_out_last_0),
		.io_out_valid_0(_mesh_16_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9905 == GlobalFiModInstNr[0]) || (9905 == GlobalFiModInstNr[1]) || (9905 == GlobalFiModInstNr[2]) || (9905 == GlobalFiModInstNr[3]))));
	Tile mesh_16_23(
		.clock(clock),
		.io_in_a_0(r_535_0),
		.io_in_b_0(b_752_0),
		.io_in_d_0(b_1776_0),
		.io_in_control_0_dataflow(mesh_16_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2800_0),
		.io_in_last_0(r_3824_0),
		.io_in_valid_0(r_1776_0),
		.io_out_a_0(_mesh_16_23_io_out_a_0),
		.io_out_c_0(_mesh_16_23_io_out_c_0),
		.io_out_b_0(_mesh_16_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_23_io_out_id_0),
		.io_out_last_0(_mesh_16_23_io_out_last_0),
		.io_out_valid_0(_mesh_16_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9906 == GlobalFiModInstNr[0]) || (9906 == GlobalFiModInstNr[1]) || (9906 == GlobalFiModInstNr[2]) || (9906 == GlobalFiModInstNr[3]))));
	Tile mesh_16_24(
		.clock(clock),
		.io_in_a_0(r_536_0),
		.io_in_b_0(b_784_0),
		.io_in_d_0(b_1808_0),
		.io_in_control_0_dataflow(mesh_16_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2832_0),
		.io_in_last_0(r_3856_0),
		.io_in_valid_0(r_1808_0),
		.io_out_a_0(_mesh_16_24_io_out_a_0),
		.io_out_c_0(_mesh_16_24_io_out_c_0),
		.io_out_b_0(_mesh_16_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_24_io_out_id_0),
		.io_out_last_0(_mesh_16_24_io_out_last_0),
		.io_out_valid_0(_mesh_16_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9907 == GlobalFiModInstNr[0]) || (9907 == GlobalFiModInstNr[1]) || (9907 == GlobalFiModInstNr[2]) || (9907 == GlobalFiModInstNr[3]))));
	Tile mesh_16_25(
		.clock(clock),
		.io_in_a_0(r_537_0),
		.io_in_b_0(b_816_0),
		.io_in_d_0(b_1840_0),
		.io_in_control_0_dataflow(mesh_16_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2864_0),
		.io_in_last_0(r_3888_0),
		.io_in_valid_0(r_1840_0),
		.io_out_a_0(_mesh_16_25_io_out_a_0),
		.io_out_c_0(_mesh_16_25_io_out_c_0),
		.io_out_b_0(_mesh_16_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_25_io_out_id_0),
		.io_out_last_0(_mesh_16_25_io_out_last_0),
		.io_out_valid_0(_mesh_16_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9908 == GlobalFiModInstNr[0]) || (9908 == GlobalFiModInstNr[1]) || (9908 == GlobalFiModInstNr[2]) || (9908 == GlobalFiModInstNr[3]))));
	Tile mesh_16_26(
		.clock(clock),
		.io_in_a_0(r_538_0),
		.io_in_b_0(b_848_0),
		.io_in_d_0(b_1872_0),
		.io_in_control_0_dataflow(mesh_16_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2896_0),
		.io_in_last_0(r_3920_0),
		.io_in_valid_0(r_1872_0),
		.io_out_a_0(_mesh_16_26_io_out_a_0),
		.io_out_c_0(_mesh_16_26_io_out_c_0),
		.io_out_b_0(_mesh_16_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_26_io_out_id_0),
		.io_out_last_0(_mesh_16_26_io_out_last_0),
		.io_out_valid_0(_mesh_16_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9909 == GlobalFiModInstNr[0]) || (9909 == GlobalFiModInstNr[1]) || (9909 == GlobalFiModInstNr[2]) || (9909 == GlobalFiModInstNr[3]))));
	Tile mesh_16_27(
		.clock(clock),
		.io_in_a_0(r_539_0),
		.io_in_b_0(b_880_0),
		.io_in_d_0(b_1904_0),
		.io_in_control_0_dataflow(mesh_16_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2928_0),
		.io_in_last_0(r_3952_0),
		.io_in_valid_0(r_1904_0),
		.io_out_a_0(_mesh_16_27_io_out_a_0),
		.io_out_c_0(_mesh_16_27_io_out_c_0),
		.io_out_b_0(_mesh_16_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_27_io_out_id_0),
		.io_out_last_0(_mesh_16_27_io_out_last_0),
		.io_out_valid_0(_mesh_16_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9910 == GlobalFiModInstNr[0]) || (9910 == GlobalFiModInstNr[1]) || (9910 == GlobalFiModInstNr[2]) || (9910 == GlobalFiModInstNr[3]))));
	Tile mesh_16_28(
		.clock(clock),
		.io_in_a_0(r_540_0),
		.io_in_b_0(b_912_0),
		.io_in_d_0(b_1936_0),
		.io_in_control_0_dataflow(mesh_16_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2960_0),
		.io_in_last_0(r_3984_0),
		.io_in_valid_0(r_1936_0),
		.io_out_a_0(_mesh_16_28_io_out_a_0),
		.io_out_c_0(_mesh_16_28_io_out_c_0),
		.io_out_b_0(_mesh_16_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_28_io_out_id_0),
		.io_out_last_0(_mesh_16_28_io_out_last_0),
		.io_out_valid_0(_mesh_16_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9911 == GlobalFiModInstNr[0]) || (9911 == GlobalFiModInstNr[1]) || (9911 == GlobalFiModInstNr[2]) || (9911 == GlobalFiModInstNr[3]))));
	Tile mesh_16_29(
		.clock(clock),
		.io_in_a_0(r_541_0),
		.io_in_b_0(b_944_0),
		.io_in_d_0(b_1968_0),
		.io_in_control_0_dataflow(mesh_16_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2992_0),
		.io_in_last_0(r_4016_0),
		.io_in_valid_0(r_1968_0),
		.io_out_a_0(_mesh_16_29_io_out_a_0),
		.io_out_c_0(_mesh_16_29_io_out_c_0),
		.io_out_b_0(_mesh_16_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_29_io_out_id_0),
		.io_out_last_0(_mesh_16_29_io_out_last_0),
		.io_out_valid_0(_mesh_16_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9912 == GlobalFiModInstNr[0]) || (9912 == GlobalFiModInstNr[1]) || (9912 == GlobalFiModInstNr[2]) || (9912 == GlobalFiModInstNr[3]))));
	Tile mesh_16_30(
		.clock(clock),
		.io_in_a_0(r_542_0),
		.io_in_b_0(b_976_0),
		.io_in_d_0(b_2000_0),
		.io_in_control_0_dataflow(mesh_16_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3024_0),
		.io_in_last_0(r_4048_0),
		.io_in_valid_0(r_2000_0),
		.io_out_a_0(_mesh_16_30_io_out_a_0),
		.io_out_c_0(_mesh_16_30_io_out_c_0),
		.io_out_b_0(_mesh_16_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_30_io_out_id_0),
		.io_out_last_0(_mesh_16_30_io_out_last_0),
		.io_out_valid_0(_mesh_16_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9913 == GlobalFiModInstNr[0]) || (9913 == GlobalFiModInstNr[1]) || (9913 == GlobalFiModInstNr[2]) || (9913 == GlobalFiModInstNr[3]))));
	Tile mesh_16_31(
		.clock(clock),
		.io_in_a_0(r_543_0),
		.io_in_b_0(b_1008_0),
		.io_in_d_0(b_2032_0),
		.io_in_control_0_dataflow(mesh_16_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_16_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_16_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3056_0),
		.io_in_last_0(r_4080_0),
		.io_in_valid_0(r_2032_0),
		.io_out_a_0(_mesh_16_31_io_out_a_0),
		.io_out_c_0(_mesh_16_31_io_out_c_0),
		.io_out_b_0(_mesh_16_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_16_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_16_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_16_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_16_31_io_out_id_0),
		.io_out_last_0(_mesh_16_31_io_out_last_0),
		.io_out_valid_0(_mesh_16_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9914 == GlobalFiModInstNr[0]) || (9914 == GlobalFiModInstNr[1]) || (9914 == GlobalFiModInstNr[2]) || (9914 == GlobalFiModInstNr[3]))));
	Tile mesh_17_0(
		.clock(clock),
		.io_in_a_0(r_544_0),
		.io_in_b_0(b_17_0),
		.io_in_d_0(b_1041_0),
		.io_in_control_0_dataflow(mesh_17_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2065_0),
		.io_in_last_0(r_3089_0),
		.io_in_valid_0(r_1041_0),
		.io_out_a_0(_mesh_17_0_io_out_a_0),
		.io_out_c_0(_mesh_17_0_io_out_c_0),
		.io_out_b_0(_mesh_17_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_0_io_out_id_0),
		.io_out_last_0(_mesh_17_0_io_out_last_0),
		.io_out_valid_0(_mesh_17_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9915 == GlobalFiModInstNr[0]) || (9915 == GlobalFiModInstNr[1]) || (9915 == GlobalFiModInstNr[2]) || (9915 == GlobalFiModInstNr[3]))));
	Tile mesh_17_1(
		.clock(clock),
		.io_in_a_0(r_545_0),
		.io_in_b_0(b_49_0),
		.io_in_d_0(b_1073_0),
		.io_in_control_0_dataflow(mesh_17_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2097_0),
		.io_in_last_0(r_3121_0),
		.io_in_valid_0(r_1073_0),
		.io_out_a_0(_mesh_17_1_io_out_a_0),
		.io_out_c_0(_mesh_17_1_io_out_c_0),
		.io_out_b_0(_mesh_17_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_1_io_out_id_0),
		.io_out_last_0(_mesh_17_1_io_out_last_0),
		.io_out_valid_0(_mesh_17_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9916 == GlobalFiModInstNr[0]) || (9916 == GlobalFiModInstNr[1]) || (9916 == GlobalFiModInstNr[2]) || (9916 == GlobalFiModInstNr[3]))));
	Tile mesh_17_2(
		.clock(clock),
		.io_in_a_0(r_546_0),
		.io_in_b_0(b_81_0),
		.io_in_d_0(b_1105_0),
		.io_in_control_0_dataflow(mesh_17_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2129_0),
		.io_in_last_0(r_3153_0),
		.io_in_valid_0(r_1105_0),
		.io_out_a_0(_mesh_17_2_io_out_a_0),
		.io_out_c_0(_mesh_17_2_io_out_c_0),
		.io_out_b_0(_mesh_17_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_2_io_out_id_0),
		.io_out_last_0(_mesh_17_2_io_out_last_0),
		.io_out_valid_0(_mesh_17_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9917 == GlobalFiModInstNr[0]) || (9917 == GlobalFiModInstNr[1]) || (9917 == GlobalFiModInstNr[2]) || (9917 == GlobalFiModInstNr[3]))));
	Tile mesh_17_3(
		.clock(clock),
		.io_in_a_0(r_547_0),
		.io_in_b_0(b_113_0),
		.io_in_d_0(b_1137_0),
		.io_in_control_0_dataflow(mesh_17_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2161_0),
		.io_in_last_0(r_3185_0),
		.io_in_valid_0(r_1137_0),
		.io_out_a_0(_mesh_17_3_io_out_a_0),
		.io_out_c_0(_mesh_17_3_io_out_c_0),
		.io_out_b_0(_mesh_17_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_3_io_out_id_0),
		.io_out_last_0(_mesh_17_3_io_out_last_0),
		.io_out_valid_0(_mesh_17_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9918 == GlobalFiModInstNr[0]) || (9918 == GlobalFiModInstNr[1]) || (9918 == GlobalFiModInstNr[2]) || (9918 == GlobalFiModInstNr[3]))));
	Tile mesh_17_4(
		.clock(clock),
		.io_in_a_0(r_548_0),
		.io_in_b_0(b_145_0),
		.io_in_d_0(b_1169_0),
		.io_in_control_0_dataflow(mesh_17_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2193_0),
		.io_in_last_0(r_3217_0),
		.io_in_valid_0(r_1169_0),
		.io_out_a_0(_mesh_17_4_io_out_a_0),
		.io_out_c_0(_mesh_17_4_io_out_c_0),
		.io_out_b_0(_mesh_17_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_4_io_out_id_0),
		.io_out_last_0(_mesh_17_4_io_out_last_0),
		.io_out_valid_0(_mesh_17_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9919 == GlobalFiModInstNr[0]) || (9919 == GlobalFiModInstNr[1]) || (9919 == GlobalFiModInstNr[2]) || (9919 == GlobalFiModInstNr[3]))));
	Tile mesh_17_5(
		.clock(clock),
		.io_in_a_0(r_549_0),
		.io_in_b_0(b_177_0),
		.io_in_d_0(b_1201_0),
		.io_in_control_0_dataflow(mesh_17_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2225_0),
		.io_in_last_0(r_3249_0),
		.io_in_valid_0(r_1201_0),
		.io_out_a_0(_mesh_17_5_io_out_a_0),
		.io_out_c_0(_mesh_17_5_io_out_c_0),
		.io_out_b_0(_mesh_17_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_5_io_out_id_0),
		.io_out_last_0(_mesh_17_5_io_out_last_0),
		.io_out_valid_0(_mesh_17_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9920 == GlobalFiModInstNr[0]) || (9920 == GlobalFiModInstNr[1]) || (9920 == GlobalFiModInstNr[2]) || (9920 == GlobalFiModInstNr[3]))));
	Tile mesh_17_6(
		.clock(clock),
		.io_in_a_0(r_550_0),
		.io_in_b_0(b_209_0),
		.io_in_d_0(b_1233_0),
		.io_in_control_0_dataflow(mesh_17_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2257_0),
		.io_in_last_0(r_3281_0),
		.io_in_valid_0(r_1233_0),
		.io_out_a_0(_mesh_17_6_io_out_a_0),
		.io_out_c_0(_mesh_17_6_io_out_c_0),
		.io_out_b_0(_mesh_17_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_6_io_out_id_0),
		.io_out_last_0(_mesh_17_6_io_out_last_0),
		.io_out_valid_0(_mesh_17_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9921 == GlobalFiModInstNr[0]) || (9921 == GlobalFiModInstNr[1]) || (9921 == GlobalFiModInstNr[2]) || (9921 == GlobalFiModInstNr[3]))));
	Tile mesh_17_7(
		.clock(clock),
		.io_in_a_0(r_551_0),
		.io_in_b_0(b_241_0),
		.io_in_d_0(b_1265_0),
		.io_in_control_0_dataflow(mesh_17_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2289_0),
		.io_in_last_0(r_3313_0),
		.io_in_valid_0(r_1265_0),
		.io_out_a_0(_mesh_17_7_io_out_a_0),
		.io_out_c_0(_mesh_17_7_io_out_c_0),
		.io_out_b_0(_mesh_17_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_7_io_out_id_0),
		.io_out_last_0(_mesh_17_7_io_out_last_0),
		.io_out_valid_0(_mesh_17_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9922 == GlobalFiModInstNr[0]) || (9922 == GlobalFiModInstNr[1]) || (9922 == GlobalFiModInstNr[2]) || (9922 == GlobalFiModInstNr[3]))));
	Tile mesh_17_8(
		.clock(clock),
		.io_in_a_0(r_552_0),
		.io_in_b_0(b_273_0),
		.io_in_d_0(b_1297_0),
		.io_in_control_0_dataflow(mesh_17_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2321_0),
		.io_in_last_0(r_3345_0),
		.io_in_valid_0(r_1297_0),
		.io_out_a_0(_mesh_17_8_io_out_a_0),
		.io_out_c_0(_mesh_17_8_io_out_c_0),
		.io_out_b_0(_mesh_17_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_8_io_out_id_0),
		.io_out_last_0(_mesh_17_8_io_out_last_0),
		.io_out_valid_0(_mesh_17_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9923 == GlobalFiModInstNr[0]) || (9923 == GlobalFiModInstNr[1]) || (9923 == GlobalFiModInstNr[2]) || (9923 == GlobalFiModInstNr[3]))));
	Tile mesh_17_9(
		.clock(clock),
		.io_in_a_0(r_553_0),
		.io_in_b_0(b_305_0),
		.io_in_d_0(b_1329_0),
		.io_in_control_0_dataflow(mesh_17_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2353_0),
		.io_in_last_0(r_3377_0),
		.io_in_valid_0(r_1329_0),
		.io_out_a_0(_mesh_17_9_io_out_a_0),
		.io_out_c_0(_mesh_17_9_io_out_c_0),
		.io_out_b_0(_mesh_17_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_9_io_out_id_0),
		.io_out_last_0(_mesh_17_9_io_out_last_0),
		.io_out_valid_0(_mesh_17_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9924 == GlobalFiModInstNr[0]) || (9924 == GlobalFiModInstNr[1]) || (9924 == GlobalFiModInstNr[2]) || (9924 == GlobalFiModInstNr[3]))));
	Tile mesh_17_10(
		.clock(clock),
		.io_in_a_0(r_554_0),
		.io_in_b_0(b_337_0),
		.io_in_d_0(b_1361_0),
		.io_in_control_0_dataflow(mesh_17_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2385_0),
		.io_in_last_0(r_3409_0),
		.io_in_valid_0(r_1361_0),
		.io_out_a_0(_mesh_17_10_io_out_a_0),
		.io_out_c_0(_mesh_17_10_io_out_c_0),
		.io_out_b_0(_mesh_17_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_10_io_out_id_0),
		.io_out_last_0(_mesh_17_10_io_out_last_0),
		.io_out_valid_0(_mesh_17_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9925 == GlobalFiModInstNr[0]) || (9925 == GlobalFiModInstNr[1]) || (9925 == GlobalFiModInstNr[2]) || (9925 == GlobalFiModInstNr[3]))));
	Tile mesh_17_11(
		.clock(clock),
		.io_in_a_0(r_555_0),
		.io_in_b_0(b_369_0),
		.io_in_d_0(b_1393_0),
		.io_in_control_0_dataflow(mesh_17_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2417_0),
		.io_in_last_0(r_3441_0),
		.io_in_valid_0(r_1393_0),
		.io_out_a_0(_mesh_17_11_io_out_a_0),
		.io_out_c_0(_mesh_17_11_io_out_c_0),
		.io_out_b_0(_mesh_17_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_11_io_out_id_0),
		.io_out_last_0(_mesh_17_11_io_out_last_0),
		.io_out_valid_0(_mesh_17_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9926 == GlobalFiModInstNr[0]) || (9926 == GlobalFiModInstNr[1]) || (9926 == GlobalFiModInstNr[2]) || (9926 == GlobalFiModInstNr[3]))));
	Tile mesh_17_12(
		.clock(clock),
		.io_in_a_0(r_556_0),
		.io_in_b_0(b_401_0),
		.io_in_d_0(b_1425_0),
		.io_in_control_0_dataflow(mesh_17_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2449_0),
		.io_in_last_0(r_3473_0),
		.io_in_valid_0(r_1425_0),
		.io_out_a_0(_mesh_17_12_io_out_a_0),
		.io_out_c_0(_mesh_17_12_io_out_c_0),
		.io_out_b_0(_mesh_17_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_12_io_out_id_0),
		.io_out_last_0(_mesh_17_12_io_out_last_0),
		.io_out_valid_0(_mesh_17_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9927 == GlobalFiModInstNr[0]) || (9927 == GlobalFiModInstNr[1]) || (9927 == GlobalFiModInstNr[2]) || (9927 == GlobalFiModInstNr[3]))));
	Tile mesh_17_13(
		.clock(clock),
		.io_in_a_0(r_557_0),
		.io_in_b_0(b_433_0),
		.io_in_d_0(b_1457_0),
		.io_in_control_0_dataflow(mesh_17_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2481_0),
		.io_in_last_0(r_3505_0),
		.io_in_valid_0(r_1457_0),
		.io_out_a_0(_mesh_17_13_io_out_a_0),
		.io_out_c_0(_mesh_17_13_io_out_c_0),
		.io_out_b_0(_mesh_17_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_13_io_out_id_0),
		.io_out_last_0(_mesh_17_13_io_out_last_0),
		.io_out_valid_0(_mesh_17_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9928 == GlobalFiModInstNr[0]) || (9928 == GlobalFiModInstNr[1]) || (9928 == GlobalFiModInstNr[2]) || (9928 == GlobalFiModInstNr[3]))));
	Tile mesh_17_14(
		.clock(clock),
		.io_in_a_0(r_558_0),
		.io_in_b_0(b_465_0),
		.io_in_d_0(b_1489_0),
		.io_in_control_0_dataflow(mesh_17_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2513_0),
		.io_in_last_0(r_3537_0),
		.io_in_valid_0(r_1489_0),
		.io_out_a_0(_mesh_17_14_io_out_a_0),
		.io_out_c_0(_mesh_17_14_io_out_c_0),
		.io_out_b_0(_mesh_17_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_14_io_out_id_0),
		.io_out_last_0(_mesh_17_14_io_out_last_0),
		.io_out_valid_0(_mesh_17_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9929 == GlobalFiModInstNr[0]) || (9929 == GlobalFiModInstNr[1]) || (9929 == GlobalFiModInstNr[2]) || (9929 == GlobalFiModInstNr[3]))));
	Tile mesh_17_15(
		.clock(clock),
		.io_in_a_0(r_559_0),
		.io_in_b_0(b_497_0),
		.io_in_d_0(b_1521_0),
		.io_in_control_0_dataflow(mesh_17_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2545_0),
		.io_in_last_0(r_3569_0),
		.io_in_valid_0(r_1521_0),
		.io_out_a_0(_mesh_17_15_io_out_a_0),
		.io_out_c_0(_mesh_17_15_io_out_c_0),
		.io_out_b_0(_mesh_17_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_15_io_out_id_0),
		.io_out_last_0(_mesh_17_15_io_out_last_0),
		.io_out_valid_0(_mesh_17_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9930 == GlobalFiModInstNr[0]) || (9930 == GlobalFiModInstNr[1]) || (9930 == GlobalFiModInstNr[2]) || (9930 == GlobalFiModInstNr[3]))));
	Tile mesh_17_16(
		.clock(clock),
		.io_in_a_0(r_560_0),
		.io_in_b_0(b_529_0),
		.io_in_d_0(b_1553_0),
		.io_in_control_0_dataflow(mesh_17_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2577_0),
		.io_in_last_0(r_3601_0),
		.io_in_valid_0(r_1553_0),
		.io_out_a_0(_mesh_17_16_io_out_a_0),
		.io_out_c_0(_mesh_17_16_io_out_c_0),
		.io_out_b_0(_mesh_17_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_16_io_out_id_0),
		.io_out_last_0(_mesh_17_16_io_out_last_0),
		.io_out_valid_0(_mesh_17_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9931 == GlobalFiModInstNr[0]) || (9931 == GlobalFiModInstNr[1]) || (9931 == GlobalFiModInstNr[2]) || (9931 == GlobalFiModInstNr[3]))));
	Tile mesh_17_17(
		.clock(clock),
		.io_in_a_0(r_561_0),
		.io_in_b_0(b_561_0),
		.io_in_d_0(b_1585_0),
		.io_in_control_0_dataflow(mesh_17_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2609_0),
		.io_in_last_0(r_3633_0),
		.io_in_valid_0(r_1585_0),
		.io_out_a_0(_mesh_17_17_io_out_a_0),
		.io_out_c_0(_mesh_17_17_io_out_c_0),
		.io_out_b_0(_mesh_17_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_17_io_out_id_0),
		.io_out_last_0(_mesh_17_17_io_out_last_0),
		.io_out_valid_0(_mesh_17_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9932 == GlobalFiModInstNr[0]) || (9932 == GlobalFiModInstNr[1]) || (9932 == GlobalFiModInstNr[2]) || (9932 == GlobalFiModInstNr[3]))));
	Tile mesh_17_18(
		.clock(clock),
		.io_in_a_0(r_562_0),
		.io_in_b_0(b_593_0),
		.io_in_d_0(b_1617_0),
		.io_in_control_0_dataflow(mesh_17_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2641_0),
		.io_in_last_0(r_3665_0),
		.io_in_valid_0(r_1617_0),
		.io_out_a_0(_mesh_17_18_io_out_a_0),
		.io_out_c_0(_mesh_17_18_io_out_c_0),
		.io_out_b_0(_mesh_17_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_18_io_out_id_0),
		.io_out_last_0(_mesh_17_18_io_out_last_0),
		.io_out_valid_0(_mesh_17_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9933 == GlobalFiModInstNr[0]) || (9933 == GlobalFiModInstNr[1]) || (9933 == GlobalFiModInstNr[2]) || (9933 == GlobalFiModInstNr[3]))));
	Tile mesh_17_19(
		.clock(clock),
		.io_in_a_0(r_563_0),
		.io_in_b_0(b_625_0),
		.io_in_d_0(b_1649_0),
		.io_in_control_0_dataflow(mesh_17_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2673_0),
		.io_in_last_0(r_3697_0),
		.io_in_valid_0(r_1649_0),
		.io_out_a_0(_mesh_17_19_io_out_a_0),
		.io_out_c_0(_mesh_17_19_io_out_c_0),
		.io_out_b_0(_mesh_17_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_19_io_out_id_0),
		.io_out_last_0(_mesh_17_19_io_out_last_0),
		.io_out_valid_0(_mesh_17_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9934 == GlobalFiModInstNr[0]) || (9934 == GlobalFiModInstNr[1]) || (9934 == GlobalFiModInstNr[2]) || (9934 == GlobalFiModInstNr[3]))));
	Tile mesh_17_20(
		.clock(clock),
		.io_in_a_0(r_564_0),
		.io_in_b_0(b_657_0),
		.io_in_d_0(b_1681_0),
		.io_in_control_0_dataflow(mesh_17_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2705_0),
		.io_in_last_0(r_3729_0),
		.io_in_valid_0(r_1681_0),
		.io_out_a_0(_mesh_17_20_io_out_a_0),
		.io_out_c_0(_mesh_17_20_io_out_c_0),
		.io_out_b_0(_mesh_17_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_20_io_out_id_0),
		.io_out_last_0(_mesh_17_20_io_out_last_0),
		.io_out_valid_0(_mesh_17_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9935 == GlobalFiModInstNr[0]) || (9935 == GlobalFiModInstNr[1]) || (9935 == GlobalFiModInstNr[2]) || (9935 == GlobalFiModInstNr[3]))));
	Tile mesh_17_21(
		.clock(clock),
		.io_in_a_0(r_565_0),
		.io_in_b_0(b_689_0),
		.io_in_d_0(b_1713_0),
		.io_in_control_0_dataflow(mesh_17_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2737_0),
		.io_in_last_0(r_3761_0),
		.io_in_valid_0(r_1713_0),
		.io_out_a_0(_mesh_17_21_io_out_a_0),
		.io_out_c_0(_mesh_17_21_io_out_c_0),
		.io_out_b_0(_mesh_17_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_21_io_out_id_0),
		.io_out_last_0(_mesh_17_21_io_out_last_0),
		.io_out_valid_0(_mesh_17_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9936 == GlobalFiModInstNr[0]) || (9936 == GlobalFiModInstNr[1]) || (9936 == GlobalFiModInstNr[2]) || (9936 == GlobalFiModInstNr[3]))));
	Tile mesh_17_22(
		.clock(clock),
		.io_in_a_0(r_566_0),
		.io_in_b_0(b_721_0),
		.io_in_d_0(b_1745_0),
		.io_in_control_0_dataflow(mesh_17_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2769_0),
		.io_in_last_0(r_3793_0),
		.io_in_valid_0(r_1745_0),
		.io_out_a_0(_mesh_17_22_io_out_a_0),
		.io_out_c_0(_mesh_17_22_io_out_c_0),
		.io_out_b_0(_mesh_17_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_22_io_out_id_0),
		.io_out_last_0(_mesh_17_22_io_out_last_0),
		.io_out_valid_0(_mesh_17_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9937 == GlobalFiModInstNr[0]) || (9937 == GlobalFiModInstNr[1]) || (9937 == GlobalFiModInstNr[2]) || (9937 == GlobalFiModInstNr[3]))));
	Tile mesh_17_23(
		.clock(clock),
		.io_in_a_0(r_567_0),
		.io_in_b_0(b_753_0),
		.io_in_d_0(b_1777_0),
		.io_in_control_0_dataflow(mesh_17_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2801_0),
		.io_in_last_0(r_3825_0),
		.io_in_valid_0(r_1777_0),
		.io_out_a_0(_mesh_17_23_io_out_a_0),
		.io_out_c_0(_mesh_17_23_io_out_c_0),
		.io_out_b_0(_mesh_17_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_23_io_out_id_0),
		.io_out_last_0(_mesh_17_23_io_out_last_0),
		.io_out_valid_0(_mesh_17_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9938 == GlobalFiModInstNr[0]) || (9938 == GlobalFiModInstNr[1]) || (9938 == GlobalFiModInstNr[2]) || (9938 == GlobalFiModInstNr[3]))));
	Tile mesh_17_24(
		.clock(clock),
		.io_in_a_0(r_568_0),
		.io_in_b_0(b_785_0),
		.io_in_d_0(b_1809_0),
		.io_in_control_0_dataflow(mesh_17_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2833_0),
		.io_in_last_0(r_3857_0),
		.io_in_valid_0(r_1809_0),
		.io_out_a_0(_mesh_17_24_io_out_a_0),
		.io_out_c_0(_mesh_17_24_io_out_c_0),
		.io_out_b_0(_mesh_17_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_24_io_out_id_0),
		.io_out_last_0(_mesh_17_24_io_out_last_0),
		.io_out_valid_0(_mesh_17_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9939 == GlobalFiModInstNr[0]) || (9939 == GlobalFiModInstNr[1]) || (9939 == GlobalFiModInstNr[2]) || (9939 == GlobalFiModInstNr[3]))));
	Tile mesh_17_25(
		.clock(clock),
		.io_in_a_0(r_569_0),
		.io_in_b_0(b_817_0),
		.io_in_d_0(b_1841_0),
		.io_in_control_0_dataflow(mesh_17_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2865_0),
		.io_in_last_0(r_3889_0),
		.io_in_valid_0(r_1841_0),
		.io_out_a_0(_mesh_17_25_io_out_a_0),
		.io_out_c_0(_mesh_17_25_io_out_c_0),
		.io_out_b_0(_mesh_17_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_25_io_out_id_0),
		.io_out_last_0(_mesh_17_25_io_out_last_0),
		.io_out_valid_0(_mesh_17_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9940 == GlobalFiModInstNr[0]) || (9940 == GlobalFiModInstNr[1]) || (9940 == GlobalFiModInstNr[2]) || (9940 == GlobalFiModInstNr[3]))));
	Tile mesh_17_26(
		.clock(clock),
		.io_in_a_0(r_570_0),
		.io_in_b_0(b_849_0),
		.io_in_d_0(b_1873_0),
		.io_in_control_0_dataflow(mesh_17_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2897_0),
		.io_in_last_0(r_3921_0),
		.io_in_valid_0(r_1873_0),
		.io_out_a_0(_mesh_17_26_io_out_a_0),
		.io_out_c_0(_mesh_17_26_io_out_c_0),
		.io_out_b_0(_mesh_17_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_26_io_out_id_0),
		.io_out_last_0(_mesh_17_26_io_out_last_0),
		.io_out_valid_0(_mesh_17_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9941 == GlobalFiModInstNr[0]) || (9941 == GlobalFiModInstNr[1]) || (9941 == GlobalFiModInstNr[2]) || (9941 == GlobalFiModInstNr[3]))));
	Tile mesh_17_27(
		.clock(clock),
		.io_in_a_0(r_571_0),
		.io_in_b_0(b_881_0),
		.io_in_d_0(b_1905_0),
		.io_in_control_0_dataflow(mesh_17_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2929_0),
		.io_in_last_0(r_3953_0),
		.io_in_valid_0(r_1905_0),
		.io_out_a_0(_mesh_17_27_io_out_a_0),
		.io_out_c_0(_mesh_17_27_io_out_c_0),
		.io_out_b_0(_mesh_17_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_27_io_out_id_0),
		.io_out_last_0(_mesh_17_27_io_out_last_0),
		.io_out_valid_0(_mesh_17_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9942 == GlobalFiModInstNr[0]) || (9942 == GlobalFiModInstNr[1]) || (9942 == GlobalFiModInstNr[2]) || (9942 == GlobalFiModInstNr[3]))));
	Tile mesh_17_28(
		.clock(clock),
		.io_in_a_0(r_572_0),
		.io_in_b_0(b_913_0),
		.io_in_d_0(b_1937_0),
		.io_in_control_0_dataflow(mesh_17_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2961_0),
		.io_in_last_0(r_3985_0),
		.io_in_valid_0(r_1937_0),
		.io_out_a_0(_mesh_17_28_io_out_a_0),
		.io_out_c_0(_mesh_17_28_io_out_c_0),
		.io_out_b_0(_mesh_17_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_28_io_out_id_0),
		.io_out_last_0(_mesh_17_28_io_out_last_0),
		.io_out_valid_0(_mesh_17_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9943 == GlobalFiModInstNr[0]) || (9943 == GlobalFiModInstNr[1]) || (9943 == GlobalFiModInstNr[2]) || (9943 == GlobalFiModInstNr[3]))));
	Tile mesh_17_29(
		.clock(clock),
		.io_in_a_0(r_573_0),
		.io_in_b_0(b_945_0),
		.io_in_d_0(b_1969_0),
		.io_in_control_0_dataflow(mesh_17_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2993_0),
		.io_in_last_0(r_4017_0),
		.io_in_valid_0(r_1969_0),
		.io_out_a_0(_mesh_17_29_io_out_a_0),
		.io_out_c_0(_mesh_17_29_io_out_c_0),
		.io_out_b_0(_mesh_17_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_29_io_out_id_0),
		.io_out_last_0(_mesh_17_29_io_out_last_0),
		.io_out_valid_0(_mesh_17_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9944 == GlobalFiModInstNr[0]) || (9944 == GlobalFiModInstNr[1]) || (9944 == GlobalFiModInstNr[2]) || (9944 == GlobalFiModInstNr[3]))));
	Tile mesh_17_30(
		.clock(clock),
		.io_in_a_0(r_574_0),
		.io_in_b_0(b_977_0),
		.io_in_d_0(b_2001_0),
		.io_in_control_0_dataflow(mesh_17_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3025_0),
		.io_in_last_0(r_4049_0),
		.io_in_valid_0(r_2001_0),
		.io_out_a_0(_mesh_17_30_io_out_a_0),
		.io_out_c_0(_mesh_17_30_io_out_c_0),
		.io_out_b_0(_mesh_17_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_30_io_out_id_0),
		.io_out_last_0(_mesh_17_30_io_out_last_0),
		.io_out_valid_0(_mesh_17_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9945 == GlobalFiModInstNr[0]) || (9945 == GlobalFiModInstNr[1]) || (9945 == GlobalFiModInstNr[2]) || (9945 == GlobalFiModInstNr[3]))));
	Tile mesh_17_31(
		.clock(clock),
		.io_in_a_0(r_575_0),
		.io_in_b_0(b_1009_0),
		.io_in_d_0(b_2033_0),
		.io_in_control_0_dataflow(mesh_17_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_17_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_17_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3057_0),
		.io_in_last_0(r_4081_0),
		.io_in_valid_0(r_2033_0),
		.io_out_a_0(_mesh_17_31_io_out_a_0),
		.io_out_c_0(_mesh_17_31_io_out_c_0),
		.io_out_b_0(_mesh_17_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_17_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_17_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_17_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_17_31_io_out_id_0),
		.io_out_last_0(_mesh_17_31_io_out_last_0),
		.io_out_valid_0(_mesh_17_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9946 == GlobalFiModInstNr[0]) || (9946 == GlobalFiModInstNr[1]) || (9946 == GlobalFiModInstNr[2]) || (9946 == GlobalFiModInstNr[3]))));
	Tile mesh_18_0(
		.clock(clock),
		.io_in_a_0(r_576_0),
		.io_in_b_0(b_18_0),
		.io_in_d_0(b_1042_0),
		.io_in_control_0_dataflow(mesh_18_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2066_0),
		.io_in_last_0(r_3090_0),
		.io_in_valid_0(r_1042_0),
		.io_out_a_0(_mesh_18_0_io_out_a_0),
		.io_out_c_0(_mesh_18_0_io_out_c_0),
		.io_out_b_0(_mesh_18_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_0_io_out_id_0),
		.io_out_last_0(_mesh_18_0_io_out_last_0),
		.io_out_valid_0(_mesh_18_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9947 == GlobalFiModInstNr[0]) || (9947 == GlobalFiModInstNr[1]) || (9947 == GlobalFiModInstNr[2]) || (9947 == GlobalFiModInstNr[3]))));
	Tile mesh_18_1(
		.clock(clock),
		.io_in_a_0(r_577_0),
		.io_in_b_0(b_50_0),
		.io_in_d_0(b_1074_0),
		.io_in_control_0_dataflow(mesh_18_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2098_0),
		.io_in_last_0(r_3122_0),
		.io_in_valid_0(r_1074_0),
		.io_out_a_0(_mesh_18_1_io_out_a_0),
		.io_out_c_0(_mesh_18_1_io_out_c_0),
		.io_out_b_0(_mesh_18_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_1_io_out_id_0),
		.io_out_last_0(_mesh_18_1_io_out_last_0),
		.io_out_valid_0(_mesh_18_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9948 == GlobalFiModInstNr[0]) || (9948 == GlobalFiModInstNr[1]) || (9948 == GlobalFiModInstNr[2]) || (9948 == GlobalFiModInstNr[3]))));
	Tile mesh_18_2(
		.clock(clock),
		.io_in_a_0(r_578_0),
		.io_in_b_0(b_82_0),
		.io_in_d_0(b_1106_0),
		.io_in_control_0_dataflow(mesh_18_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2130_0),
		.io_in_last_0(r_3154_0),
		.io_in_valid_0(r_1106_0),
		.io_out_a_0(_mesh_18_2_io_out_a_0),
		.io_out_c_0(_mesh_18_2_io_out_c_0),
		.io_out_b_0(_mesh_18_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_2_io_out_id_0),
		.io_out_last_0(_mesh_18_2_io_out_last_0),
		.io_out_valid_0(_mesh_18_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9949 == GlobalFiModInstNr[0]) || (9949 == GlobalFiModInstNr[1]) || (9949 == GlobalFiModInstNr[2]) || (9949 == GlobalFiModInstNr[3]))));
	Tile mesh_18_3(
		.clock(clock),
		.io_in_a_0(r_579_0),
		.io_in_b_0(b_114_0),
		.io_in_d_0(b_1138_0),
		.io_in_control_0_dataflow(mesh_18_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2162_0),
		.io_in_last_0(r_3186_0),
		.io_in_valid_0(r_1138_0),
		.io_out_a_0(_mesh_18_3_io_out_a_0),
		.io_out_c_0(_mesh_18_3_io_out_c_0),
		.io_out_b_0(_mesh_18_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_3_io_out_id_0),
		.io_out_last_0(_mesh_18_3_io_out_last_0),
		.io_out_valid_0(_mesh_18_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9950 == GlobalFiModInstNr[0]) || (9950 == GlobalFiModInstNr[1]) || (9950 == GlobalFiModInstNr[2]) || (9950 == GlobalFiModInstNr[3]))));
	Tile mesh_18_4(
		.clock(clock),
		.io_in_a_0(r_580_0),
		.io_in_b_0(b_146_0),
		.io_in_d_0(b_1170_0),
		.io_in_control_0_dataflow(mesh_18_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2194_0),
		.io_in_last_0(r_3218_0),
		.io_in_valid_0(r_1170_0),
		.io_out_a_0(_mesh_18_4_io_out_a_0),
		.io_out_c_0(_mesh_18_4_io_out_c_0),
		.io_out_b_0(_mesh_18_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_4_io_out_id_0),
		.io_out_last_0(_mesh_18_4_io_out_last_0),
		.io_out_valid_0(_mesh_18_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9951 == GlobalFiModInstNr[0]) || (9951 == GlobalFiModInstNr[1]) || (9951 == GlobalFiModInstNr[2]) || (9951 == GlobalFiModInstNr[3]))));
	Tile mesh_18_5(
		.clock(clock),
		.io_in_a_0(r_581_0),
		.io_in_b_0(b_178_0),
		.io_in_d_0(b_1202_0),
		.io_in_control_0_dataflow(mesh_18_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2226_0),
		.io_in_last_0(r_3250_0),
		.io_in_valid_0(r_1202_0),
		.io_out_a_0(_mesh_18_5_io_out_a_0),
		.io_out_c_0(_mesh_18_5_io_out_c_0),
		.io_out_b_0(_mesh_18_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_5_io_out_id_0),
		.io_out_last_0(_mesh_18_5_io_out_last_0),
		.io_out_valid_0(_mesh_18_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9952 == GlobalFiModInstNr[0]) || (9952 == GlobalFiModInstNr[1]) || (9952 == GlobalFiModInstNr[2]) || (9952 == GlobalFiModInstNr[3]))));
	Tile mesh_18_6(
		.clock(clock),
		.io_in_a_0(r_582_0),
		.io_in_b_0(b_210_0),
		.io_in_d_0(b_1234_0),
		.io_in_control_0_dataflow(mesh_18_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2258_0),
		.io_in_last_0(r_3282_0),
		.io_in_valid_0(r_1234_0),
		.io_out_a_0(_mesh_18_6_io_out_a_0),
		.io_out_c_0(_mesh_18_6_io_out_c_0),
		.io_out_b_0(_mesh_18_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_6_io_out_id_0),
		.io_out_last_0(_mesh_18_6_io_out_last_0),
		.io_out_valid_0(_mesh_18_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9953 == GlobalFiModInstNr[0]) || (9953 == GlobalFiModInstNr[1]) || (9953 == GlobalFiModInstNr[2]) || (9953 == GlobalFiModInstNr[3]))));
	Tile mesh_18_7(
		.clock(clock),
		.io_in_a_0(r_583_0),
		.io_in_b_0(b_242_0),
		.io_in_d_0(b_1266_0),
		.io_in_control_0_dataflow(mesh_18_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2290_0),
		.io_in_last_0(r_3314_0),
		.io_in_valid_0(r_1266_0),
		.io_out_a_0(_mesh_18_7_io_out_a_0),
		.io_out_c_0(_mesh_18_7_io_out_c_0),
		.io_out_b_0(_mesh_18_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_7_io_out_id_0),
		.io_out_last_0(_mesh_18_7_io_out_last_0),
		.io_out_valid_0(_mesh_18_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9954 == GlobalFiModInstNr[0]) || (9954 == GlobalFiModInstNr[1]) || (9954 == GlobalFiModInstNr[2]) || (9954 == GlobalFiModInstNr[3]))));
	Tile mesh_18_8(
		.clock(clock),
		.io_in_a_0(r_584_0),
		.io_in_b_0(b_274_0),
		.io_in_d_0(b_1298_0),
		.io_in_control_0_dataflow(mesh_18_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2322_0),
		.io_in_last_0(r_3346_0),
		.io_in_valid_0(r_1298_0),
		.io_out_a_0(_mesh_18_8_io_out_a_0),
		.io_out_c_0(_mesh_18_8_io_out_c_0),
		.io_out_b_0(_mesh_18_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_8_io_out_id_0),
		.io_out_last_0(_mesh_18_8_io_out_last_0),
		.io_out_valid_0(_mesh_18_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9955 == GlobalFiModInstNr[0]) || (9955 == GlobalFiModInstNr[1]) || (9955 == GlobalFiModInstNr[2]) || (9955 == GlobalFiModInstNr[3]))));
	Tile mesh_18_9(
		.clock(clock),
		.io_in_a_0(r_585_0),
		.io_in_b_0(b_306_0),
		.io_in_d_0(b_1330_0),
		.io_in_control_0_dataflow(mesh_18_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2354_0),
		.io_in_last_0(r_3378_0),
		.io_in_valid_0(r_1330_0),
		.io_out_a_0(_mesh_18_9_io_out_a_0),
		.io_out_c_0(_mesh_18_9_io_out_c_0),
		.io_out_b_0(_mesh_18_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_9_io_out_id_0),
		.io_out_last_0(_mesh_18_9_io_out_last_0),
		.io_out_valid_0(_mesh_18_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9956 == GlobalFiModInstNr[0]) || (9956 == GlobalFiModInstNr[1]) || (9956 == GlobalFiModInstNr[2]) || (9956 == GlobalFiModInstNr[3]))));
	Tile mesh_18_10(
		.clock(clock),
		.io_in_a_0(r_586_0),
		.io_in_b_0(b_338_0),
		.io_in_d_0(b_1362_0),
		.io_in_control_0_dataflow(mesh_18_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2386_0),
		.io_in_last_0(r_3410_0),
		.io_in_valid_0(r_1362_0),
		.io_out_a_0(_mesh_18_10_io_out_a_0),
		.io_out_c_0(_mesh_18_10_io_out_c_0),
		.io_out_b_0(_mesh_18_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_10_io_out_id_0),
		.io_out_last_0(_mesh_18_10_io_out_last_0),
		.io_out_valid_0(_mesh_18_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9957 == GlobalFiModInstNr[0]) || (9957 == GlobalFiModInstNr[1]) || (9957 == GlobalFiModInstNr[2]) || (9957 == GlobalFiModInstNr[3]))));
	Tile mesh_18_11(
		.clock(clock),
		.io_in_a_0(r_587_0),
		.io_in_b_0(b_370_0),
		.io_in_d_0(b_1394_0),
		.io_in_control_0_dataflow(mesh_18_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2418_0),
		.io_in_last_0(r_3442_0),
		.io_in_valid_0(r_1394_0),
		.io_out_a_0(_mesh_18_11_io_out_a_0),
		.io_out_c_0(_mesh_18_11_io_out_c_0),
		.io_out_b_0(_mesh_18_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_11_io_out_id_0),
		.io_out_last_0(_mesh_18_11_io_out_last_0),
		.io_out_valid_0(_mesh_18_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9958 == GlobalFiModInstNr[0]) || (9958 == GlobalFiModInstNr[1]) || (9958 == GlobalFiModInstNr[2]) || (9958 == GlobalFiModInstNr[3]))));
	Tile mesh_18_12(
		.clock(clock),
		.io_in_a_0(r_588_0),
		.io_in_b_0(b_402_0),
		.io_in_d_0(b_1426_0),
		.io_in_control_0_dataflow(mesh_18_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2450_0),
		.io_in_last_0(r_3474_0),
		.io_in_valid_0(r_1426_0),
		.io_out_a_0(_mesh_18_12_io_out_a_0),
		.io_out_c_0(_mesh_18_12_io_out_c_0),
		.io_out_b_0(_mesh_18_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_12_io_out_id_0),
		.io_out_last_0(_mesh_18_12_io_out_last_0),
		.io_out_valid_0(_mesh_18_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9959 == GlobalFiModInstNr[0]) || (9959 == GlobalFiModInstNr[1]) || (9959 == GlobalFiModInstNr[2]) || (9959 == GlobalFiModInstNr[3]))));
	Tile mesh_18_13(
		.clock(clock),
		.io_in_a_0(r_589_0),
		.io_in_b_0(b_434_0),
		.io_in_d_0(b_1458_0),
		.io_in_control_0_dataflow(mesh_18_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2482_0),
		.io_in_last_0(r_3506_0),
		.io_in_valid_0(r_1458_0),
		.io_out_a_0(_mesh_18_13_io_out_a_0),
		.io_out_c_0(_mesh_18_13_io_out_c_0),
		.io_out_b_0(_mesh_18_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_13_io_out_id_0),
		.io_out_last_0(_mesh_18_13_io_out_last_0),
		.io_out_valid_0(_mesh_18_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9960 == GlobalFiModInstNr[0]) || (9960 == GlobalFiModInstNr[1]) || (9960 == GlobalFiModInstNr[2]) || (9960 == GlobalFiModInstNr[3]))));
	Tile mesh_18_14(
		.clock(clock),
		.io_in_a_0(r_590_0),
		.io_in_b_0(b_466_0),
		.io_in_d_0(b_1490_0),
		.io_in_control_0_dataflow(mesh_18_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2514_0),
		.io_in_last_0(r_3538_0),
		.io_in_valid_0(r_1490_0),
		.io_out_a_0(_mesh_18_14_io_out_a_0),
		.io_out_c_0(_mesh_18_14_io_out_c_0),
		.io_out_b_0(_mesh_18_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_14_io_out_id_0),
		.io_out_last_0(_mesh_18_14_io_out_last_0),
		.io_out_valid_0(_mesh_18_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9961 == GlobalFiModInstNr[0]) || (9961 == GlobalFiModInstNr[1]) || (9961 == GlobalFiModInstNr[2]) || (9961 == GlobalFiModInstNr[3]))));
	Tile mesh_18_15(
		.clock(clock),
		.io_in_a_0(r_591_0),
		.io_in_b_0(b_498_0),
		.io_in_d_0(b_1522_0),
		.io_in_control_0_dataflow(mesh_18_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2546_0),
		.io_in_last_0(r_3570_0),
		.io_in_valid_0(r_1522_0),
		.io_out_a_0(_mesh_18_15_io_out_a_0),
		.io_out_c_0(_mesh_18_15_io_out_c_0),
		.io_out_b_0(_mesh_18_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_15_io_out_id_0),
		.io_out_last_0(_mesh_18_15_io_out_last_0),
		.io_out_valid_0(_mesh_18_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9962 == GlobalFiModInstNr[0]) || (9962 == GlobalFiModInstNr[1]) || (9962 == GlobalFiModInstNr[2]) || (9962 == GlobalFiModInstNr[3]))));
	Tile mesh_18_16(
		.clock(clock),
		.io_in_a_0(r_592_0),
		.io_in_b_0(b_530_0),
		.io_in_d_0(b_1554_0),
		.io_in_control_0_dataflow(mesh_18_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2578_0),
		.io_in_last_0(r_3602_0),
		.io_in_valid_0(r_1554_0),
		.io_out_a_0(_mesh_18_16_io_out_a_0),
		.io_out_c_0(_mesh_18_16_io_out_c_0),
		.io_out_b_0(_mesh_18_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_16_io_out_id_0),
		.io_out_last_0(_mesh_18_16_io_out_last_0),
		.io_out_valid_0(_mesh_18_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9963 == GlobalFiModInstNr[0]) || (9963 == GlobalFiModInstNr[1]) || (9963 == GlobalFiModInstNr[2]) || (9963 == GlobalFiModInstNr[3]))));
	Tile mesh_18_17(
		.clock(clock),
		.io_in_a_0(r_593_0),
		.io_in_b_0(b_562_0),
		.io_in_d_0(b_1586_0),
		.io_in_control_0_dataflow(mesh_18_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2610_0),
		.io_in_last_0(r_3634_0),
		.io_in_valid_0(r_1586_0),
		.io_out_a_0(_mesh_18_17_io_out_a_0),
		.io_out_c_0(_mesh_18_17_io_out_c_0),
		.io_out_b_0(_mesh_18_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_17_io_out_id_0),
		.io_out_last_0(_mesh_18_17_io_out_last_0),
		.io_out_valid_0(_mesh_18_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9964 == GlobalFiModInstNr[0]) || (9964 == GlobalFiModInstNr[1]) || (9964 == GlobalFiModInstNr[2]) || (9964 == GlobalFiModInstNr[3]))));
	Tile mesh_18_18(
		.clock(clock),
		.io_in_a_0(r_594_0),
		.io_in_b_0(b_594_0),
		.io_in_d_0(b_1618_0),
		.io_in_control_0_dataflow(mesh_18_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2642_0),
		.io_in_last_0(r_3666_0),
		.io_in_valid_0(r_1618_0),
		.io_out_a_0(_mesh_18_18_io_out_a_0),
		.io_out_c_0(_mesh_18_18_io_out_c_0),
		.io_out_b_0(_mesh_18_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_18_io_out_id_0),
		.io_out_last_0(_mesh_18_18_io_out_last_0),
		.io_out_valid_0(_mesh_18_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9965 == GlobalFiModInstNr[0]) || (9965 == GlobalFiModInstNr[1]) || (9965 == GlobalFiModInstNr[2]) || (9965 == GlobalFiModInstNr[3]))));
	Tile mesh_18_19(
		.clock(clock),
		.io_in_a_0(r_595_0),
		.io_in_b_0(b_626_0),
		.io_in_d_0(b_1650_0),
		.io_in_control_0_dataflow(mesh_18_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2674_0),
		.io_in_last_0(r_3698_0),
		.io_in_valid_0(r_1650_0),
		.io_out_a_0(_mesh_18_19_io_out_a_0),
		.io_out_c_0(_mesh_18_19_io_out_c_0),
		.io_out_b_0(_mesh_18_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_19_io_out_id_0),
		.io_out_last_0(_mesh_18_19_io_out_last_0),
		.io_out_valid_0(_mesh_18_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9966 == GlobalFiModInstNr[0]) || (9966 == GlobalFiModInstNr[1]) || (9966 == GlobalFiModInstNr[2]) || (9966 == GlobalFiModInstNr[3]))));
	Tile mesh_18_20(
		.clock(clock),
		.io_in_a_0(r_596_0),
		.io_in_b_0(b_658_0),
		.io_in_d_0(b_1682_0),
		.io_in_control_0_dataflow(mesh_18_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2706_0),
		.io_in_last_0(r_3730_0),
		.io_in_valid_0(r_1682_0),
		.io_out_a_0(_mesh_18_20_io_out_a_0),
		.io_out_c_0(_mesh_18_20_io_out_c_0),
		.io_out_b_0(_mesh_18_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_20_io_out_id_0),
		.io_out_last_0(_mesh_18_20_io_out_last_0),
		.io_out_valid_0(_mesh_18_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9967 == GlobalFiModInstNr[0]) || (9967 == GlobalFiModInstNr[1]) || (9967 == GlobalFiModInstNr[2]) || (9967 == GlobalFiModInstNr[3]))));
	Tile mesh_18_21(
		.clock(clock),
		.io_in_a_0(r_597_0),
		.io_in_b_0(b_690_0),
		.io_in_d_0(b_1714_0),
		.io_in_control_0_dataflow(mesh_18_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2738_0),
		.io_in_last_0(r_3762_0),
		.io_in_valid_0(r_1714_0),
		.io_out_a_0(_mesh_18_21_io_out_a_0),
		.io_out_c_0(_mesh_18_21_io_out_c_0),
		.io_out_b_0(_mesh_18_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_21_io_out_id_0),
		.io_out_last_0(_mesh_18_21_io_out_last_0),
		.io_out_valid_0(_mesh_18_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9968 == GlobalFiModInstNr[0]) || (9968 == GlobalFiModInstNr[1]) || (9968 == GlobalFiModInstNr[2]) || (9968 == GlobalFiModInstNr[3]))));
	Tile mesh_18_22(
		.clock(clock),
		.io_in_a_0(r_598_0),
		.io_in_b_0(b_722_0),
		.io_in_d_0(b_1746_0),
		.io_in_control_0_dataflow(mesh_18_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2770_0),
		.io_in_last_0(r_3794_0),
		.io_in_valid_0(r_1746_0),
		.io_out_a_0(_mesh_18_22_io_out_a_0),
		.io_out_c_0(_mesh_18_22_io_out_c_0),
		.io_out_b_0(_mesh_18_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_22_io_out_id_0),
		.io_out_last_0(_mesh_18_22_io_out_last_0),
		.io_out_valid_0(_mesh_18_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9969 == GlobalFiModInstNr[0]) || (9969 == GlobalFiModInstNr[1]) || (9969 == GlobalFiModInstNr[2]) || (9969 == GlobalFiModInstNr[3]))));
	Tile mesh_18_23(
		.clock(clock),
		.io_in_a_0(r_599_0),
		.io_in_b_0(b_754_0),
		.io_in_d_0(b_1778_0),
		.io_in_control_0_dataflow(mesh_18_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2802_0),
		.io_in_last_0(r_3826_0),
		.io_in_valid_0(r_1778_0),
		.io_out_a_0(_mesh_18_23_io_out_a_0),
		.io_out_c_0(_mesh_18_23_io_out_c_0),
		.io_out_b_0(_mesh_18_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_23_io_out_id_0),
		.io_out_last_0(_mesh_18_23_io_out_last_0),
		.io_out_valid_0(_mesh_18_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9970 == GlobalFiModInstNr[0]) || (9970 == GlobalFiModInstNr[1]) || (9970 == GlobalFiModInstNr[2]) || (9970 == GlobalFiModInstNr[3]))));
	Tile mesh_18_24(
		.clock(clock),
		.io_in_a_0(r_600_0),
		.io_in_b_0(b_786_0),
		.io_in_d_0(b_1810_0),
		.io_in_control_0_dataflow(mesh_18_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2834_0),
		.io_in_last_0(r_3858_0),
		.io_in_valid_0(r_1810_0),
		.io_out_a_0(_mesh_18_24_io_out_a_0),
		.io_out_c_0(_mesh_18_24_io_out_c_0),
		.io_out_b_0(_mesh_18_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_24_io_out_id_0),
		.io_out_last_0(_mesh_18_24_io_out_last_0),
		.io_out_valid_0(_mesh_18_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9971 == GlobalFiModInstNr[0]) || (9971 == GlobalFiModInstNr[1]) || (9971 == GlobalFiModInstNr[2]) || (9971 == GlobalFiModInstNr[3]))));
	Tile mesh_18_25(
		.clock(clock),
		.io_in_a_0(r_601_0),
		.io_in_b_0(b_818_0),
		.io_in_d_0(b_1842_0),
		.io_in_control_0_dataflow(mesh_18_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2866_0),
		.io_in_last_0(r_3890_0),
		.io_in_valid_0(r_1842_0),
		.io_out_a_0(_mesh_18_25_io_out_a_0),
		.io_out_c_0(_mesh_18_25_io_out_c_0),
		.io_out_b_0(_mesh_18_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_25_io_out_id_0),
		.io_out_last_0(_mesh_18_25_io_out_last_0),
		.io_out_valid_0(_mesh_18_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9972 == GlobalFiModInstNr[0]) || (9972 == GlobalFiModInstNr[1]) || (9972 == GlobalFiModInstNr[2]) || (9972 == GlobalFiModInstNr[3]))));
	Tile mesh_18_26(
		.clock(clock),
		.io_in_a_0(r_602_0),
		.io_in_b_0(b_850_0),
		.io_in_d_0(b_1874_0),
		.io_in_control_0_dataflow(mesh_18_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2898_0),
		.io_in_last_0(r_3922_0),
		.io_in_valid_0(r_1874_0),
		.io_out_a_0(_mesh_18_26_io_out_a_0),
		.io_out_c_0(_mesh_18_26_io_out_c_0),
		.io_out_b_0(_mesh_18_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_26_io_out_id_0),
		.io_out_last_0(_mesh_18_26_io_out_last_0),
		.io_out_valid_0(_mesh_18_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9973 == GlobalFiModInstNr[0]) || (9973 == GlobalFiModInstNr[1]) || (9973 == GlobalFiModInstNr[2]) || (9973 == GlobalFiModInstNr[3]))));
	Tile mesh_18_27(
		.clock(clock),
		.io_in_a_0(r_603_0),
		.io_in_b_0(b_882_0),
		.io_in_d_0(b_1906_0),
		.io_in_control_0_dataflow(mesh_18_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2930_0),
		.io_in_last_0(r_3954_0),
		.io_in_valid_0(r_1906_0),
		.io_out_a_0(_mesh_18_27_io_out_a_0),
		.io_out_c_0(_mesh_18_27_io_out_c_0),
		.io_out_b_0(_mesh_18_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_27_io_out_id_0),
		.io_out_last_0(_mesh_18_27_io_out_last_0),
		.io_out_valid_0(_mesh_18_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9974 == GlobalFiModInstNr[0]) || (9974 == GlobalFiModInstNr[1]) || (9974 == GlobalFiModInstNr[2]) || (9974 == GlobalFiModInstNr[3]))));
	Tile mesh_18_28(
		.clock(clock),
		.io_in_a_0(r_604_0),
		.io_in_b_0(b_914_0),
		.io_in_d_0(b_1938_0),
		.io_in_control_0_dataflow(mesh_18_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2962_0),
		.io_in_last_0(r_3986_0),
		.io_in_valid_0(r_1938_0),
		.io_out_a_0(_mesh_18_28_io_out_a_0),
		.io_out_c_0(_mesh_18_28_io_out_c_0),
		.io_out_b_0(_mesh_18_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_28_io_out_id_0),
		.io_out_last_0(_mesh_18_28_io_out_last_0),
		.io_out_valid_0(_mesh_18_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9975 == GlobalFiModInstNr[0]) || (9975 == GlobalFiModInstNr[1]) || (9975 == GlobalFiModInstNr[2]) || (9975 == GlobalFiModInstNr[3]))));
	Tile mesh_18_29(
		.clock(clock),
		.io_in_a_0(r_605_0),
		.io_in_b_0(b_946_0),
		.io_in_d_0(b_1970_0),
		.io_in_control_0_dataflow(mesh_18_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2994_0),
		.io_in_last_0(r_4018_0),
		.io_in_valid_0(r_1970_0),
		.io_out_a_0(_mesh_18_29_io_out_a_0),
		.io_out_c_0(_mesh_18_29_io_out_c_0),
		.io_out_b_0(_mesh_18_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_29_io_out_id_0),
		.io_out_last_0(_mesh_18_29_io_out_last_0),
		.io_out_valid_0(_mesh_18_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9976 == GlobalFiModInstNr[0]) || (9976 == GlobalFiModInstNr[1]) || (9976 == GlobalFiModInstNr[2]) || (9976 == GlobalFiModInstNr[3]))));
	Tile mesh_18_30(
		.clock(clock),
		.io_in_a_0(r_606_0),
		.io_in_b_0(b_978_0),
		.io_in_d_0(b_2002_0),
		.io_in_control_0_dataflow(mesh_18_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3026_0),
		.io_in_last_0(r_4050_0),
		.io_in_valid_0(r_2002_0),
		.io_out_a_0(_mesh_18_30_io_out_a_0),
		.io_out_c_0(_mesh_18_30_io_out_c_0),
		.io_out_b_0(_mesh_18_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_30_io_out_id_0),
		.io_out_last_0(_mesh_18_30_io_out_last_0),
		.io_out_valid_0(_mesh_18_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9977 == GlobalFiModInstNr[0]) || (9977 == GlobalFiModInstNr[1]) || (9977 == GlobalFiModInstNr[2]) || (9977 == GlobalFiModInstNr[3]))));
	Tile mesh_18_31(
		.clock(clock),
		.io_in_a_0(r_607_0),
		.io_in_b_0(b_1010_0),
		.io_in_d_0(b_2034_0),
		.io_in_control_0_dataflow(mesh_18_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_18_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_18_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3058_0),
		.io_in_last_0(r_4082_0),
		.io_in_valid_0(r_2034_0),
		.io_out_a_0(_mesh_18_31_io_out_a_0),
		.io_out_c_0(_mesh_18_31_io_out_c_0),
		.io_out_b_0(_mesh_18_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_18_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_18_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_18_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_18_31_io_out_id_0),
		.io_out_last_0(_mesh_18_31_io_out_last_0),
		.io_out_valid_0(_mesh_18_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9978 == GlobalFiModInstNr[0]) || (9978 == GlobalFiModInstNr[1]) || (9978 == GlobalFiModInstNr[2]) || (9978 == GlobalFiModInstNr[3]))));
	Tile mesh_19_0(
		.clock(clock),
		.io_in_a_0(r_608_0),
		.io_in_b_0(b_19_0),
		.io_in_d_0(b_1043_0),
		.io_in_control_0_dataflow(mesh_19_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2067_0),
		.io_in_last_0(r_3091_0),
		.io_in_valid_0(r_1043_0),
		.io_out_a_0(_mesh_19_0_io_out_a_0),
		.io_out_c_0(_mesh_19_0_io_out_c_0),
		.io_out_b_0(_mesh_19_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_0_io_out_id_0),
		.io_out_last_0(_mesh_19_0_io_out_last_0),
		.io_out_valid_0(_mesh_19_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9979 == GlobalFiModInstNr[0]) || (9979 == GlobalFiModInstNr[1]) || (9979 == GlobalFiModInstNr[2]) || (9979 == GlobalFiModInstNr[3]))));
	Tile mesh_19_1(
		.clock(clock),
		.io_in_a_0(r_609_0),
		.io_in_b_0(b_51_0),
		.io_in_d_0(b_1075_0),
		.io_in_control_0_dataflow(mesh_19_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2099_0),
		.io_in_last_0(r_3123_0),
		.io_in_valid_0(r_1075_0),
		.io_out_a_0(_mesh_19_1_io_out_a_0),
		.io_out_c_0(_mesh_19_1_io_out_c_0),
		.io_out_b_0(_mesh_19_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_1_io_out_id_0),
		.io_out_last_0(_mesh_19_1_io_out_last_0),
		.io_out_valid_0(_mesh_19_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9980 == GlobalFiModInstNr[0]) || (9980 == GlobalFiModInstNr[1]) || (9980 == GlobalFiModInstNr[2]) || (9980 == GlobalFiModInstNr[3]))));
	Tile mesh_19_2(
		.clock(clock),
		.io_in_a_0(r_610_0),
		.io_in_b_0(b_83_0),
		.io_in_d_0(b_1107_0),
		.io_in_control_0_dataflow(mesh_19_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2131_0),
		.io_in_last_0(r_3155_0),
		.io_in_valid_0(r_1107_0),
		.io_out_a_0(_mesh_19_2_io_out_a_0),
		.io_out_c_0(_mesh_19_2_io_out_c_0),
		.io_out_b_0(_mesh_19_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_2_io_out_id_0),
		.io_out_last_0(_mesh_19_2_io_out_last_0),
		.io_out_valid_0(_mesh_19_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9981 == GlobalFiModInstNr[0]) || (9981 == GlobalFiModInstNr[1]) || (9981 == GlobalFiModInstNr[2]) || (9981 == GlobalFiModInstNr[3]))));
	Tile mesh_19_3(
		.clock(clock),
		.io_in_a_0(r_611_0),
		.io_in_b_0(b_115_0),
		.io_in_d_0(b_1139_0),
		.io_in_control_0_dataflow(mesh_19_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2163_0),
		.io_in_last_0(r_3187_0),
		.io_in_valid_0(r_1139_0),
		.io_out_a_0(_mesh_19_3_io_out_a_0),
		.io_out_c_0(_mesh_19_3_io_out_c_0),
		.io_out_b_0(_mesh_19_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_3_io_out_id_0),
		.io_out_last_0(_mesh_19_3_io_out_last_0),
		.io_out_valid_0(_mesh_19_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9982 == GlobalFiModInstNr[0]) || (9982 == GlobalFiModInstNr[1]) || (9982 == GlobalFiModInstNr[2]) || (9982 == GlobalFiModInstNr[3]))));
	Tile mesh_19_4(
		.clock(clock),
		.io_in_a_0(r_612_0),
		.io_in_b_0(b_147_0),
		.io_in_d_0(b_1171_0),
		.io_in_control_0_dataflow(mesh_19_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2195_0),
		.io_in_last_0(r_3219_0),
		.io_in_valid_0(r_1171_0),
		.io_out_a_0(_mesh_19_4_io_out_a_0),
		.io_out_c_0(_mesh_19_4_io_out_c_0),
		.io_out_b_0(_mesh_19_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_4_io_out_id_0),
		.io_out_last_0(_mesh_19_4_io_out_last_0),
		.io_out_valid_0(_mesh_19_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9983 == GlobalFiModInstNr[0]) || (9983 == GlobalFiModInstNr[1]) || (9983 == GlobalFiModInstNr[2]) || (9983 == GlobalFiModInstNr[3]))));
	Tile mesh_19_5(
		.clock(clock),
		.io_in_a_0(r_613_0),
		.io_in_b_0(b_179_0),
		.io_in_d_0(b_1203_0),
		.io_in_control_0_dataflow(mesh_19_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2227_0),
		.io_in_last_0(r_3251_0),
		.io_in_valid_0(r_1203_0),
		.io_out_a_0(_mesh_19_5_io_out_a_0),
		.io_out_c_0(_mesh_19_5_io_out_c_0),
		.io_out_b_0(_mesh_19_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_5_io_out_id_0),
		.io_out_last_0(_mesh_19_5_io_out_last_0),
		.io_out_valid_0(_mesh_19_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9984 == GlobalFiModInstNr[0]) || (9984 == GlobalFiModInstNr[1]) || (9984 == GlobalFiModInstNr[2]) || (9984 == GlobalFiModInstNr[3]))));
	Tile mesh_19_6(
		.clock(clock),
		.io_in_a_0(r_614_0),
		.io_in_b_0(b_211_0),
		.io_in_d_0(b_1235_0),
		.io_in_control_0_dataflow(mesh_19_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2259_0),
		.io_in_last_0(r_3283_0),
		.io_in_valid_0(r_1235_0),
		.io_out_a_0(_mesh_19_6_io_out_a_0),
		.io_out_c_0(_mesh_19_6_io_out_c_0),
		.io_out_b_0(_mesh_19_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_6_io_out_id_0),
		.io_out_last_0(_mesh_19_6_io_out_last_0),
		.io_out_valid_0(_mesh_19_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9985 == GlobalFiModInstNr[0]) || (9985 == GlobalFiModInstNr[1]) || (9985 == GlobalFiModInstNr[2]) || (9985 == GlobalFiModInstNr[3]))));
	Tile mesh_19_7(
		.clock(clock),
		.io_in_a_0(r_615_0),
		.io_in_b_0(b_243_0),
		.io_in_d_0(b_1267_0),
		.io_in_control_0_dataflow(mesh_19_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2291_0),
		.io_in_last_0(r_3315_0),
		.io_in_valid_0(r_1267_0),
		.io_out_a_0(_mesh_19_7_io_out_a_0),
		.io_out_c_0(_mesh_19_7_io_out_c_0),
		.io_out_b_0(_mesh_19_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_7_io_out_id_0),
		.io_out_last_0(_mesh_19_7_io_out_last_0),
		.io_out_valid_0(_mesh_19_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9986 == GlobalFiModInstNr[0]) || (9986 == GlobalFiModInstNr[1]) || (9986 == GlobalFiModInstNr[2]) || (9986 == GlobalFiModInstNr[3]))));
	Tile mesh_19_8(
		.clock(clock),
		.io_in_a_0(r_616_0),
		.io_in_b_0(b_275_0),
		.io_in_d_0(b_1299_0),
		.io_in_control_0_dataflow(mesh_19_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2323_0),
		.io_in_last_0(r_3347_0),
		.io_in_valid_0(r_1299_0),
		.io_out_a_0(_mesh_19_8_io_out_a_0),
		.io_out_c_0(_mesh_19_8_io_out_c_0),
		.io_out_b_0(_mesh_19_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_8_io_out_id_0),
		.io_out_last_0(_mesh_19_8_io_out_last_0),
		.io_out_valid_0(_mesh_19_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9987 == GlobalFiModInstNr[0]) || (9987 == GlobalFiModInstNr[1]) || (9987 == GlobalFiModInstNr[2]) || (9987 == GlobalFiModInstNr[3]))));
	Tile mesh_19_9(
		.clock(clock),
		.io_in_a_0(r_617_0),
		.io_in_b_0(b_307_0),
		.io_in_d_0(b_1331_0),
		.io_in_control_0_dataflow(mesh_19_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2355_0),
		.io_in_last_0(r_3379_0),
		.io_in_valid_0(r_1331_0),
		.io_out_a_0(_mesh_19_9_io_out_a_0),
		.io_out_c_0(_mesh_19_9_io_out_c_0),
		.io_out_b_0(_mesh_19_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_9_io_out_id_0),
		.io_out_last_0(_mesh_19_9_io_out_last_0),
		.io_out_valid_0(_mesh_19_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9988 == GlobalFiModInstNr[0]) || (9988 == GlobalFiModInstNr[1]) || (9988 == GlobalFiModInstNr[2]) || (9988 == GlobalFiModInstNr[3]))));
	Tile mesh_19_10(
		.clock(clock),
		.io_in_a_0(r_618_0),
		.io_in_b_0(b_339_0),
		.io_in_d_0(b_1363_0),
		.io_in_control_0_dataflow(mesh_19_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2387_0),
		.io_in_last_0(r_3411_0),
		.io_in_valid_0(r_1363_0),
		.io_out_a_0(_mesh_19_10_io_out_a_0),
		.io_out_c_0(_mesh_19_10_io_out_c_0),
		.io_out_b_0(_mesh_19_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_10_io_out_id_0),
		.io_out_last_0(_mesh_19_10_io_out_last_0),
		.io_out_valid_0(_mesh_19_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9989 == GlobalFiModInstNr[0]) || (9989 == GlobalFiModInstNr[1]) || (9989 == GlobalFiModInstNr[2]) || (9989 == GlobalFiModInstNr[3]))));
	Tile mesh_19_11(
		.clock(clock),
		.io_in_a_0(r_619_0),
		.io_in_b_0(b_371_0),
		.io_in_d_0(b_1395_0),
		.io_in_control_0_dataflow(mesh_19_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2419_0),
		.io_in_last_0(r_3443_0),
		.io_in_valid_0(r_1395_0),
		.io_out_a_0(_mesh_19_11_io_out_a_0),
		.io_out_c_0(_mesh_19_11_io_out_c_0),
		.io_out_b_0(_mesh_19_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_11_io_out_id_0),
		.io_out_last_0(_mesh_19_11_io_out_last_0),
		.io_out_valid_0(_mesh_19_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9990 == GlobalFiModInstNr[0]) || (9990 == GlobalFiModInstNr[1]) || (9990 == GlobalFiModInstNr[2]) || (9990 == GlobalFiModInstNr[3]))));
	Tile mesh_19_12(
		.clock(clock),
		.io_in_a_0(r_620_0),
		.io_in_b_0(b_403_0),
		.io_in_d_0(b_1427_0),
		.io_in_control_0_dataflow(mesh_19_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2451_0),
		.io_in_last_0(r_3475_0),
		.io_in_valid_0(r_1427_0),
		.io_out_a_0(_mesh_19_12_io_out_a_0),
		.io_out_c_0(_mesh_19_12_io_out_c_0),
		.io_out_b_0(_mesh_19_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_12_io_out_id_0),
		.io_out_last_0(_mesh_19_12_io_out_last_0),
		.io_out_valid_0(_mesh_19_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9991 == GlobalFiModInstNr[0]) || (9991 == GlobalFiModInstNr[1]) || (9991 == GlobalFiModInstNr[2]) || (9991 == GlobalFiModInstNr[3]))));
	Tile mesh_19_13(
		.clock(clock),
		.io_in_a_0(r_621_0),
		.io_in_b_0(b_435_0),
		.io_in_d_0(b_1459_0),
		.io_in_control_0_dataflow(mesh_19_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2483_0),
		.io_in_last_0(r_3507_0),
		.io_in_valid_0(r_1459_0),
		.io_out_a_0(_mesh_19_13_io_out_a_0),
		.io_out_c_0(_mesh_19_13_io_out_c_0),
		.io_out_b_0(_mesh_19_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_13_io_out_id_0),
		.io_out_last_0(_mesh_19_13_io_out_last_0),
		.io_out_valid_0(_mesh_19_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9992 == GlobalFiModInstNr[0]) || (9992 == GlobalFiModInstNr[1]) || (9992 == GlobalFiModInstNr[2]) || (9992 == GlobalFiModInstNr[3]))));
	Tile mesh_19_14(
		.clock(clock),
		.io_in_a_0(r_622_0),
		.io_in_b_0(b_467_0),
		.io_in_d_0(b_1491_0),
		.io_in_control_0_dataflow(mesh_19_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2515_0),
		.io_in_last_0(r_3539_0),
		.io_in_valid_0(r_1491_0),
		.io_out_a_0(_mesh_19_14_io_out_a_0),
		.io_out_c_0(_mesh_19_14_io_out_c_0),
		.io_out_b_0(_mesh_19_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_14_io_out_id_0),
		.io_out_last_0(_mesh_19_14_io_out_last_0),
		.io_out_valid_0(_mesh_19_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9993 == GlobalFiModInstNr[0]) || (9993 == GlobalFiModInstNr[1]) || (9993 == GlobalFiModInstNr[2]) || (9993 == GlobalFiModInstNr[3]))));
	Tile mesh_19_15(
		.clock(clock),
		.io_in_a_0(r_623_0),
		.io_in_b_0(b_499_0),
		.io_in_d_0(b_1523_0),
		.io_in_control_0_dataflow(mesh_19_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2547_0),
		.io_in_last_0(r_3571_0),
		.io_in_valid_0(r_1523_0),
		.io_out_a_0(_mesh_19_15_io_out_a_0),
		.io_out_c_0(_mesh_19_15_io_out_c_0),
		.io_out_b_0(_mesh_19_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_15_io_out_id_0),
		.io_out_last_0(_mesh_19_15_io_out_last_0),
		.io_out_valid_0(_mesh_19_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9994 == GlobalFiModInstNr[0]) || (9994 == GlobalFiModInstNr[1]) || (9994 == GlobalFiModInstNr[2]) || (9994 == GlobalFiModInstNr[3]))));
	Tile mesh_19_16(
		.clock(clock),
		.io_in_a_0(r_624_0),
		.io_in_b_0(b_531_0),
		.io_in_d_0(b_1555_0),
		.io_in_control_0_dataflow(mesh_19_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2579_0),
		.io_in_last_0(r_3603_0),
		.io_in_valid_0(r_1555_0),
		.io_out_a_0(_mesh_19_16_io_out_a_0),
		.io_out_c_0(_mesh_19_16_io_out_c_0),
		.io_out_b_0(_mesh_19_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_16_io_out_id_0),
		.io_out_last_0(_mesh_19_16_io_out_last_0),
		.io_out_valid_0(_mesh_19_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9995 == GlobalFiModInstNr[0]) || (9995 == GlobalFiModInstNr[1]) || (9995 == GlobalFiModInstNr[2]) || (9995 == GlobalFiModInstNr[3]))));
	Tile mesh_19_17(
		.clock(clock),
		.io_in_a_0(r_625_0),
		.io_in_b_0(b_563_0),
		.io_in_d_0(b_1587_0),
		.io_in_control_0_dataflow(mesh_19_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2611_0),
		.io_in_last_0(r_3635_0),
		.io_in_valid_0(r_1587_0),
		.io_out_a_0(_mesh_19_17_io_out_a_0),
		.io_out_c_0(_mesh_19_17_io_out_c_0),
		.io_out_b_0(_mesh_19_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_17_io_out_id_0),
		.io_out_last_0(_mesh_19_17_io_out_last_0),
		.io_out_valid_0(_mesh_19_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9996 == GlobalFiModInstNr[0]) || (9996 == GlobalFiModInstNr[1]) || (9996 == GlobalFiModInstNr[2]) || (9996 == GlobalFiModInstNr[3]))));
	Tile mesh_19_18(
		.clock(clock),
		.io_in_a_0(r_626_0),
		.io_in_b_0(b_595_0),
		.io_in_d_0(b_1619_0),
		.io_in_control_0_dataflow(mesh_19_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2643_0),
		.io_in_last_0(r_3667_0),
		.io_in_valid_0(r_1619_0),
		.io_out_a_0(_mesh_19_18_io_out_a_0),
		.io_out_c_0(_mesh_19_18_io_out_c_0),
		.io_out_b_0(_mesh_19_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_18_io_out_id_0),
		.io_out_last_0(_mesh_19_18_io_out_last_0),
		.io_out_valid_0(_mesh_19_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9997 == GlobalFiModInstNr[0]) || (9997 == GlobalFiModInstNr[1]) || (9997 == GlobalFiModInstNr[2]) || (9997 == GlobalFiModInstNr[3]))));
	Tile mesh_19_19(
		.clock(clock),
		.io_in_a_0(r_627_0),
		.io_in_b_0(b_627_0),
		.io_in_d_0(b_1651_0),
		.io_in_control_0_dataflow(mesh_19_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2675_0),
		.io_in_last_0(r_3699_0),
		.io_in_valid_0(r_1651_0),
		.io_out_a_0(_mesh_19_19_io_out_a_0),
		.io_out_c_0(_mesh_19_19_io_out_c_0),
		.io_out_b_0(_mesh_19_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_19_io_out_id_0),
		.io_out_last_0(_mesh_19_19_io_out_last_0),
		.io_out_valid_0(_mesh_19_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9998 == GlobalFiModInstNr[0]) || (9998 == GlobalFiModInstNr[1]) || (9998 == GlobalFiModInstNr[2]) || (9998 == GlobalFiModInstNr[3]))));
	Tile mesh_19_20(
		.clock(clock),
		.io_in_a_0(r_628_0),
		.io_in_b_0(b_659_0),
		.io_in_d_0(b_1683_0),
		.io_in_control_0_dataflow(mesh_19_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2707_0),
		.io_in_last_0(r_3731_0),
		.io_in_valid_0(r_1683_0),
		.io_out_a_0(_mesh_19_20_io_out_a_0),
		.io_out_c_0(_mesh_19_20_io_out_c_0),
		.io_out_b_0(_mesh_19_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_20_io_out_id_0),
		.io_out_last_0(_mesh_19_20_io_out_last_0),
		.io_out_valid_0(_mesh_19_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((9999 == GlobalFiModInstNr[0]) || (9999 == GlobalFiModInstNr[1]) || (9999 == GlobalFiModInstNr[2]) || (9999 == GlobalFiModInstNr[3]))));
	Tile mesh_19_21(
		.clock(clock),
		.io_in_a_0(r_629_0),
		.io_in_b_0(b_691_0),
		.io_in_d_0(b_1715_0),
		.io_in_control_0_dataflow(mesh_19_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2739_0),
		.io_in_last_0(r_3763_0),
		.io_in_valid_0(r_1715_0),
		.io_out_a_0(_mesh_19_21_io_out_a_0),
		.io_out_c_0(_mesh_19_21_io_out_c_0),
		.io_out_b_0(_mesh_19_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_21_io_out_id_0),
		.io_out_last_0(_mesh_19_21_io_out_last_0),
		.io_out_valid_0(_mesh_19_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10000 == GlobalFiModInstNr[0]) || (10000 == GlobalFiModInstNr[1]) || (10000 == GlobalFiModInstNr[2]) || (10000 == GlobalFiModInstNr[3]))));
	Tile mesh_19_22(
		.clock(clock),
		.io_in_a_0(r_630_0),
		.io_in_b_0(b_723_0),
		.io_in_d_0(b_1747_0),
		.io_in_control_0_dataflow(mesh_19_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2771_0),
		.io_in_last_0(r_3795_0),
		.io_in_valid_0(r_1747_0),
		.io_out_a_0(_mesh_19_22_io_out_a_0),
		.io_out_c_0(_mesh_19_22_io_out_c_0),
		.io_out_b_0(_mesh_19_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_22_io_out_id_0),
		.io_out_last_0(_mesh_19_22_io_out_last_0),
		.io_out_valid_0(_mesh_19_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10001 == GlobalFiModInstNr[0]) || (10001 == GlobalFiModInstNr[1]) || (10001 == GlobalFiModInstNr[2]) || (10001 == GlobalFiModInstNr[3]))));
	Tile mesh_19_23(
		.clock(clock),
		.io_in_a_0(r_631_0),
		.io_in_b_0(b_755_0),
		.io_in_d_0(b_1779_0),
		.io_in_control_0_dataflow(mesh_19_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2803_0),
		.io_in_last_0(r_3827_0),
		.io_in_valid_0(r_1779_0),
		.io_out_a_0(_mesh_19_23_io_out_a_0),
		.io_out_c_0(_mesh_19_23_io_out_c_0),
		.io_out_b_0(_mesh_19_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_23_io_out_id_0),
		.io_out_last_0(_mesh_19_23_io_out_last_0),
		.io_out_valid_0(_mesh_19_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10002 == GlobalFiModInstNr[0]) || (10002 == GlobalFiModInstNr[1]) || (10002 == GlobalFiModInstNr[2]) || (10002 == GlobalFiModInstNr[3]))));
	Tile mesh_19_24(
		.clock(clock),
		.io_in_a_0(r_632_0),
		.io_in_b_0(b_787_0),
		.io_in_d_0(b_1811_0),
		.io_in_control_0_dataflow(mesh_19_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2835_0),
		.io_in_last_0(r_3859_0),
		.io_in_valid_0(r_1811_0),
		.io_out_a_0(_mesh_19_24_io_out_a_0),
		.io_out_c_0(_mesh_19_24_io_out_c_0),
		.io_out_b_0(_mesh_19_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_24_io_out_id_0),
		.io_out_last_0(_mesh_19_24_io_out_last_0),
		.io_out_valid_0(_mesh_19_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10003 == GlobalFiModInstNr[0]) || (10003 == GlobalFiModInstNr[1]) || (10003 == GlobalFiModInstNr[2]) || (10003 == GlobalFiModInstNr[3]))));
	Tile mesh_19_25(
		.clock(clock),
		.io_in_a_0(r_633_0),
		.io_in_b_0(b_819_0),
		.io_in_d_0(b_1843_0),
		.io_in_control_0_dataflow(mesh_19_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2867_0),
		.io_in_last_0(r_3891_0),
		.io_in_valid_0(r_1843_0),
		.io_out_a_0(_mesh_19_25_io_out_a_0),
		.io_out_c_0(_mesh_19_25_io_out_c_0),
		.io_out_b_0(_mesh_19_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_25_io_out_id_0),
		.io_out_last_0(_mesh_19_25_io_out_last_0),
		.io_out_valid_0(_mesh_19_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10004 == GlobalFiModInstNr[0]) || (10004 == GlobalFiModInstNr[1]) || (10004 == GlobalFiModInstNr[2]) || (10004 == GlobalFiModInstNr[3]))));
	Tile mesh_19_26(
		.clock(clock),
		.io_in_a_0(r_634_0),
		.io_in_b_0(b_851_0),
		.io_in_d_0(b_1875_0),
		.io_in_control_0_dataflow(mesh_19_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2899_0),
		.io_in_last_0(r_3923_0),
		.io_in_valid_0(r_1875_0),
		.io_out_a_0(_mesh_19_26_io_out_a_0),
		.io_out_c_0(_mesh_19_26_io_out_c_0),
		.io_out_b_0(_mesh_19_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_26_io_out_id_0),
		.io_out_last_0(_mesh_19_26_io_out_last_0),
		.io_out_valid_0(_mesh_19_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10005 == GlobalFiModInstNr[0]) || (10005 == GlobalFiModInstNr[1]) || (10005 == GlobalFiModInstNr[2]) || (10005 == GlobalFiModInstNr[3]))));
	Tile mesh_19_27(
		.clock(clock),
		.io_in_a_0(r_635_0),
		.io_in_b_0(b_883_0),
		.io_in_d_0(b_1907_0),
		.io_in_control_0_dataflow(mesh_19_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2931_0),
		.io_in_last_0(r_3955_0),
		.io_in_valid_0(r_1907_0),
		.io_out_a_0(_mesh_19_27_io_out_a_0),
		.io_out_c_0(_mesh_19_27_io_out_c_0),
		.io_out_b_0(_mesh_19_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_27_io_out_id_0),
		.io_out_last_0(_mesh_19_27_io_out_last_0),
		.io_out_valid_0(_mesh_19_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10006 == GlobalFiModInstNr[0]) || (10006 == GlobalFiModInstNr[1]) || (10006 == GlobalFiModInstNr[2]) || (10006 == GlobalFiModInstNr[3]))));
	Tile mesh_19_28(
		.clock(clock),
		.io_in_a_0(r_636_0),
		.io_in_b_0(b_915_0),
		.io_in_d_0(b_1939_0),
		.io_in_control_0_dataflow(mesh_19_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2963_0),
		.io_in_last_0(r_3987_0),
		.io_in_valid_0(r_1939_0),
		.io_out_a_0(_mesh_19_28_io_out_a_0),
		.io_out_c_0(_mesh_19_28_io_out_c_0),
		.io_out_b_0(_mesh_19_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_28_io_out_id_0),
		.io_out_last_0(_mesh_19_28_io_out_last_0),
		.io_out_valid_0(_mesh_19_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10007 == GlobalFiModInstNr[0]) || (10007 == GlobalFiModInstNr[1]) || (10007 == GlobalFiModInstNr[2]) || (10007 == GlobalFiModInstNr[3]))));
	Tile mesh_19_29(
		.clock(clock),
		.io_in_a_0(r_637_0),
		.io_in_b_0(b_947_0),
		.io_in_d_0(b_1971_0),
		.io_in_control_0_dataflow(mesh_19_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2995_0),
		.io_in_last_0(r_4019_0),
		.io_in_valid_0(r_1971_0),
		.io_out_a_0(_mesh_19_29_io_out_a_0),
		.io_out_c_0(_mesh_19_29_io_out_c_0),
		.io_out_b_0(_mesh_19_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_29_io_out_id_0),
		.io_out_last_0(_mesh_19_29_io_out_last_0),
		.io_out_valid_0(_mesh_19_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10008 == GlobalFiModInstNr[0]) || (10008 == GlobalFiModInstNr[1]) || (10008 == GlobalFiModInstNr[2]) || (10008 == GlobalFiModInstNr[3]))));
	Tile mesh_19_30(
		.clock(clock),
		.io_in_a_0(r_638_0),
		.io_in_b_0(b_979_0),
		.io_in_d_0(b_2003_0),
		.io_in_control_0_dataflow(mesh_19_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3027_0),
		.io_in_last_0(r_4051_0),
		.io_in_valid_0(r_2003_0),
		.io_out_a_0(_mesh_19_30_io_out_a_0),
		.io_out_c_0(_mesh_19_30_io_out_c_0),
		.io_out_b_0(_mesh_19_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_30_io_out_id_0),
		.io_out_last_0(_mesh_19_30_io_out_last_0),
		.io_out_valid_0(_mesh_19_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10009 == GlobalFiModInstNr[0]) || (10009 == GlobalFiModInstNr[1]) || (10009 == GlobalFiModInstNr[2]) || (10009 == GlobalFiModInstNr[3]))));
	Tile mesh_19_31(
		.clock(clock),
		.io_in_a_0(r_639_0),
		.io_in_b_0(b_1011_0),
		.io_in_d_0(b_2035_0),
		.io_in_control_0_dataflow(mesh_19_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_19_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_19_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3059_0),
		.io_in_last_0(r_4083_0),
		.io_in_valid_0(r_2035_0),
		.io_out_a_0(_mesh_19_31_io_out_a_0),
		.io_out_c_0(_mesh_19_31_io_out_c_0),
		.io_out_b_0(_mesh_19_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_19_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_19_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_19_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_19_31_io_out_id_0),
		.io_out_last_0(_mesh_19_31_io_out_last_0),
		.io_out_valid_0(_mesh_19_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10010 == GlobalFiModInstNr[0]) || (10010 == GlobalFiModInstNr[1]) || (10010 == GlobalFiModInstNr[2]) || (10010 == GlobalFiModInstNr[3]))));
	Tile mesh_20_0(
		.clock(clock),
		.io_in_a_0(r_640_0),
		.io_in_b_0(b_20_0),
		.io_in_d_0(b_1044_0),
		.io_in_control_0_dataflow(mesh_20_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2068_0),
		.io_in_last_0(r_3092_0),
		.io_in_valid_0(r_1044_0),
		.io_out_a_0(_mesh_20_0_io_out_a_0),
		.io_out_c_0(_mesh_20_0_io_out_c_0),
		.io_out_b_0(_mesh_20_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_0_io_out_id_0),
		.io_out_last_0(_mesh_20_0_io_out_last_0),
		.io_out_valid_0(_mesh_20_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10011 == GlobalFiModInstNr[0]) || (10011 == GlobalFiModInstNr[1]) || (10011 == GlobalFiModInstNr[2]) || (10011 == GlobalFiModInstNr[3]))));
	Tile mesh_20_1(
		.clock(clock),
		.io_in_a_0(r_641_0),
		.io_in_b_0(b_52_0),
		.io_in_d_0(b_1076_0),
		.io_in_control_0_dataflow(mesh_20_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2100_0),
		.io_in_last_0(r_3124_0),
		.io_in_valid_0(r_1076_0),
		.io_out_a_0(_mesh_20_1_io_out_a_0),
		.io_out_c_0(_mesh_20_1_io_out_c_0),
		.io_out_b_0(_mesh_20_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_1_io_out_id_0),
		.io_out_last_0(_mesh_20_1_io_out_last_0),
		.io_out_valid_0(_mesh_20_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10012 == GlobalFiModInstNr[0]) || (10012 == GlobalFiModInstNr[1]) || (10012 == GlobalFiModInstNr[2]) || (10012 == GlobalFiModInstNr[3]))));
	Tile mesh_20_2(
		.clock(clock),
		.io_in_a_0(r_642_0),
		.io_in_b_0(b_84_0),
		.io_in_d_0(b_1108_0),
		.io_in_control_0_dataflow(mesh_20_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2132_0),
		.io_in_last_0(r_3156_0),
		.io_in_valid_0(r_1108_0),
		.io_out_a_0(_mesh_20_2_io_out_a_0),
		.io_out_c_0(_mesh_20_2_io_out_c_0),
		.io_out_b_0(_mesh_20_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_2_io_out_id_0),
		.io_out_last_0(_mesh_20_2_io_out_last_0),
		.io_out_valid_0(_mesh_20_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10013 == GlobalFiModInstNr[0]) || (10013 == GlobalFiModInstNr[1]) || (10013 == GlobalFiModInstNr[2]) || (10013 == GlobalFiModInstNr[3]))));
	Tile mesh_20_3(
		.clock(clock),
		.io_in_a_0(r_643_0),
		.io_in_b_0(b_116_0),
		.io_in_d_0(b_1140_0),
		.io_in_control_0_dataflow(mesh_20_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2164_0),
		.io_in_last_0(r_3188_0),
		.io_in_valid_0(r_1140_0),
		.io_out_a_0(_mesh_20_3_io_out_a_0),
		.io_out_c_0(_mesh_20_3_io_out_c_0),
		.io_out_b_0(_mesh_20_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_3_io_out_id_0),
		.io_out_last_0(_mesh_20_3_io_out_last_0),
		.io_out_valid_0(_mesh_20_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10014 == GlobalFiModInstNr[0]) || (10014 == GlobalFiModInstNr[1]) || (10014 == GlobalFiModInstNr[2]) || (10014 == GlobalFiModInstNr[3]))));
	Tile mesh_20_4(
		.clock(clock),
		.io_in_a_0(r_644_0),
		.io_in_b_0(b_148_0),
		.io_in_d_0(b_1172_0),
		.io_in_control_0_dataflow(mesh_20_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2196_0),
		.io_in_last_0(r_3220_0),
		.io_in_valid_0(r_1172_0),
		.io_out_a_0(_mesh_20_4_io_out_a_0),
		.io_out_c_0(_mesh_20_4_io_out_c_0),
		.io_out_b_0(_mesh_20_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_4_io_out_id_0),
		.io_out_last_0(_mesh_20_4_io_out_last_0),
		.io_out_valid_0(_mesh_20_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10015 == GlobalFiModInstNr[0]) || (10015 == GlobalFiModInstNr[1]) || (10015 == GlobalFiModInstNr[2]) || (10015 == GlobalFiModInstNr[3]))));
	Tile mesh_20_5(
		.clock(clock),
		.io_in_a_0(r_645_0),
		.io_in_b_0(b_180_0),
		.io_in_d_0(b_1204_0),
		.io_in_control_0_dataflow(mesh_20_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2228_0),
		.io_in_last_0(r_3252_0),
		.io_in_valid_0(r_1204_0),
		.io_out_a_0(_mesh_20_5_io_out_a_0),
		.io_out_c_0(_mesh_20_5_io_out_c_0),
		.io_out_b_0(_mesh_20_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_5_io_out_id_0),
		.io_out_last_0(_mesh_20_5_io_out_last_0),
		.io_out_valid_0(_mesh_20_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10016 == GlobalFiModInstNr[0]) || (10016 == GlobalFiModInstNr[1]) || (10016 == GlobalFiModInstNr[2]) || (10016 == GlobalFiModInstNr[3]))));
	Tile mesh_20_6(
		.clock(clock),
		.io_in_a_0(r_646_0),
		.io_in_b_0(b_212_0),
		.io_in_d_0(b_1236_0),
		.io_in_control_0_dataflow(mesh_20_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2260_0),
		.io_in_last_0(r_3284_0),
		.io_in_valid_0(r_1236_0),
		.io_out_a_0(_mesh_20_6_io_out_a_0),
		.io_out_c_0(_mesh_20_6_io_out_c_0),
		.io_out_b_0(_mesh_20_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_6_io_out_id_0),
		.io_out_last_0(_mesh_20_6_io_out_last_0),
		.io_out_valid_0(_mesh_20_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10017 == GlobalFiModInstNr[0]) || (10017 == GlobalFiModInstNr[1]) || (10017 == GlobalFiModInstNr[2]) || (10017 == GlobalFiModInstNr[3]))));
	Tile mesh_20_7(
		.clock(clock),
		.io_in_a_0(r_647_0),
		.io_in_b_0(b_244_0),
		.io_in_d_0(b_1268_0),
		.io_in_control_0_dataflow(mesh_20_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2292_0),
		.io_in_last_0(r_3316_0),
		.io_in_valid_0(r_1268_0),
		.io_out_a_0(_mesh_20_7_io_out_a_0),
		.io_out_c_0(_mesh_20_7_io_out_c_0),
		.io_out_b_0(_mesh_20_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_7_io_out_id_0),
		.io_out_last_0(_mesh_20_7_io_out_last_0),
		.io_out_valid_0(_mesh_20_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10018 == GlobalFiModInstNr[0]) || (10018 == GlobalFiModInstNr[1]) || (10018 == GlobalFiModInstNr[2]) || (10018 == GlobalFiModInstNr[3]))));
	Tile mesh_20_8(
		.clock(clock),
		.io_in_a_0(r_648_0),
		.io_in_b_0(b_276_0),
		.io_in_d_0(b_1300_0),
		.io_in_control_0_dataflow(mesh_20_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2324_0),
		.io_in_last_0(r_3348_0),
		.io_in_valid_0(r_1300_0),
		.io_out_a_0(_mesh_20_8_io_out_a_0),
		.io_out_c_0(_mesh_20_8_io_out_c_0),
		.io_out_b_0(_mesh_20_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_8_io_out_id_0),
		.io_out_last_0(_mesh_20_8_io_out_last_0),
		.io_out_valid_0(_mesh_20_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10019 == GlobalFiModInstNr[0]) || (10019 == GlobalFiModInstNr[1]) || (10019 == GlobalFiModInstNr[2]) || (10019 == GlobalFiModInstNr[3]))));
	Tile mesh_20_9(
		.clock(clock),
		.io_in_a_0(r_649_0),
		.io_in_b_0(b_308_0),
		.io_in_d_0(b_1332_0),
		.io_in_control_0_dataflow(mesh_20_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2356_0),
		.io_in_last_0(r_3380_0),
		.io_in_valid_0(r_1332_0),
		.io_out_a_0(_mesh_20_9_io_out_a_0),
		.io_out_c_0(_mesh_20_9_io_out_c_0),
		.io_out_b_0(_mesh_20_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_9_io_out_id_0),
		.io_out_last_0(_mesh_20_9_io_out_last_0),
		.io_out_valid_0(_mesh_20_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10020 == GlobalFiModInstNr[0]) || (10020 == GlobalFiModInstNr[1]) || (10020 == GlobalFiModInstNr[2]) || (10020 == GlobalFiModInstNr[3]))));
	Tile mesh_20_10(
		.clock(clock),
		.io_in_a_0(r_650_0),
		.io_in_b_0(b_340_0),
		.io_in_d_0(b_1364_0),
		.io_in_control_0_dataflow(mesh_20_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2388_0),
		.io_in_last_0(r_3412_0),
		.io_in_valid_0(r_1364_0),
		.io_out_a_0(_mesh_20_10_io_out_a_0),
		.io_out_c_0(_mesh_20_10_io_out_c_0),
		.io_out_b_0(_mesh_20_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_10_io_out_id_0),
		.io_out_last_0(_mesh_20_10_io_out_last_0),
		.io_out_valid_0(_mesh_20_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10021 == GlobalFiModInstNr[0]) || (10021 == GlobalFiModInstNr[1]) || (10021 == GlobalFiModInstNr[2]) || (10021 == GlobalFiModInstNr[3]))));
	Tile mesh_20_11(
		.clock(clock),
		.io_in_a_0(r_651_0),
		.io_in_b_0(b_372_0),
		.io_in_d_0(b_1396_0),
		.io_in_control_0_dataflow(mesh_20_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2420_0),
		.io_in_last_0(r_3444_0),
		.io_in_valid_0(r_1396_0),
		.io_out_a_0(_mesh_20_11_io_out_a_0),
		.io_out_c_0(_mesh_20_11_io_out_c_0),
		.io_out_b_0(_mesh_20_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_11_io_out_id_0),
		.io_out_last_0(_mesh_20_11_io_out_last_0),
		.io_out_valid_0(_mesh_20_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10022 == GlobalFiModInstNr[0]) || (10022 == GlobalFiModInstNr[1]) || (10022 == GlobalFiModInstNr[2]) || (10022 == GlobalFiModInstNr[3]))));
	Tile mesh_20_12(
		.clock(clock),
		.io_in_a_0(r_652_0),
		.io_in_b_0(b_404_0),
		.io_in_d_0(b_1428_0),
		.io_in_control_0_dataflow(mesh_20_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2452_0),
		.io_in_last_0(r_3476_0),
		.io_in_valid_0(r_1428_0),
		.io_out_a_0(_mesh_20_12_io_out_a_0),
		.io_out_c_0(_mesh_20_12_io_out_c_0),
		.io_out_b_0(_mesh_20_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_12_io_out_id_0),
		.io_out_last_0(_mesh_20_12_io_out_last_0),
		.io_out_valid_0(_mesh_20_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10023 == GlobalFiModInstNr[0]) || (10023 == GlobalFiModInstNr[1]) || (10023 == GlobalFiModInstNr[2]) || (10023 == GlobalFiModInstNr[3]))));
	Tile mesh_20_13(
		.clock(clock),
		.io_in_a_0(r_653_0),
		.io_in_b_0(b_436_0),
		.io_in_d_0(b_1460_0),
		.io_in_control_0_dataflow(mesh_20_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2484_0),
		.io_in_last_0(r_3508_0),
		.io_in_valid_0(r_1460_0),
		.io_out_a_0(_mesh_20_13_io_out_a_0),
		.io_out_c_0(_mesh_20_13_io_out_c_0),
		.io_out_b_0(_mesh_20_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_13_io_out_id_0),
		.io_out_last_0(_mesh_20_13_io_out_last_0),
		.io_out_valid_0(_mesh_20_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10024 == GlobalFiModInstNr[0]) || (10024 == GlobalFiModInstNr[1]) || (10024 == GlobalFiModInstNr[2]) || (10024 == GlobalFiModInstNr[3]))));
	Tile mesh_20_14(
		.clock(clock),
		.io_in_a_0(r_654_0),
		.io_in_b_0(b_468_0),
		.io_in_d_0(b_1492_0),
		.io_in_control_0_dataflow(mesh_20_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2516_0),
		.io_in_last_0(r_3540_0),
		.io_in_valid_0(r_1492_0),
		.io_out_a_0(_mesh_20_14_io_out_a_0),
		.io_out_c_0(_mesh_20_14_io_out_c_0),
		.io_out_b_0(_mesh_20_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_14_io_out_id_0),
		.io_out_last_0(_mesh_20_14_io_out_last_0),
		.io_out_valid_0(_mesh_20_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10025 == GlobalFiModInstNr[0]) || (10025 == GlobalFiModInstNr[1]) || (10025 == GlobalFiModInstNr[2]) || (10025 == GlobalFiModInstNr[3]))));
	Tile mesh_20_15(
		.clock(clock),
		.io_in_a_0(r_655_0),
		.io_in_b_0(b_500_0),
		.io_in_d_0(b_1524_0),
		.io_in_control_0_dataflow(mesh_20_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2548_0),
		.io_in_last_0(r_3572_0),
		.io_in_valid_0(r_1524_0),
		.io_out_a_0(_mesh_20_15_io_out_a_0),
		.io_out_c_0(_mesh_20_15_io_out_c_0),
		.io_out_b_0(_mesh_20_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_15_io_out_id_0),
		.io_out_last_0(_mesh_20_15_io_out_last_0),
		.io_out_valid_0(_mesh_20_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10026 == GlobalFiModInstNr[0]) || (10026 == GlobalFiModInstNr[1]) || (10026 == GlobalFiModInstNr[2]) || (10026 == GlobalFiModInstNr[3]))));
	Tile mesh_20_16(
		.clock(clock),
		.io_in_a_0(r_656_0),
		.io_in_b_0(b_532_0),
		.io_in_d_0(b_1556_0),
		.io_in_control_0_dataflow(mesh_20_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2580_0),
		.io_in_last_0(r_3604_0),
		.io_in_valid_0(r_1556_0),
		.io_out_a_0(_mesh_20_16_io_out_a_0),
		.io_out_c_0(_mesh_20_16_io_out_c_0),
		.io_out_b_0(_mesh_20_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_16_io_out_id_0),
		.io_out_last_0(_mesh_20_16_io_out_last_0),
		.io_out_valid_0(_mesh_20_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10027 == GlobalFiModInstNr[0]) || (10027 == GlobalFiModInstNr[1]) || (10027 == GlobalFiModInstNr[2]) || (10027 == GlobalFiModInstNr[3]))));
	Tile mesh_20_17(
		.clock(clock),
		.io_in_a_0(r_657_0),
		.io_in_b_0(b_564_0),
		.io_in_d_0(b_1588_0),
		.io_in_control_0_dataflow(mesh_20_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2612_0),
		.io_in_last_0(r_3636_0),
		.io_in_valid_0(r_1588_0),
		.io_out_a_0(_mesh_20_17_io_out_a_0),
		.io_out_c_0(_mesh_20_17_io_out_c_0),
		.io_out_b_0(_mesh_20_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_17_io_out_id_0),
		.io_out_last_0(_mesh_20_17_io_out_last_0),
		.io_out_valid_0(_mesh_20_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10028 == GlobalFiModInstNr[0]) || (10028 == GlobalFiModInstNr[1]) || (10028 == GlobalFiModInstNr[2]) || (10028 == GlobalFiModInstNr[3]))));
	Tile mesh_20_18(
		.clock(clock),
		.io_in_a_0(r_658_0),
		.io_in_b_0(b_596_0),
		.io_in_d_0(b_1620_0),
		.io_in_control_0_dataflow(mesh_20_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2644_0),
		.io_in_last_0(r_3668_0),
		.io_in_valid_0(r_1620_0),
		.io_out_a_0(_mesh_20_18_io_out_a_0),
		.io_out_c_0(_mesh_20_18_io_out_c_0),
		.io_out_b_0(_mesh_20_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_18_io_out_id_0),
		.io_out_last_0(_mesh_20_18_io_out_last_0),
		.io_out_valid_0(_mesh_20_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10029 == GlobalFiModInstNr[0]) || (10029 == GlobalFiModInstNr[1]) || (10029 == GlobalFiModInstNr[2]) || (10029 == GlobalFiModInstNr[3]))));
	Tile mesh_20_19(
		.clock(clock),
		.io_in_a_0(r_659_0),
		.io_in_b_0(b_628_0),
		.io_in_d_0(b_1652_0),
		.io_in_control_0_dataflow(mesh_20_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2676_0),
		.io_in_last_0(r_3700_0),
		.io_in_valid_0(r_1652_0),
		.io_out_a_0(_mesh_20_19_io_out_a_0),
		.io_out_c_0(_mesh_20_19_io_out_c_0),
		.io_out_b_0(_mesh_20_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_19_io_out_id_0),
		.io_out_last_0(_mesh_20_19_io_out_last_0),
		.io_out_valid_0(_mesh_20_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10030 == GlobalFiModInstNr[0]) || (10030 == GlobalFiModInstNr[1]) || (10030 == GlobalFiModInstNr[2]) || (10030 == GlobalFiModInstNr[3]))));
	Tile mesh_20_20(
		.clock(clock),
		.io_in_a_0(r_660_0),
		.io_in_b_0(b_660_0),
		.io_in_d_0(b_1684_0),
		.io_in_control_0_dataflow(mesh_20_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2708_0),
		.io_in_last_0(r_3732_0),
		.io_in_valid_0(r_1684_0),
		.io_out_a_0(_mesh_20_20_io_out_a_0),
		.io_out_c_0(_mesh_20_20_io_out_c_0),
		.io_out_b_0(_mesh_20_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_20_io_out_id_0),
		.io_out_last_0(_mesh_20_20_io_out_last_0),
		.io_out_valid_0(_mesh_20_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10031 == GlobalFiModInstNr[0]) || (10031 == GlobalFiModInstNr[1]) || (10031 == GlobalFiModInstNr[2]) || (10031 == GlobalFiModInstNr[3]))));
	Tile mesh_20_21(
		.clock(clock),
		.io_in_a_0(r_661_0),
		.io_in_b_0(b_692_0),
		.io_in_d_0(b_1716_0),
		.io_in_control_0_dataflow(mesh_20_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2740_0),
		.io_in_last_0(r_3764_0),
		.io_in_valid_0(r_1716_0),
		.io_out_a_0(_mesh_20_21_io_out_a_0),
		.io_out_c_0(_mesh_20_21_io_out_c_0),
		.io_out_b_0(_mesh_20_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_21_io_out_id_0),
		.io_out_last_0(_mesh_20_21_io_out_last_0),
		.io_out_valid_0(_mesh_20_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10032 == GlobalFiModInstNr[0]) || (10032 == GlobalFiModInstNr[1]) || (10032 == GlobalFiModInstNr[2]) || (10032 == GlobalFiModInstNr[3]))));
	Tile mesh_20_22(
		.clock(clock),
		.io_in_a_0(r_662_0),
		.io_in_b_0(b_724_0),
		.io_in_d_0(b_1748_0),
		.io_in_control_0_dataflow(mesh_20_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2772_0),
		.io_in_last_0(r_3796_0),
		.io_in_valid_0(r_1748_0),
		.io_out_a_0(_mesh_20_22_io_out_a_0),
		.io_out_c_0(_mesh_20_22_io_out_c_0),
		.io_out_b_0(_mesh_20_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_22_io_out_id_0),
		.io_out_last_0(_mesh_20_22_io_out_last_0),
		.io_out_valid_0(_mesh_20_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10033 == GlobalFiModInstNr[0]) || (10033 == GlobalFiModInstNr[1]) || (10033 == GlobalFiModInstNr[2]) || (10033 == GlobalFiModInstNr[3]))));
	Tile mesh_20_23(
		.clock(clock),
		.io_in_a_0(r_663_0),
		.io_in_b_0(b_756_0),
		.io_in_d_0(b_1780_0),
		.io_in_control_0_dataflow(mesh_20_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2804_0),
		.io_in_last_0(r_3828_0),
		.io_in_valid_0(r_1780_0),
		.io_out_a_0(_mesh_20_23_io_out_a_0),
		.io_out_c_0(_mesh_20_23_io_out_c_0),
		.io_out_b_0(_mesh_20_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_23_io_out_id_0),
		.io_out_last_0(_mesh_20_23_io_out_last_0),
		.io_out_valid_0(_mesh_20_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10034 == GlobalFiModInstNr[0]) || (10034 == GlobalFiModInstNr[1]) || (10034 == GlobalFiModInstNr[2]) || (10034 == GlobalFiModInstNr[3]))));
	Tile mesh_20_24(
		.clock(clock),
		.io_in_a_0(r_664_0),
		.io_in_b_0(b_788_0),
		.io_in_d_0(b_1812_0),
		.io_in_control_0_dataflow(mesh_20_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2836_0),
		.io_in_last_0(r_3860_0),
		.io_in_valid_0(r_1812_0),
		.io_out_a_0(_mesh_20_24_io_out_a_0),
		.io_out_c_0(_mesh_20_24_io_out_c_0),
		.io_out_b_0(_mesh_20_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_24_io_out_id_0),
		.io_out_last_0(_mesh_20_24_io_out_last_0),
		.io_out_valid_0(_mesh_20_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10035 == GlobalFiModInstNr[0]) || (10035 == GlobalFiModInstNr[1]) || (10035 == GlobalFiModInstNr[2]) || (10035 == GlobalFiModInstNr[3]))));
	Tile mesh_20_25(
		.clock(clock),
		.io_in_a_0(r_665_0),
		.io_in_b_0(b_820_0),
		.io_in_d_0(b_1844_0),
		.io_in_control_0_dataflow(mesh_20_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2868_0),
		.io_in_last_0(r_3892_0),
		.io_in_valid_0(r_1844_0),
		.io_out_a_0(_mesh_20_25_io_out_a_0),
		.io_out_c_0(_mesh_20_25_io_out_c_0),
		.io_out_b_0(_mesh_20_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_25_io_out_id_0),
		.io_out_last_0(_mesh_20_25_io_out_last_0),
		.io_out_valid_0(_mesh_20_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10036 == GlobalFiModInstNr[0]) || (10036 == GlobalFiModInstNr[1]) || (10036 == GlobalFiModInstNr[2]) || (10036 == GlobalFiModInstNr[3]))));
	Tile mesh_20_26(
		.clock(clock),
		.io_in_a_0(r_666_0),
		.io_in_b_0(b_852_0),
		.io_in_d_0(b_1876_0),
		.io_in_control_0_dataflow(mesh_20_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2900_0),
		.io_in_last_0(r_3924_0),
		.io_in_valid_0(r_1876_0),
		.io_out_a_0(_mesh_20_26_io_out_a_0),
		.io_out_c_0(_mesh_20_26_io_out_c_0),
		.io_out_b_0(_mesh_20_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_26_io_out_id_0),
		.io_out_last_0(_mesh_20_26_io_out_last_0),
		.io_out_valid_0(_mesh_20_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10037 == GlobalFiModInstNr[0]) || (10037 == GlobalFiModInstNr[1]) || (10037 == GlobalFiModInstNr[2]) || (10037 == GlobalFiModInstNr[3]))));
	Tile mesh_20_27(
		.clock(clock),
		.io_in_a_0(r_667_0),
		.io_in_b_0(b_884_0),
		.io_in_d_0(b_1908_0),
		.io_in_control_0_dataflow(mesh_20_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2932_0),
		.io_in_last_0(r_3956_0),
		.io_in_valid_0(r_1908_0),
		.io_out_a_0(_mesh_20_27_io_out_a_0),
		.io_out_c_0(_mesh_20_27_io_out_c_0),
		.io_out_b_0(_mesh_20_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_27_io_out_id_0),
		.io_out_last_0(_mesh_20_27_io_out_last_0),
		.io_out_valid_0(_mesh_20_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10038 == GlobalFiModInstNr[0]) || (10038 == GlobalFiModInstNr[1]) || (10038 == GlobalFiModInstNr[2]) || (10038 == GlobalFiModInstNr[3]))));
	Tile mesh_20_28(
		.clock(clock),
		.io_in_a_0(r_668_0),
		.io_in_b_0(b_916_0),
		.io_in_d_0(b_1940_0),
		.io_in_control_0_dataflow(mesh_20_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2964_0),
		.io_in_last_0(r_3988_0),
		.io_in_valid_0(r_1940_0),
		.io_out_a_0(_mesh_20_28_io_out_a_0),
		.io_out_c_0(_mesh_20_28_io_out_c_0),
		.io_out_b_0(_mesh_20_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_28_io_out_id_0),
		.io_out_last_0(_mesh_20_28_io_out_last_0),
		.io_out_valid_0(_mesh_20_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10039 == GlobalFiModInstNr[0]) || (10039 == GlobalFiModInstNr[1]) || (10039 == GlobalFiModInstNr[2]) || (10039 == GlobalFiModInstNr[3]))));
	Tile mesh_20_29(
		.clock(clock),
		.io_in_a_0(r_669_0),
		.io_in_b_0(b_948_0),
		.io_in_d_0(b_1972_0),
		.io_in_control_0_dataflow(mesh_20_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2996_0),
		.io_in_last_0(r_4020_0),
		.io_in_valid_0(r_1972_0),
		.io_out_a_0(_mesh_20_29_io_out_a_0),
		.io_out_c_0(_mesh_20_29_io_out_c_0),
		.io_out_b_0(_mesh_20_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_29_io_out_id_0),
		.io_out_last_0(_mesh_20_29_io_out_last_0),
		.io_out_valid_0(_mesh_20_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10040 == GlobalFiModInstNr[0]) || (10040 == GlobalFiModInstNr[1]) || (10040 == GlobalFiModInstNr[2]) || (10040 == GlobalFiModInstNr[3]))));
	Tile mesh_20_30(
		.clock(clock),
		.io_in_a_0(r_670_0),
		.io_in_b_0(b_980_0),
		.io_in_d_0(b_2004_0),
		.io_in_control_0_dataflow(mesh_20_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3028_0),
		.io_in_last_0(r_4052_0),
		.io_in_valid_0(r_2004_0),
		.io_out_a_0(_mesh_20_30_io_out_a_0),
		.io_out_c_0(_mesh_20_30_io_out_c_0),
		.io_out_b_0(_mesh_20_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_30_io_out_id_0),
		.io_out_last_0(_mesh_20_30_io_out_last_0),
		.io_out_valid_0(_mesh_20_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10041 == GlobalFiModInstNr[0]) || (10041 == GlobalFiModInstNr[1]) || (10041 == GlobalFiModInstNr[2]) || (10041 == GlobalFiModInstNr[3]))));
	Tile mesh_20_31(
		.clock(clock),
		.io_in_a_0(r_671_0),
		.io_in_b_0(b_1012_0),
		.io_in_d_0(b_2036_0),
		.io_in_control_0_dataflow(mesh_20_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_20_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_20_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3060_0),
		.io_in_last_0(r_4084_0),
		.io_in_valid_0(r_2036_0),
		.io_out_a_0(_mesh_20_31_io_out_a_0),
		.io_out_c_0(_mesh_20_31_io_out_c_0),
		.io_out_b_0(_mesh_20_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_20_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_20_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_20_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_20_31_io_out_id_0),
		.io_out_last_0(_mesh_20_31_io_out_last_0),
		.io_out_valid_0(_mesh_20_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10042 == GlobalFiModInstNr[0]) || (10042 == GlobalFiModInstNr[1]) || (10042 == GlobalFiModInstNr[2]) || (10042 == GlobalFiModInstNr[3]))));
	Tile mesh_21_0(
		.clock(clock),
		.io_in_a_0(r_672_0),
		.io_in_b_0(b_21_0),
		.io_in_d_0(b_1045_0),
		.io_in_control_0_dataflow(mesh_21_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2069_0),
		.io_in_last_0(r_3093_0),
		.io_in_valid_0(r_1045_0),
		.io_out_a_0(_mesh_21_0_io_out_a_0),
		.io_out_c_0(_mesh_21_0_io_out_c_0),
		.io_out_b_0(_mesh_21_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_0_io_out_id_0),
		.io_out_last_0(_mesh_21_0_io_out_last_0),
		.io_out_valid_0(_mesh_21_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10043 == GlobalFiModInstNr[0]) || (10043 == GlobalFiModInstNr[1]) || (10043 == GlobalFiModInstNr[2]) || (10043 == GlobalFiModInstNr[3]))));
	Tile mesh_21_1(
		.clock(clock),
		.io_in_a_0(r_673_0),
		.io_in_b_0(b_53_0),
		.io_in_d_0(b_1077_0),
		.io_in_control_0_dataflow(mesh_21_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2101_0),
		.io_in_last_0(r_3125_0),
		.io_in_valid_0(r_1077_0),
		.io_out_a_0(_mesh_21_1_io_out_a_0),
		.io_out_c_0(_mesh_21_1_io_out_c_0),
		.io_out_b_0(_mesh_21_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_1_io_out_id_0),
		.io_out_last_0(_mesh_21_1_io_out_last_0),
		.io_out_valid_0(_mesh_21_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10044 == GlobalFiModInstNr[0]) || (10044 == GlobalFiModInstNr[1]) || (10044 == GlobalFiModInstNr[2]) || (10044 == GlobalFiModInstNr[3]))));
	Tile mesh_21_2(
		.clock(clock),
		.io_in_a_0(r_674_0),
		.io_in_b_0(b_85_0),
		.io_in_d_0(b_1109_0),
		.io_in_control_0_dataflow(mesh_21_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2133_0),
		.io_in_last_0(r_3157_0),
		.io_in_valid_0(r_1109_0),
		.io_out_a_0(_mesh_21_2_io_out_a_0),
		.io_out_c_0(_mesh_21_2_io_out_c_0),
		.io_out_b_0(_mesh_21_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_2_io_out_id_0),
		.io_out_last_0(_mesh_21_2_io_out_last_0),
		.io_out_valid_0(_mesh_21_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10045 == GlobalFiModInstNr[0]) || (10045 == GlobalFiModInstNr[1]) || (10045 == GlobalFiModInstNr[2]) || (10045 == GlobalFiModInstNr[3]))));
	Tile mesh_21_3(
		.clock(clock),
		.io_in_a_0(r_675_0),
		.io_in_b_0(b_117_0),
		.io_in_d_0(b_1141_0),
		.io_in_control_0_dataflow(mesh_21_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2165_0),
		.io_in_last_0(r_3189_0),
		.io_in_valid_0(r_1141_0),
		.io_out_a_0(_mesh_21_3_io_out_a_0),
		.io_out_c_0(_mesh_21_3_io_out_c_0),
		.io_out_b_0(_mesh_21_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_3_io_out_id_0),
		.io_out_last_0(_mesh_21_3_io_out_last_0),
		.io_out_valid_0(_mesh_21_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10046 == GlobalFiModInstNr[0]) || (10046 == GlobalFiModInstNr[1]) || (10046 == GlobalFiModInstNr[2]) || (10046 == GlobalFiModInstNr[3]))));
	Tile mesh_21_4(
		.clock(clock),
		.io_in_a_0(r_676_0),
		.io_in_b_0(b_149_0),
		.io_in_d_0(b_1173_0),
		.io_in_control_0_dataflow(mesh_21_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2197_0),
		.io_in_last_0(r_3221_0),
		.io_in_valid_0(r_1173_0),
		.io_out_a_0(_mesh_21_4_io_out_a_0),
		.io_out_c_0(_mesh_21_4_io_out_c_0),
		.io_out_b_0(_mesh_21_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_4_io_out_id_0),
		.io_out_last_0(_mesh_21_4_io_out_last_0),
		.io_out_valid_0(_mesh_21_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10047 == GlobalFiModInstNr[0]) || (10047 == GlobalFiModInstNr[1]) || (10047 == GlobalFiModInstNr[2]) || (10047 == GlobalFiModInstNr[3]))));
	Tile mesh_21_5(
		.clock(clock),
		.io_in_a_0(r_677_0),
		.io_in_b_0(b_181_0),
		.io_in_d_0(b_1205_0),
		.io_in_control_0_dataflow(mesh_21_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2229_0),
		.io_in_last_0(r_3253_0),
		.io_in_valid_0(r_1205_0),
		.io_out_a_0(_mesh_21_5_io_out_a_0),
		.io_out_c_0(_mesh_21_5_io_out_c_0),
		.io_out_b_0(_mesh_21_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_5_io_out_id_0),
		.io_out_last_0(_mesh_21_5_io_out_last_0),
		.io_out_valid_0(_mesh_21_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10048 == GlobalFiModInstNr[0]) || (10048 == GlobalFiModInstNr[1]) || (10048 == GlobalFiModInstNr[2]) || (10048 == GlobalFiModInstNr[3]))));
	Tile mesh_21_6(
		.clock(clock),
		.io_in_a_0(r_678_0),
		.io_in_b_0(b_213_0),
		.io_in_d_0(b_1237_0),
		.io_in_control_0_dataflow(mesh_21_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2261_0),
		.io_in_last_0(r_3285_0),
		.io_in_valid_0(r_1237_0),
		.io_out_a_0(_mesh_21_6_io_out_a_0),
		.io_out_c_0(_mesh_21_6_io_out_c_0),
		.io_out_b_0(_mesh_21_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_6_io_out_id_0),
		.io_out_last_0(_mesh_21_6_io_out_last_0),
		.io_out_valid_0(_mesh_21_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10049 == GlobalFiModInstNr[0]) || (10049 == GlobalFiModInstNr[1]) || (10049 == GlobalFiModInstNr[2]) || (10049 == GlobalFiModInstNr[3]))));
	Tile mesh_21_7(
		.clock(clock),
		.io_in_a_0(r_679_0),
		.io_in_b_0(b_245_0),
		.io_in_d_0(b_1269_0),
		.io_in_control_0_dataflow(mesh_21_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2293_0),
		.io_in_last_0(r_3317_0),
		.io_in_valid_0(r_1269_0),
		.io_out_a_0(_mesh_21_7_io_out_a_0),
		.io_out_c_0(_mesh_21_7_io_out_c_0),
		.io_out_b_0(_mesh_21_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_7_io_out_id_0),
		.io_out_last_0(_mesh_21_7_io_out_last_0),
		.io_out_valid_0(_mesh_21_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10050 == GlobalFiModInstNr[0]) || (10050 == GlobalFiModInstNr[1]) || (10050 == GlobalFiModInstNr[2]) || (10050 == GlobalFiModInstNr[3]))));
	Tile mesh_21_8(
		.clock(clock),
		.io_in_a_0(r_680_0),
		.io_in_b_0(b_277_0),
		.io_in_d_0(b_1301_0),
		.io_in_control_0_dataflow(mesh_21_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2325_0),
		.io_in_last_0(r_3349_0),
		.io_in_valid_0(r_1301_0),
		.io_out_a_0(_mesh_21_8_io_out_a_0),
		.io_out_c_0(_mesh_21_8_io_out_c_0),
		.io_out_b_0(_mesh_21_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_8_io_out_id_0),
		.io_out_last_0(_mesh_21_8_io_out_last_0),
		.io_out_valid_0(_mesh_21_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10051 == GlobalFiModInstNr[0]) || (10051 == GlobalFiModInstNr[1]) || (10051 == GlobalFiModInstNr[2]) || (10051 == GlobalFiModInstNr[3]))));
	Tile mesh_21_9(
		.clock(clock),
		.io_in_a_0(r_681_0),
		.io_in_b_0(b_309_0),
		.io_in_d_0(b_1333_0),
		.io_in_control_0_dataflow(mesh_21_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2357_0),
		.io_in_last_0(r_3381_0),
		.io_in_valid_0(r_1333_0),
		.io_out_a_0(_mesh_21_9_io_out_a_0),
		.io_out_c_0(_mesh_21_9_io_out_c_0),
		.io_out_b_0(_mesh_21_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_9_io_out_id_0),
		.io_out_last_0(_mesh_21_9_io_out_last_0),
		.io_out_valid_0(_mesh_21_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10052 == GlobalFiModInstNr[0]) || (10052 == GlobalFiModInstNr[1]) || (10052 == GlobalFiModInstNr[2]) || (10052 == GlobalFiModInstNr[3]))));
	Tile mesh_21_10(
		.clock(clock),
		.io_in_a_0(r_682_0),
		.io_in_b_0(b_341_0),
		.io_in_d_0(b_1365_0),
		.io_in_control_0_dataflow(mesh_21_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2389_0),
		.io_in_last_0(r_3413_0),
		.io_in_valid_0(r_1365_0),
		.io_out_a_0(_mesh_21_10_io_out_a_0),
		.io_out_c_0(_mesh_21_10_io_out_c_0),
		.io_out_b_0(_mesh_21_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_10_io_out_id_0),
		.io_out_last_0(_mesh_21_10_io_out_last_0),
		.io_out_valid_0(_mesh_21_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10053 == GlobalFiModInstNr[0]) || (10053 == GlobalFiModInstNr[1]) || (10053 == GlobalFiModInstNr[2]) || (10053 == GlobalFiModInstNr[3]))));
	Tile mesh_21_11(
		.clock(clock),
		.io_in_a_0(r_683_0),
		.io_in_b_0(b_373_0),
		.io_in_d_0(b_1397_0),
		.io_in_control_0_dataflow(mesh_21_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2421_0),
		.io_in_last_0(r_3445_0),
		.io_in_valid_0(r_1397_0),
		.io_out_a_0(_mesh_21_11_io_out_a_0),
		.io_out_c_0(_mesh_21_11_io_out_c_0),
		.io_out_b_0(_mesh_21_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_11_io_out_id_0),
		.io_out_last_0(_mesh_21_11_io_out_last_0),
		.io_out_valid_0(_mesh_21_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10054 == GlobalFiModInstNr[0]) || (10054 == GlobalFiModInstNr[1]) || (10054 == GlobalFiModInstNr[2]) || (10054 == GlobalFiModInstNr[3]))));
	Tile mesh_21_12(
		.clock(clock),
		.io_in_a_0(r_684_0),
		.io_in_b_0(b_405_0),
		.io_in_d_0(b_1429_0),
		.io_in_control_0_dataflow(mesh_21_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2453_0),
		.io_in_last_0(r_3477_0),
		.io_in_valid_0(r_1429_0),
		.io_out_a_0(_mesh_21_12_io_out_a_0),
		.io_out_c_0(_mesh_21_12_io_out_c_0),
		.io_out_b_0(_mesh_21_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_12_io_out_id_0),
		.io_out_last_0(_mesh_21_12_io_out_last_0),
		.io_out_valid_0(_mesh_21_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10055 == GlobalFiModInstNr[0]) || (10055 == GlobalFiModInstNr[1]) || (10055 == GlobalFiModInstNr[2]) || (10055 == GlobalFiModInstNr[3]))));
	Tile mesh_21_13(
		.clock(clock),
		.io_in_a_0(r_685_0),
		.io_in_b_0(b_437_0),
		.io_in_d_0(b_1461_0),
		.io_in_control_0_dataflow(mesh_21_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2485_0),
		.io_in_last_0(r_3509_0),
		.io_in_valid_0(r_1461_0),
		.io_out_a_0(_mesh_21_13_io_out_a_0),
		.io_out_c_0(_mesh_21_13_io_out_c_0),
		.io_out_b_0(_mesh_21_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_13_io_out_id_0),
		.io_out_last_0(_mesh_21_13_io_out_last_0),
		.io_out_valid_0(_mesh_21_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10056 == GlobalFiModInstNr[0]) || (10056 == GlobalFiModInstNr[1]) || (10056 == GlobalFiModInstNr[2]) || (10056 == GlobalFiModInstNr[3]))));
	Tile mesh_21_14(
		.clock(clock),
		.io_in_a_0(r_686_0),
		.io_in_b_0(b_469_0),
		.io_in_d_0(b_1493_0),
		.io_in_control_0_dataflow(mesh_21_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2517_0),
		.io_in_last_0(r_3541_0),
		.io_in_valid_0(r_1493_0),
		.io_out_a_0(_mesh_21_14_io_out_a_0),
		.io_out_c_0(_mesh_21_14_io_out_c_0),
		.io_out_b_0(_mesh_21_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_14_io_out_id_0),
		.io_out_last_0(_mesh_21_14_io_out_last_0),
		.io_out_valid_0(_mesh_21_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10057 == GlobalFiModInstNr[0]) || (10057 == GlobalFiModInstNr[1]) || (10057 == GlobalFiModInstNr[2]) || (10057 == GlobalFiModInstNr[3]))));
	Tile mesh_21_15(
		.clock(clock),
		.io_in_a_0(r_687_0),
		.io_in_b_0(b_501_0),
		.io_in_d_0(b_1525_0),
		.io_in_control_0_dataflow(mesh_21_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2549_0),
		.io_in_last_0(r_3573_0),
		.io_in_valid_0(r_1525_0),
		.io_out_a_0(_mesh_21_15_io_out_a_0),
		.io_out_c_0(_mesh_21_15_io_out_c_0),
		.io_out_b_0(_mesh_21_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_15_io_out_id_0),
		.io_out_last_0(_mesh_21_15_io_out_last_0),
		.io_out_valid_0(_mesh_21_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10058 == GlobalFiModInstNr[0]) || (10058 == GlobalFiModInstNr[1]) || (10058 == GlobalFiModInstNr[2]) || (10058 == GlobalFiModInstNr[3]))));
	Tile mesh_21_16(
		.clock(clock),
		.io_in_a_0(r_688_0),
		.io_in_b_0(b_533_0),
		.io_in_d_0(b_1557_0),
		.io_in_control_0_dataflow(mesh_21_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2581_0),
		.io_in_last_0(r_3605_0),
		.io_in_valid_0(r_1557_0),
		.io_out_a_0(_mesh_21_16_io_out_a_0),
		.io_out_c_0(_mesh_21_16_io_out_c_0),
		.io_out_b_0(_mesh_21_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_16_io_out_id_0),
		.io_out_last_0(_mesh_21_16_io_out_last_0),
		.io_out_valid_0(_mesh_21_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10059 == GlobalFiModInstNr[0]) || (10059 == GlobalFiModInstNr[1]) || (10059 == GlobalFiModInstNr[2]) || (10059 == GlobalFiModInstNr[3]))));
	Tile mesh_21_17(
		.clock(clock),
		.io_in_a_0(r_689_0),
		.io_in_b_0(b_565_0),
		.io_in_d_0(b_1589_0),
		.io_in_control_0_dataflow(mesh_21_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2613_0),
		.io_in_last_0(r_3637_0),
		.io_in_valid_0(r_1589_0),
		.io_out_a_0(_mesh_21_17_io_out_a_0),
		.io_out_c_0(_mesh_21_17_io_out_c_0),
		.io_out_b_0(_mesh_21_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_17_io_out_id_0),
		.io_out_last_0(_mesh_21_17_io_out_last_0),
		.io_out_valid_0(_mesh_21_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10060 == GlobalFiModInstNr[0]) || (10060 == GlobalFiModInstNr[1]) || (10060 == GlobalFiModInstNr[2]) || (10060 == GlobalFiModInstNr[3]))));
	Tile mesh_21_18(
		.clock(clock),
		.io_in_a_0(r_690_0),
		.io_in_b_0(b_597_0),
		.io_in_d_0(b_1621_0),
		.io_in_control_0_dataflow(mesh_21_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2645_0),
		.io_in_last_0(r_3669_0),
		.io_in_valid_0(r_1621_0),
		.io_out_a_0(_mesh_21_18_io_out_a_0),
		.io_out_c_0(_mesh_21_18_io_out_c_0),
		.io_out_b_0(_mesh_21_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_18_io_out_id_0),
		.io_out_last_0(_mesh_21_18_io_out_last_0),
		.io_out_valid_0(_mesh_21_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10061 == GlobalFiModInstNr[0]) || (10061 == GlobalFiModInstNr[1]) || (10061 == GlobalFiModInstNr[2]) || (10061 == GlobalFiModInstNr[3]))));
	Tile mesh_21_19(
		.clock(clock),
		.io_in_a_0(r_691_0),
		.io_in_b_0(b_629_0),
		.io_in_d_0(b_1653_0),
		.io_in_control_0_dataflow(mesh_21_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2677_0),
		.io_in_last_0(r_3701_0),
		.io_in_valid_0(r_1653_0),
		.io_out_a_0(_mesh_21_19_io_out_a_0),
		.io_out_c_0(_mesh_21_19_io_out_c_0),
		.io_out_b_0(_mesh_21_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_19_io_out_id_0),
		.io_out_last_0(_mesh_21_19_io_out_last_0),
		.io_out_valid_0(_mesh_21_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10062 == GlobalFiModInstNr[0]) || (10062 == GlobalFiModInstNr[1]) || (10062 == GlobalFiModInstNr[2]) || (10062 == GlobalFiModInstNr[3]))));
	Tile mesh_21_20(
		.clock(clock),
		.io_in_a_0(r_692_0),
		.io_in_b_0(b_661_0),
		.io_in_d_0(b_1685_0),
		.io_in_control_0_dataflow(mesh_21_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2709_0),
		.io_in_last_0(r_3733_0),
		.io_in_valid_0(r_1685_0),
		.io_out_a_0(_mesh_21_20_io_out_a_0),
		.io_out_c_0(_mesh_21_20_io_out_c_0),
		.io_out_b_0(_mesh_21_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_20_io_out_id_0),
		.io_out_last_0(_mesh_21_20_io_out_last_0),
		.io_out_valid_0(_mesh_21_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10063 == GlobalFiModInstNr[0]) || (10063 == GlobalFiModInstNr[1]) || (10063 == GlobalFiModInstNr[2]) || (10063 == GlobalFiModInstNr[3]))));
	Tile mesh_21_21(
		.clock(clock),
		.io_in_a_0(r_693_0),
		.io_in_b_0(b_693_0),
		.io_in_d_0(b_1717_0),
		.io_in_control_0_dataflow(mesh_21_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2741_0),
		.io_in_last_0(r_3765_0),
		.io_in_valid_0(r_1717_0),
		.io_out_a_0(_mesh_21_21_io_out_a_0),
		.io_out_c_0(_mesh_21_21_io_out_c_0),
		.io_out_b_0(_mesh_21_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_21_io_out_id_0),
		.io_out_last_0(_mesh_21_21_io_out_last_0),
		.io_out_valid_0(_mesh_21_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10064 == GlobalFiModInstNr[0]) || (10064 == GlobalFiModInstNr[1]) || (10064 == GlobalFiModInstNr[2]) || (10064 == GlobalFiModInstNr[3]))));
	Tile mesh_21_22(
		.clock(clock),
		.io_in_a_0(r_694_0),
		.io_in_b_0(b_725_0),
		.io_in_d_0(b_1749_0),
		.io_in_control_0_dataflow(mesh_21_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2773_0),
		.io_in_last_0(r_3797_0),
		.io_in_valid_0(r_1749_0),
		.io_out_a_0(_mesh_21_22_io_out_a_0),
		.io_out_c_0(_mesh_21_22_io_out_c_0),
		.io_out_b_0(_mesh_21_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_22_io_out_id_0),
		.io_out_last_0(_mesh_21_22_io_out_last_0),
		.io_out_valid_0(_mesh_21_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10065 == GlobalFiModInstNr[0]) || (10065 == GlobalFiModInstNr[1]) || (10065 == GlobalFiModInstNr[2]) || (10065 == GlobalFiModInstNr[3]))));
	Tile mesh_21_23(
		.clock(clock),
		.io_in_a_0(r_695_0),
		.io_in_b_0(b_757_0),
		.io_in_d_0(b_1781_0),
		.io_in_control_0_dataflow(mesh_21_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2805_0),
		.io_in_last_0(r_3829_0),
		.io_in_valid_0(r_1781_0),
		.io_out_a_0(_mesh_21_23_io_out_a_0),
		.io_out_c_0(_mesh_21_23_io_out_c_0),
		.io_out_b_0(_mesh_21_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_23_io_out_id_0),
		.io_out_last_0(_mesh_21_23_io_out_last_0),
		.io_out_valid_0(_mesh_21_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10066 == GlobalFiModInstNr[0]) || (10066 == GlobalFiModInstNr[1]) || (10066 == GlobalFiModInstNr[2]) || (10066 == GlobalFiModInstNr[3]))));
	Tile mesh_21_24(
		.clock(clock),
		.io_in_a_0(r_696_0),
		.io_in_b_0(b_789_0),
		.io_in_d_0(b_1813_0),
		.io_in_control_0_dataflow(mesh_21_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2837_0),
		.io_in_last_0(r_3861_0),
		.io_in_valid_0(r_1813_0),
		.io_out_a_0(_mesh_21_24_io_out_a_0),
		.io_out_c_0(_mesh_21_24_io_out_c_0),
		.io_out_b_0(_mesh_21_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_24_io_out_id_0),
		.io_out_last_0(_mesh_21_24_io_out_last_0),
		.io_out_valid_0(_mesh_21_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10067 == GlobalFiModInstNr[0]) || (10067 == GlobalFiModInstNr[1]) || (10067 == GlobalFiModInstNr[2]) || (10067 == GlobalFiModInstNr[3]))));
	Tile mesh_21_25(
		.clock(clock),
		.io_in_a_0(r_697_0),
		.io_in_b_0(b_821_0),
		.io_in_d_0(b_1845_0),
		.io_in_control_0_dataflow(mesh_21_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2869_0),
		.io_in_last_0(r_3893_0),
		.io_in_valid_0(r_1845_0),
		.io_out_a_0(_mesh_21_25_io_out_a_0),
		.io_out_c_0(_mesh_21_25_io_out_c_0),
		.io_out_b_0(_mesh_21_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_25_io_out_id_0),
		.io_out_last_0(_mesh_21_25_io_out_last_0),
		.io_out_valid_0(_mesh_21_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10068 == GlobalFiModInstNr[0]) || (10068 == GlobalFiModInstNr[1]) || (10068 == GlobalFiModInstNr[2]) || (10068 == GlobalFiModInstNr[3]))));
	Tile mesh_21_26(
		.clock(clock),
		.io_in_a_0(r_698_0),
		.io_in_b_0(b_853_0),
		.io_in_d_0(b_1877_0),
		.io_in_control_0_dataflow(mesh_21_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2901_0),
		.io_in_last_0(r_3925_0),
		.io_in_valid_0(r_1877_0),
		.io_out_a_0(_mesh_21_26_io_out_a_0),
		.io_out_c_0(_mesh_21_26_io_out_c_0),
		.io_out_b_0(_mesh_21_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_26_io_out_id_0),
		.io_out_last_0(_mesh_21_26_io_out_last_0),
		.io_out_valid_0(_mesh_21_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10069 == GlobalFiModInstNr[0]) || (10069 == GlobalFiModInstNr[1]) || (10069 == GlobalFiModInstNr[2]) || (10069 == GlobalFiModInstNr[3]))));
	Tile mesh_21_27(
		.clock(clock),
		.io_in_a_0(r_699_0),
		.io_in_b_0(b_885_0),
		.io_in_d_0(b_1909_0),
		.io_in_control_0_dataflow(mesh_21_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2933_0),
		.io_in_last_0(r_3957_0),
		.io_in_valid_0(r_1909_0),
		.io_out_a_0(_mesh_21_27_io_out_a_0),
		.io_out_c_0(_mesh_21_27_io_out_c_0),
		.io_out_b_0(_mesh_21_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_27_io_out_id_0),
		.io_out_last_0(_mesh_21_27_io_out_last_0),
		.io_out_valid_0(_mesh_21_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10070 == GlobalFiModInstNr[0]) || (10070 == GlobalFiModInstNr[1]) || (10070 == GlobalFiModInstNr[2]) || (10070 == GlobalFiModInstNr[3]))));
	Tile mesh_21_28(
		.clock(clock),
		.io_in_a_0(r_700_0),
		.io_in_b_0(b_917_0),
		.io_in_d_0(b_1941_0),
		.io_in_control_0_dataflow(mesh_21_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2965_0),
		.io_in_last_0(r_3989_0),
		.io_in_valid_0(r_1941_0),
		.io_out_a_0(_mesh_21_28_io_out_a_0),
		.io_out_c_0(_mesh_21_28_io_out_c_0),
		.io_out_b_0(_mesh_21_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_28_io_out_id_0),
		.io_out_last_0(_mesh_21_28_io_out_last_0),
		.io_out_valid_0(_mesh_21_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10071 == GlobalFiModInstNr[0]) || (10071 == GlobalFiModInstNr[1]) || (10071 == GlobalFiModInstNr[2]) || (10071 == GlobalFiModInstNr[3]))));
	Tile mesh_21_29(
		.clock(clock),
		.io_in_a_0(r_701_0),
		.io_in_b_0(b_949_0),
		.io_in_d_0(b_1973_0),
		.io_in_control_0_dataflow(mesh_21_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2997_0),
		.io_in_last_0(r_4021_0),
		.io_in_valid_0(r_1973_0),
		.io_out_a_0(_mesh_21_29_io_out_a_0),
		.io_out_c_0(_mesh_21_29_io_out_c_0),
		.io_out_b_0(_mesh_21_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_29_io_out_id_0),
		.io_out_last_0(_mesh_21_29_io_out_last_0),
		.io_out_valid_0(_mesh_21_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10072 == GlobalFiModInstNr[0]) || (10072 == GlobalFiModInstNr[1]) || (10072 == GlobalFiModInstNr[2]) || (10072 == GlobalFiModInstNr[3]))));
	Tile mesh_21_30(
		.clock(clock),
		.io_in_a_0(r_702_0),
		.io_in_b_0(b_981_0),
		.io_in_d_0(b_2005_0),
		.io_in_control_0_dataflow(mesh_21_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3029_0),
		.io_in_last_0(r_4053_0),
		.io_in_valid_0(r_2005_0),
		.io_out_a_0(_mesh_21_30_io_out_a_0),
		.io_out_c_0(_mesh_21_30_io_out_c_0),
		.io_out_b_0(_mesh_21_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_30_io_out_id_0),
		.io_out_last_0(_mesh_21_30_io_out_last_0),
		.io_out_valid_0(_mesh_21_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10073 == GlobalFiModInstNr[0]) || (10073 == GlobalFiModInstNr[1]) || (10073 == GlobalFiModInstNr[2]) || (10073 == GlobalFiModInstNr[3]))));
	Tile mesh_21_31(
		.clock(clock),
		.io_in_a_0(r_703_0),
		.io_in_b_0(b_1013_0),
		.io_in_d_0(b_2037_0),
		.io_in_control_0_dataflow(mesh_21_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_21_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_21_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3061_0),
		.io_in_last_0(r_4085_0),
		.io_in_valid_0(r_2037_0),
		.io_out_a_0(_mesh_21_31_io_out_a_0),
		.io_out_c_0(_mesh_21_31_io_out_c_0),
		.io_out_b_0(_mesh_21_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_21_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_21_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_21_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_21_31_io_out_id_0),
		.io_out_last_0(_mesh_21_31_io_out_last_0),
		.io_out_valid_0(_mesh_21_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10074 == GlobalFiModInstNr[0]) || (10074 == GlobalFiModInstNr[1]) || (10074 == GlobalFiModInstNr[2]) || (10074 == GlobalFiModInstNr[3]))));
	Tile mesh_22_0(
		.clock(clock),
		.io_in_a_0(r_704_0),
		.io_in_b_0(b_22_0),
		.io_in_d_0(b_1046_0),
		.io_in_control_0_dataflow(mesh_22_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2070_0),
		.io_in_last_0(r_3094_0),
		.io_in_valid_0(r_1046_0),
		.io_out_a_0(_mesh_22_0_io_out_a_0),
		.io_out_c_0(_mesh_22_0_io_out_c_0),
		.io_out_b_0(_mesh_22_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_0_io_out_id_0),
		.io_out_last_0(_mesh_22_0_io_out_last_0),
		.io_out_valid_0(_mesh_22_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10075 == GlobalFiModInstNr[0]) || (10075 == GlobalFiModInstNr[1]) || (10075 == GlobalFiModInstNr[2]) || (10075 == GlobalFiModInstNr[3]))));
	Tile mesh_22_1(
		.clock(clock),
		.io_in_a_0(r_705_0),
		.io_in_b_0(b_54_0),
		.io_in_d_0(b_1078_0),
		.io_in_control_0_dataflow(mesh_22_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2102_0),
		.io_in_last_0(r_3126_0),
		.io_in_valid_0(r_1078_0),
		.io_out_a_0(_mesh_22_1_io_out_a_0),
		.io_out_c_0(_mesh_22_1_io_out_c_0),
		.io_out_b_0(_mesh_22_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_1_io_out_id_0),
		.io_out_last_0(_mesh_22_1_io_out_last_0),
		.io_out_valid_0(_mesh_22_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10076 == GlobalFiModInstNr[0]) || (10076 == GlobalFiModInstNr[1]) || (10076 == GlobalFiModInstNr[2]) || (10076 == GlobalFiModInstNr[3]))));
	Tile mesh_22_2(
		.clock(clock),
		.io_in_a_0(r_706_0),
		.io_in_b_0(b_86_0),
		.io_in_d_0(b_1110_0),
		.io_in_control_0_dataflow(mesh_22_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2134_0),
		.io_in_last_0(r_3158_0),
		.io_in_valid_0(r_1110_0),
		.io_out_a_0(_mesh_22_2_io_out_a_0),
		.io_out_c_0(_mesh_22_2_io_out_c_0),
		.io_out_b_0(_mesh_22_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_2_io_out_id_0),
		.io_out_last_0(_mesh_22_2_io_out_last_0),
		.io_out_valid_0(_mesh_22_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10077 == GlobalFiModInstNr[0]) || (10077 == GlobalFiModInstNr[1]) || (10077 == GlobalFiModInstNr[2]) || (10077 == GlobalFiModInstNr[3]))));
	Tile mesh_22_3(
		.clock(clock),
		.io_in_a_0(r_707_0),
		.io_in_b_0(b_118_0),
		.io_in_d_0(b_1142_0),
		.io_in_control_0_dataflow(mesh_22_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2166_0),
		.io_in_last_0(r_3190_0),
		.io_in_valid_0(r_1142_0),
		.io_out_a_0(_mesh_22_3_io_out_a_0),
		.io_out_c_0(_mesh_22_3_io_out_c_0),
		.io_out_b_0(_mesh_22_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_3_io_out_id_0),
		.io_out_last_0(_mesh_22_3_io_out_last_0),
		.io_out_valid_0(_mesh_22_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10078 == GlobalFiModInstNr[0]) || (10078 == GlobalFiModInstNr[1]) || (10078 == GlobalFiModInstNr[2]) || (10078 == GlobalFiModInstNr[3]))));
	Tile mesh_22_4(
		.clock(clock),
		.io_in_a_0(r_708_0),
		.io_in_b_0(b_150_0),
		.io_in_d_0(b_1174_0),
		.io_in_control_0_dataflow(mesh_22_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2198_0),
		.io_in_last_0(r_3222_0),
		.io_in_valid_0(r_1174_0),
		.io_out_a_0(_mesh_22_4_io_out_a_0),
		.io_out_c_0(_mesh_22_4_io_out_c_0),
		.io_out_b_0(_mesh_22_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_4_io_out_id_0),
		.io_out_last_0(_mesh_22_4_io_out_last_0),
		.io_out_valid_0(_mesh_22_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10079 == GlobalFiModInstNr[0]) || (10079 == GlobalFiModInstNr[1]) || (10079 == GlobalFiModInstNr[2]) || (10079 == GlobalFiModInstNr[3]))));
	Tile mesh_22_5(
		.clock(clock),
		.io_in_a_0(r_709_0),
		.io_in_b_0(b_182_0),
		.io_in_d_0(b_1206_0),
		.io_in_control_0_dataflow(mesh_22_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2230_0),
		.io_in_last_0(r_3254_0),
		.io_in_valid_0(r_1206_0),
		.io_out_a_0(_mesh_22_5_io_out_a_0),
		.io_out_c_0(_mesh_22_5_io_out_c_0),
		.io_out_b_0(_mesh_22_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_5_io_out_id_0),
		.io_out_last_0(_mesh_22_5_io_out_last_0),
		.io_out_valid_0(_mesh_22_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10080 == GlobalFiModInstNr[0]) || (10080 == GlobalFiModInstNr[1]) || (10080 == GlobalFiModInstNr[2]) || (10080 == GlobalFiModInstNr[3]))));
	Tile mesh_22_6(
		.clock(clock),
		.io_in_a_0(r_710_0),
		.io_in_b_0(b_214_0),
		.io_in_d_0(b_1238_0),
		.io_in_control_0_dataflow(mesh_22_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2262_0),
		.io_in_last_0(r_3286_0),
		.io_in_valid_0(r_1238_0),
		.io_out_a_0(_mesh_22_6_io_out_a_0),
		.io_out_c_0(_mesh_22_6_io_out_c_0),
		.io_out_b_0(_mesh_22_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_6_io_out_id_0),
		.io_out_last_0(_mesh_22_6_io_out_last_0),
		.io_out_valid_0(_mesh_22_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10081 == GlobalFiModInstNr[0]) || (10081 == GlobalFiModInstNr[1]) || (10081 == GlobalFiModInstNr[2]) || (10081 == GlobalFiModInstNr[3]))));
	Tile mesh_22_7(
		.clock(clock),
		.io_in_a_0(r_711_0),
		.io_in_b_0(b_246_0),
		.io_in_d_0(b_1270_0),
		.io_in_control_0_dataflow(mesh_22_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2294_0),
		.io_in_last_0(r_3318_0),
		.io_in_valid_0(r_1270_0),
		.io_out_a_0(_mesh_22_7_io_out_a_0),
		.io_out_c_0(_mesh_22_7_io_out_c_0),
		.io_out_b_0(_mesh_22_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_7_io_out_id_0),
		.io_out_last_0(_mesh_22_7_io_out_last_0),
		.io_out_valid_0(_mesh_22_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10082 == GlobalFiModInstNr[0]) || (10082 == GlobalFiModInstNr[1]) || (10082 == GlobalFiModInstNr[2]) || (10082 == GlobalFiModInstNr[3]))));
	Tile mesh_22_8(
		.clock(clock),
		.io_in_a_0(r_712_0),
		.io_in_b_0(b_278_0),
		.io_in_d_0(b_1302_0),
		.io_in_control_0_dataflow(mesh_22_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2326_0),
		.io_in_last_0(r_3350_0),
		.io_in_valid_0(r_1302_0),
		.io_out_a_0(_mesh_22_8_io_out_a_0),
		.io_out_c_0(_mesh_22_8_io_out_c_0),
		.io_out_b_0(_mesh_22_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_8_io_out_id_0),
		.io_out_last_0(_mesh_22_8_io_out_last_0),
		.io_out_valid_0(_mesh_22_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10083 == GlobalFiModInstNr[0]) || (10083 == GlobalFiModInstNr[1]) || (10083 == GlobalFiModInstNr[2]) || (10083 == GlobalFiModInstNr[3]))));
	Tile mesh_22_9(
		.clock(clock),
		.io_in_a_0(r_713_0),
		.io_in_b_0(b_310_0),
		.io_in_d_0(b_1334_0),
		.io_in_control_0_dataflow(mesh_22_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2358_0),
		.io_in_last_0(r_3382_0),
		.io_in_valid_0(r_1334_0),
		.io_out_a_0(_mesh_22_9_io_out_a_0),
		.io_out_c_0(_mesh_22_9_io_out_c_0),
		.io_out_b_0(_mesh_22_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_9_io_out_id_0),
		.io_out_last_0(_mesh_22_9_io_out_last_0),
		.io_out_valid_0(_mesh_22_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10084 == GlobalFiModInstNr[0]) || (10084 == GlobalFiModInstNr[1]) || (10084 == GlobalFiModInstNr[2]) || (10084 == GlobalFiModInstNr[3]))));
	Tile mesh_22_10(
		.clock(clock),
		.io_in_a_0(r_714_0),
		.io_in_b_0(b_342_0),
		.io_in_d_0(b_1366_0),
		.io_in_control_0_dataflow(mesh_22_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2390_0),
		.io_in_last_0(r_3414_0),
		.io_in_valid_0(r_1366_0),
		.io_out_a_0(_mesh_22_10_io_out_a_0),
		.io_out_c_0(_mesh_22_10_io_out_c_0),
		.io_out_b_0(_mesh_22_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_10_io_out_id_0),
		.io_out_last_0(_mesh_22_10_io_out_last_0),
		.io_out_valid_0(_mesh_22_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10085 == GlobalFiModInstNr[0]) || (10085 == GlobalFiModInstNr[1]) || (10085 == GlobalFiModInstNr[2]) || (10085 == GlobalFiModInstNr[3]))));
	Tile mesh_22_11(
		.clock(clock),
		.io_in_a_0(r_715_0),
		.io_in_b_0(b_374_0),
		.io_in_d_0(b_1398_0),
		.io_in_control_0_dataflow(mesh_22_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2422_0),
		.io_in_last_0(r_3446_0),
		.io_in_valid_0(r_1398_0),
		.io_out_a_0(_mesh_22_11_io_out_a_0),
		.io_out_c_0(_mesh_22_11_io_out_c_0),
		.io_out_b_0(_mesh_22_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_11_io_out_id_0),
		.io_out_last_0(_mesh_22_11_io_out_last_0),
		.io_out_valid_0(_mesh_22_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10086 == GlobalFiModInstNr[0]) || (10086 == GlobalFiModInstNr[1]) || (10086 == GlobalFiModInstNr[2]) || (10086 == GlobalFiModInstNr[3]))));
	Tile mesh_22_12(
		.clock(clock),
		.io_in_a_0(r_716_0),
		.io_in_b_0(b_406_0),
		.io_in_d_0(b_1430_0),
		.io_in_control_0_dataflow(mesh_22_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2454_0),
		.io_in_last_0(r_3478_0),
		.io_in_valid_0(r_1430_0),
		.io_out_a_0(_mesh_22_12_io_out_a_0),
		.io_out_c_0(_mesh_22_12_io_out_c_0),
		.io_out_b_0(_mesh_22_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_12_io_out_id_0),
		.io_out_last_0(_mesh_22_12_io_out_last_0),
		.io_out_valid_0(_mesh_22_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10087 == GlobalFiModInstNr[0]) || (10087 == GlobalFiModInstNr[1]) || (10087 == GlobalFiModInstNr[2]) || (10087 == GlobalFiModInstNr[3]))));
	Tile mesh_22_13(
		.clock(clock),
		.io_in_a_0(r_717_0),
		.io_in_b_0(b_438_0),
		.io_in_d_0(b_1462_0),
		.io_in_control_0_dataflow(mesh_22_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2486_0),
		.io_in_last_0(r_3510_0),
		.io_in_valid_0(r_1462_0),
		.io_out_a_0(_mesh_22_13_io_out_a_0),
		.io_out_c_0(_mesh_22_13_io_out_c_0),
		.io_out_b_0(_mesh_22_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_13_io_out_id_0),
		.io_out_last_0(_mesh_22_13_io_out_last_0),
		.io_out_valid_0(_mesh_22_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10088 == GlobalFiModInstNr[0]) || (10088 == GlobalFiModInstNr[1]) || (10088 == GlobalFiModInstNr[2]) || (10088 == GlobalFiModInstNr[3]))));
	Tile mesh_22_14(
		.clock(clock),
		.io_in_a_0(r_718_0),
		.io_in_b_0(b_470_0),
		.io_in_d_0(b_1494_0),
		.io_in_control_0_dataflow(mesh_22_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2518_0),
		.io_in_last_0(r_3542_0),
		.io_in_valid_0(r_1494_0),
		.io_out_a_0(_mesh_22_14_io_out_a_0),
		.io_out_c_0(_mesh_22_14_io_out_c_0),
		.io_out_b_0(_mesh_22_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_14_io_out_id_0),
		.io_out_last_0(_mesh_22_14_io_out_last_0),
		.io_out_valid_0(_mesh_22_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10089 == GlobalFiModInstNr[0]) || (10089 == GlobalFiModInstNr[1]) || (10089 == GlobalFiModInstNr[2]) || (10089 == GlobalFiModInstNr[3]))));
	Tile mesh_22_15(
		.clock(clock),
		.io_in_a_0(r_719_0),
		.io_in_b_0(b_502_0),
		.io_in_d_0(b_1526_0),
		.io_in_control_0_dataflow(mesh_22_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2550_0),
		.io_in_last_0(r_3574_0),
		.io_in_valid_0(r_1526_0),
		.io_out_a_0(_mesh_22_15_io_out_a_0),
		.io_out_c_0(_mesh_22_15_io_out_c_0),
		.io_out_b_0(_mesh_22_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_15_io_out_id_0),
		.io_out_last_0(_mesh_22_15_io_out_last_0),
		.io_out_valid_0(_mesh_22_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10090 == GlobalFiModInstNr[0]) || (10090 == GlobalFiModInstNr[1]) || (10090 == GlobalFiModInstNr[2]) || (10090 == GlobalFiModInstNr[3]))));
	Tile mesh_22_16(
		.clock(clock),
		.io_in_a_0(r_720_0),
		.io_in_b_0(b_534_0),
		.io_in_d_0(b_1558_0),
		.io_in_control_0_dataflow(mesh_22_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2582_0),
		.io_in_last_0(r_3606_0),
		.io_in_valid_0(r_1558_0),
		.io_out_a_0(_mesh_22_16_io_out_a_0),
		.io_out_c_0(_mesh_22_16_io_out_c_0),
		.io_out_b_0(_mesh_22_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_16_io_out_id_0),
		.io_out_last_0(_mesh_22_16_io_out_last_0),
		.io_out_valid_0(_mesh_22_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10091 == GlobalFiModInstNr[0]) || (10091 == GlobalFiModInstNr[1]) || (10091 == GlobalFiModInstNr[2]) || (10091 == GlobalFiModInstNr[3]))));
	Tile mesh_22_17(
		.clock(clock),
		.io_in_a_0(r_721_0),
		.io_in_b_0(b_566_0),
		.io_in_d_0(b_1590_0),
		.io_in_control_0_dataflow(mesh_22_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2614_0),
		.io_in_last_0(r_3638_0),
		.io_in_valid_0(r_1590_0),
		.io_out_a_0(_mesh_22_17_io_out_a_0),
		.io_out_c_0(_mesh_22_17_io_out_c_0),
		.io_out_b_0(_mesh_22_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_17_io_out_id_0),
		.io_out_last_0(_mesh_22_17_io_out_last_0),
		.io_out_valid_0(_mesh_22_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10092 == GlobalFiModInstNr[0]) || (10092 == GlobalFiModInstNr[1]) || (10092 == GlobalFiModInstNr[2]) || (10092 == GlobalFiModInstNr[3]))));
	Tile mesh_22_18(
		.clock(clock),
		.io_in_a_0(r_722_0),
		.io_in_b_0(b_598_0),
		.io_in_d_0(b_1622_0),
		.io_in_control_0_dataflow(mesh_22_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2646_0),
		.io_in_last_0(r_3670_0),
		.io_in_valid_0(r_1622_0),
		.io_out_a_0(_mesh_22_18_io_out_a_0),
		.io_out_c_0(_mesh_22_18_io_out_c_0),
		.io_out_b_0(_mesh_22_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_18_io_out_id_0),
		.io_out_last_0(_mesh_22_18_io_out_last_0),
		.io_out_valid_0(_mesh_22_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10093 == GlobalFiModInstNr[0]) || (10093 == GlobalFiModInstNr[1]) || (10093 == GlobalFiModInstNr[2]) || (10093 == GlobalFiModInstNr[3]))));
	Tile mesh_22_19(
		.clock(clock),
		.io_in_a_0(r_723_0),
		.io_in_b_0(b_630_0),
		.io_in_d_0(b_1654_0),
		.io_in_control_0_dataflow(mesh_22_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2678_0),
		.io_in_last_0(r_3702_0),
		.io_in_valid_0(r_1654_0),
		.io_out_a_0(_mesh_22_19_io_out_a_0),
		.io_out_c_0(_mesh_22_19_io_out_c_0),
		.io_out_b_0(_mesh_22_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_19_io_out_id_0),
		.io_out_last_0(_mesh_22_19_io_out_last_0),
		.io_out_valid_0(_mesh_22_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10094 == GlobalFiModInstNr[0]) || (10094 == GlobalFiModInstNr[1]) || (10094 == GlobalFiModInstNr[2]) || (10094 == GlobalFiModInstNr[3]))));
	Tile mesh_22_20(
		.clock(clock),
		.io_in_a_0(r_724_0),
		.io_in_b_0(b_662_0),
		.io_in_d_0(b_1686_0),
		.io_in_control_0_dataflow(mesh_22_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2710_0),
		.io_in_last_0(r_3734_0),
		.io_in_valid_0(r_1686_0),
		.io_out_a_0(_mesh_22_20_io_out_a_0),
		.io_out_c_0(_mesh_22_20_io_out_c_0),
		.io_out_b_0(_mesh_22_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_20_io_out_id_0),
		.io_out_last_0(_mesh_22_20_io_out_last_0),
		.io_out_valid_0(_mesh_22_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10095 == GlobalFiModInstNr[0]) || (10095 == GlobalFiModInstNr[1]) || (10095 == GlobalFiModInstNr[2]) || (10095 == GlobalFiModInstNr[3]))));
	Tile mesh_22_21(
		.clock(clock),
		.io_in_a_0(r_725_0),
		.io_in_b_0(b_694_0),
		.io_in_d_0(b_1718_0),
		.io_in_control_0_dataflow(mesh_22_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2742_0),
		.io_in_last_0(r_3766_0),
		.io_in_valid_0(r_1718_0),
		.io_out_a_0(_mesh_22_21_io_out_a_0),
		.io_out_c_0(_mesh_22_21_io_out_c_0),
		.io_out_b_0(_mesh_22_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_21_io_out_id_0),
		.io_out_last_0(_mesh_22_21_io_out_last_0),
		.io_out_valid_0(_mesh_22_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10096 == GlobalFiModInstNr[0]) || (10096 == GlobalFiModInstNr[1]) || (10096 == GlobalFiModInstNr[2]) || (10096 == GlobalFiModInstNr[3]))));
	Tile mesh_22_22(
		.clock(clock),
		.io_in_a_0(r_726_0),
		.io_in_b_0(b_726_0),
		.io_in_d_0(b_1750_0),
		.io_in_control_0_dataflow(mesh_22_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2774_0),
		.io_in_last_0(r_3798_0),
		.io_in_valid_0(r_1750_0),
		.io_out_a_0(_mesh_22_22_io_out_a_0),
		.io_out_c_0(_mesh_22_22_io_out_c_0),
		.io_out_b_0(_mesh_22_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_22_io_out_id_0),
		.io_out_last_0(_mesh_22_22_io_out_last_0),
		.io_out_valid_0(_mesh_22_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10097 == GlobalFiModInstNr[0]) || (10097 == GlobalFiModInstNr[1]) || (10097 == GlobalFiModInstNr[2]) || (10097 == GlobalFiModInstNr[3]))));
	Tile mesh_22_23(
		.clock(clock),
		.io_in_a_0(r_727_0),
		.io_in_b_0(b_758_0),
		.io_in_d_0(b_1782_0),
		.io_in_control_0_dataflow(mesh_22_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2806_0),
		.io_in_last_0(r_3830_0),
		.io_in_valid_0(r_1782_0),
		.io_out_a_0(_mesh_22_23_io_out_a_0),
		.io_out_c_0(_mesh_22_23_io_out_c_0),
		.io_out_b_0(_mesh_22_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_23_io_out_id_0),
		.io_out_last_0(_mesh_22_23_io_out_last_0),
		.io_out_valid_0(_mesh_22_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10098 == GlobalFiModInstNr[0]) || (10098 == GlobalFiModInstNr[1]) || (10098 == GlobalFiModInstNr[2]) || (10098 == GlobalFiModInstNr[3]))));
	Tile mesh_22_24(
		.clock(clock),
		.io_in_a_0(r_728_0),
		.io_in_b_0(b_790_0),
		.io_in_d_0(b_1814_0),
		.io_in_control_0_dataflow(mesh_22_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2838_0),
		.io_in_last_0(r_3862_0),
		.io_in_valid_0(r_1814_0),
		.io_out_a_0(_mesh_22_24_io_out_a_0),
		.io_out_c_0(_mesh_22_24_io_out_c_0),
		.io_out_b_0(_mesh_22_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_24_io_out_id_0),
		.io_out_last_0(_mesh_22_24_io_out_last_0),
		.io_out_valid_0(_mesh_22_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10099 == GlobalFiModInstNr[0]) || (10099 == GlobalFiModInstNr[1]) || (10099 == GlobalFiModInstNr[2]) || (10099 == GlobalFiModInstNr[3]))));
	Tile mesh_22_25(
		.clock(clock),
		.io_in_a_0(r_729_0),
		.io_in_b_0(b_822_0),
		.io_in_d_0(b_1846_0),
		.io_in_control_0_dataflow(mesh_22_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2870_0),
		.io_in_last_0(r_3894_0),
		.io_in_valid_0(r_1846_0),
		.io_out_a_0(_mesh_22_25_io_out_a_0),
		.io_out_c_0(_mesh_22_25_io_out_c_0),
		.io_out_b_0(_mesh_22_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_25_io_out_id_0),
		.io_out_last_0(_mesh_22_25_io_out_last_0),
		.io_out_valid_0(_mesh_22_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10100 == GlobalFiModInstNr[0]) || (10100 == GlobalFiModInstNr[1]) || (10100 == GlobalFiModInstNr[2]) || (10100 == GlobalFiModInstNr[3]))));
	Tile mesh_22_26(
		.clock(clock),
		.io_in_a_0(r_730_0),
		.io_in_b_0(b_854_0),
		.io_in_d_0(b_1878_0),
		.io_in_control_0_dataflow(mesh_22_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2902_0),
		.io_in_last_0(r_3926_0),
		.io_in_valid_0(r_1878_0),
		.io_out_a_0(_mesh_22_26_io_out_a_0),
		.io_out_c_0(_mesh_22_26_io_out_c_0),
		.io_out_b_0(_mesh_22_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_26_io_out_id_0),
		.io_out_last_0(_mesh_22_26_io_out_last_0),
		.io_out_valid_0(_mesh_22_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10101 == GlobalFiModInstNr[0]) || (10101 == GlobalFiModInstNr[1]) || (10101 == GlobalFiModInstNr[2]) || (10101 == GlobalFiModInstNr[3]))));
	Tile mesh_22_27(
		.clock(clock),
		.io_in_a_0(r_731_0),
		.io_in_b_0(b_886_0),
		.io_in_d_0(b_1910_0),
		.io_in_control_0_dataflow(mesh_22_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2934_0),
		.io_in_last_0(r_3958_0),
		.io_in_valid_0(r_1910_0),
		.io_out_a_0(_mesh_22_27_io_out_a_0),
		.io_out_c_0(_mesh_22_27_io_out_c_0),
		.io_out_b_0(_mesh_22_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_27_io_out_id_0),
		.io_out_last_0(_mesh_22_27_io_out_last_0),
		.io_out_valid_0(_mesh_22_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10102 == GlobalFiModInstNr[0]) || (10102 == GlobalFiModInstNr[1]) || (10102 == GlobalFiModInstNr[2]) || (10102 == GlobalFiModInstNr[3]))));
	Tile mesh_22_28(
		.clock(clock),
		.io_in_a_0(r_732_0),
		.io_in_b_0(b_918_0),
		.io_in_d_0(b_1942_0),
		.io_in_control_0_dataflow(mesh_22_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2966_0),
		.io_in_last_0(r_3990_0),
		.io_in_valid_0(r_1942_0),
		.io_out_a_0(_mesh_22_28_io_out_a_0),
		.io_out_c_0(_mesh_22_28_io_out_c_0),
		.io_out_b_0(_mesh_22_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_28_io_out_id_0),
		.io_out_last_0(_mesh_22_28_io_out_last_0),
		.io_out_valid_0(_mesh_22_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10103 == GlobalFiModInstNr[0]) || (10103 == GlobalFiModInstNr[1]) || (10103 == GlobalFiModInstNr[2]) || (10103 == GlobalFiModInstNr[3]))));
	Tile mesh_22_29(
		.clock(clock),
		.io_in_a_0(r_733_0),
		.io_in_b_0(b_950_0),
		.io_in_d_0(b_1974_0),
		.io_in_control_0_dataflow(mesh_22_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2998_0),
		.io_in_last_0(r_4022_0),
		.io_in_valid_0(r_1974_0),
		.io_out_a_0(_mesh_22_29_io_out_a_0),
		.io_out_c_0(_mesh_22_29_io_out_c_0),
		.io_out_b_0(_mesh_22_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_29_io_out_id_0),
		.io_out_last_0(_mesh_22_29_io_out_last_0),
		.io_out_valid_0(_mesh_22_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10104 == GlobalFiModInstNr[0]) || (10104 == GlobalFiModInstNr[1]) || (10104 == GlobalFiModInstNr[2]) || (10104 == GlobalFiModInstNr[3]))));
	Tile mesh_22_30(
		.clock(clock),
		.io_in_a_0(r_734_0),
		.io_in_b_0(b_982_0),
		.io_in_d_0(b_2006_0),
		.io_in_control_0_dataflow(mesh_22_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3030_0),
		.io_in_last_0(r_4054_0),
		.io_in_valid_0(r_2006_0),
		.io_out_a_0(_mesh_22_30_io_out_a_0),
		.io_out_c_0(_mesh_22_30_io_out_c_0),
		.io_out_b_0(_mesh_22_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_30_io_out_id_0),
		.io_out_last_0(_mesh_22_30_io_out_last_0),
		.io_out_valid_0(_mesh_22_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10105 == GlobalFiModInstNr[0]) || (10105 == GlobalFiModInstNr[1]) || (10105 == GlobalFiModInstNr[2]) || (10105 == GlobalFiModInstNr[3]))));
	Tile mesh_22_31(
		.clock(clock),
		.io_in_a_0(r_735_0),
		.io_in_b_0(b_1014_0),
		.io_in_d_0(b_2038_0),
		.io_in_control_0_dataflow(mesh_22_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_22_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_22_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3062_0),
		.io_in_last_0(r_4086_0),
		.io_in_valid_0(r_2038_0),
		.io_out_a_0(_mesh_22_31_io_out_a_0),
		.io_out_c_0(_mesh_22_31_io_out_c_0),
		.io_out_b_0(_mesh_22_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_22_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_22_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_22_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_22_31_io_out_id_0),
		.io_out_last_0(_mesh_22_31_io_out_last_0),
		.io_out_valid_0(_mesh_22_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10106 == GlobalFiModInstNr[0]) || (10106 == GlobalFiModInstNr[1]) || (10106 == GlobalFiModInstNr[2]) || (10106 == GlobalFiModInstNr[3]))));
	Tile mesh_23_0(
		.clock(clock),
		.io_in_a_0(r_736_0),
		.io_in_b_0(b_23_0),
		.io_in_d_0(b_1047_0),
		.io_in_control_0_dataflow(mesh_23_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2071_0),
		.io_in_last_0(r_3095_0),
		.io_in_valid_0(r_1047_0),
		.io_out_a_0(_mesh_23_0_io_out_a_0),
		.io_out_c_0(_mesh_23_0_io_out_c_0),
		.io_out_b_0(_mesh_23_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_0_io_out_id_0),
		.io_out_last_0(_mesh_23_0_io_out_last_0),
		.io_out_valid_0(_mesh_23_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10107 == GlobalFiModInstNr[0]) || (10107 == GlobalFiModInstNr[1]) || (10107 == GlobalFiModInstNr[2]) || (10107 == GlobalFiModInstNr[3]))));
	Tile mesh_23_1(
		.clock(clock),
		.io_in_a_0(r_737_0),
		.io_in_b_0(b_55_0),
		.io_in_d_0(b_1079_0),
		.io_in_control_0_dataflow(mesh_23_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2103_0),
		.io_in_last_0(r_3127_0),
		.io_in_valid_0(r_1079_0),
		.io_out_a_0(_mesh_23_1_io_out_a_0),
		.io_out_c_0(_mesh_23_1_io_out_c_0),
		.io_out_b_0(_mesh_23_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_1_io_out_id_0),
		.io_out_last_0(_mesh_23_1_io_out_last_0),
		.io_out_valid_0(_mesh_23_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10108 == GlobalFiModInstNr[0]) || (10108 == GlobalFiModInstNr[1]) || (10108 == GlobalFiModInstNr[2]) || (10108 == GlobalFiModInstNr[3]))));
	Tile mesh_23_2(
		.clock(clock),
		.io_in_a_0(r_738_0),
		.io_in_b_0(b_87_0),
		.io_in_d_0(b_1111_0),
		.io_in_control_0_dataflow(mesh_23_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2135_0),
		.io_in_last_0(r_3159_0),
		.io_in_valid_0(r_1111_0),
		.io_out_a_0(_mesh_23_2_io_out_a_0),
		.io_out_c_0(_mesh_23_2_io_out_c_0),
		.io_out_b_0(_mesh_23_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_2_io_out_id_0),
		.io_out_last_0(_mesh_23_2_io_out_last_0),
		.io_out_valid_0(_mesh_23_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10109 == GlobalFiModInstNr[0]) || (10109 == GlobalFiModInstNr[1]) || (10109 == GlobalFiModInstNr[2]) || (10109 == GlobalFiModInstNr[3]))));
	Tile mesh_23_3(
		.clock(clock),
		.io_in_a_0(r_739_0),
		.io_in_b_0(b_119_0),
		.io_in_d_0(b_1143_0),
		.io_in_control_0_dataflow(mesh_23_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2167_0),
		.io_in_last_0(r_3191_0),
		.io_in_valid_0(r_1143_0),
		.io_out_a_0(_mesh_23_3_io_out_a_0),
		.io_out_c_0(_mesh_23_3_io_out_c_0),
		.io_out_b_0(_mesh_23_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_3_io_out_id_0),
		.io_out_last_0(_mesh_23_3_io_out_last_0),
		.io_out_valid_0(_mesh_23_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10110 == GlobalFiModInstNr[0]) || (10110 == GlobalFiModInstNr[1]) || (10110 == GlobalFiModInstNr[2]) || (10110 == GlobalFiModInstNr[3]))));
	Tile mesh_23_4(
		.clock(clock),
		.io_in_a_0(r_740_0),
		.io_in_b_0(b_151_0),
		.io_in_d_0(b_1175_0),
		.io_in_control_0_dataflow(mesh_23_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2199_0),
		.io_in_last_0(r_3223_0),
		.io_in_valid_0(r_1175_0),
		.io_out_a_0(_mesh_23_4_io_out_a_0),
		.io_out_c_0(_mesh_23_4_io_out_c_0),
		.io_out_b_0(_mesh_23_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_4_io_out_id_0),
		.io_out_last_0(_mesh_23_4_io_out_last_0),
		.io_out_valid_0(_mesh_23_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10111 == GlobalFiModInstNr[0]) || (10111 == GlobalFiModInstNr[1]) || (10111 == GlobalFiModInstNr[2]) || (10111 == GlobalFiModInstNr[3]))));
	Tile mesh_23_5(
		.clock(clock),
		.io_in_a_0(r_741_0),
		.io_in_b_0(b_183_0),
		.io_in_d_0(b_1207_0),
		.io_in_control_0_dataflow(mesh_23_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2231_0),
		.io_in_last_0(r_3255_0),
		.io_in_valid_0(r_1207_0),
		.io_out_a_0(_mesh_23_5_io_out_a_0),
		.io_out_c_0(_mesh_23_5_io_out_c_0),
		.io_out_b_0(_mesh_23_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_5_io_out_id_0),
		.io_out_last_0(_mesh_23_5_io_out_last_0),
		.io_out_valid_0(_mesh_23_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10112 == GlobalFiModInstNr[0]) || (10112 == GlobalFiModInstNr[1]) || (10112 == GlobalFiModInstNr[2]) || (10112 == GlobalFiModInstNr[3]))));
	Tile mesh_23_6(
		.clock(clock),
		.io_in_a_0(r_742_0),
		.io_in_b_0(b_215_0),
		.io_in_d_0(b_1239_0),
		.io_in_control_0_dataflow(mesh_23_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2263_0),
		.io_in_last_0(r_3287_0),
		.io_in_valid_0(r_1239_0),
		.io_out_a_0(_mesh_23_6_io_out_a_0),
		.io_out_c_0(_mesh_23_6_io_out_c_0),
		.io_out_b_0(_mesh_23_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_6_io_out_id_0),
		.io_out_last_0(_mesh_23_6_io_out_last_0),
		.io_out_valid_0(_mesh_23_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10113 == GlobalFiModInstNr[0]) || (10113 == GlobalFiModInstNr[1]) || (10113 == GlobalFiModInstNr[2]) || (10113 == GlobalFiModInstNr[3]))));
	Tile mesh_23_7(
		.clock(clock),
		.io_in_a_0(r_743_0),
		.io_in_b_0(b_247_0),
		.io_in_d_0(b_1271_0),
		.io_in_control_0_dataflow(mesh_23_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2295_0),
		.io_in_last_0(r_3319_0),
		.io_in_valid_0(r_1271_0),
		.io_out_a_0(_mesh_23_7_io_out_a_0),
		.io_out_c_0(_mesh_23_7_io_out_c_0),
		.io_out_b_0(_mesh_23_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_7_io_out_id_0),
		.io_out_last_0(_mesh_23_7_io_out_last_0),
		.io_out_valid_0(_mesh_23_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10114 == GlobalFiModInstNr[0]) || (10114 == GlobalFiModInstNr[1]) || (10114 == GlobalFiModInstNr[2]) || (10114 == GlobalFiModInstNr[3]))));
	Tile mesh_23_8(
		.clock(clock),
		.io_in_a_0(r_744_0),
		.io_in_b_0(b_279_0),
		.io_in_d_0(b_1303_0),
		.io_in_control_0_dataflow(mesh_23_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2327_0),
		.io_in_last_0(r_3351_0),
		.io_in_valid_0(r_1303_0),
		.io_out_a_0(_mesh_23_8_io_out_a_0),
		.io_out_c_0(_mesh_23_8_io_out_c_0),
		.io_out_b_0(_mesh_23_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_8_io_out_id_0),
		.io_out_last_0(_mesh_23_8_io_out_last_0),
		.io_out_valid_0(_mesh_23_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10115 == GlobalFiModInstNr[0]) || (10115 == GlobalFiModInstNr[1]) || (10115 == GlobalFiModInstNr[2]) || (10115 == GlobalFiModInstNr[3]))));
	Tile mesh_23_9(
		.clock(clock),
		.io_in_a_0(r_745_0),
		.io_in_b_0(b_311_0),
		.io_in_d_0(b_1335_0),
		.io_in_control_0_dataflow(mesh_23_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2359_0),
		.io_in_last_0(r_3383_0),
		.io_in_valid_0(r_1335_0),
		.io_out_a_0(_mesh_23_9_io_out_a_0),
		.io_out_c_0(_mesh_23_9_io_out_c_0),
		.io_out_b_0(_mesh_23_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_9_io_out_id_0),
		.io_out_last_0(_mesh_23_9_io_out_last_0),
		.io_out_valid_0(_mesh_23_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10116 == GlobalFiModInstNr[0]) || (10116 == GlobalFiModInstNr[1]) || (10116 == GlobalFiModInstNr[2]) || (10116 == GlobalFiModInstNr[3]))));
	Tile mesh_23_10(
		.clock(clock),
		.io_in_a_0(r_746_0),
		.io_in_b_0(b_343_0),
		.io_in_d_0(b_1367_0),
		.io_in_control_0_dataflow(mesh_23_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2391_0),
		.io_in_last_0(r_3415_0),
		.io_in_valid_0(r_1367_0),
		.io_out_a_0(_mesh_23_10_io_out_a_0),
		.io_out_c_0(_mesh_23_10_io_out_c_0),
		.io_out_b_0(_mesh_23_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_10_io_out_id_0),
		.io_out_last_0(_mesh_23_10_io_out_last_0),
		.io_out_valid_0(_mesh_23_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10117 == GlobalFiModInstNr[0]) || (10117 == GlobalFiModInstNr[1]) || (10117 == GlobalFiModInstNr[2]) || (10117 == GlobalFiModInstNr[3]))));
	Tile mesh_23_11(
		.clock(clock),
		.io_in_a_0(r_747_0),
		.io_in_b_0(b_375_0),
		.io_in_d_0(b_1399_0),
		.io_in_control_0_dataflow(mesh_23_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2423_0),
		.io_in_last_0(r_3447_0),
		.io_in_valid_0(r_1399_0),
		.io_out_a_0(_mesh_23_11_io_out_a_0),
		.io_out_c_0(_mesh_23_11_io_out_c_0),
		.io_out_b_0(_mesh_23_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_11_io_out_id_0),
		.io_out_last_0(_mesh_23_11_io_out_last_0),
		.io_out_valid_0(_mesh_23_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10118 == GlobalFiModInstNr[0]) || (10118 == GlobalFiModInstNr[1]) || (10118 == GlobalFiModInstNr[2]) || (10118 == GlobalFiModInstNr[3]))));
	Tile mesh_23_12(
		.clock(clock),
		.io_in_a_0(r_748_0),
		.io_in_b_0(b_407_0),
		.io_in_d_0(b_1431_0),
		.io_in_control_0_dataflow(mesh_23_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2455_0),
		.io_in_last_0(r_3479_0),
		.io_in_valid_0(r_1431_0),
		.io_out_a_0(_mesh_23_12_io_out_a_0),
		.io_out_c_0(_mesh_23_12_io_out_c_0),
		.io_out_b_0(_mesh_23_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_12_io_out_id_0),
		.io_out_last_0(_mesh_23_12_io_out_last_0),
		.io_out_valid_0(_mesh_23_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10119 == GlobalFiModInstNr[0]) || (10119 == GlobalFiModInstNr[1]) || (10119 == GlobalFiModInstNr[2]) || (10119 == GlobalFiModInstNr[3]))));
	Tile mesh_23_13(
		.clock(clock),
		.io_in_a_0(r_749_0),
		.io_in_b_0(b_439_0),
		.io_in_d_0(b_1463_0),
		.io_in_control_0_dataflow(mesh_23_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2487_0),
		.io_in_last_0(r_3511_0),
		.io_in_valid_0(r_1463_0),
		.io_out_a_0(_mesh_23_13_io_out_a_0),
		.io_out_c_0(_mesh_23_13_io_out_c_0),
		.io_out_b_0(_mesh_23_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_13_io_out_id_0),
		.io_out_last_0(_mesh_23_13_io_out_last_0),
		.io_out_valid_0(_mesh_23_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10120 == GlobalFiModInstNr[0]) || (10120 == GlobalFiModInstNr[1]) || (10120 == GlobalFiModInstNr[2]) || (10120 == GlobalFiModInstNr[3]))));
	Tile mesh_23_14(
		.clock(clock),
		.io_in_a_0(r_750_0),
		.io_in_b_0(b_471_0),
		.io_in_d_0(b_1495_0),
		.io_in_control_0_dataflow(mesh_23_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2519_0),
		.io_in_last_0(r_3543_0),
		.io_in_valid_0(r_1495_0),
		.io_out_a_0(_mesh_23_14_io_out_a_0),
		.io_out_c_0(_mesh_23_14_io_out_c_0),
		.io_out_b_0(_mesh_23_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_14_io_out_id_0),
		.io_out_last_0(_mesh_23_14_io_out_last_0),
		.io_out_valid_0(_mesh_23_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10121 == GlobalFiModInstNr[0]) || (10121 == GlobalFiModInstNr[1]) || (10121 == GlobalFiModInstNr[2]) || (10121 == GlobalFiModInstNr[3]))));
	Tile mesh_23_15(
		.clock(clock),
		.io_in_a_0(r_751_0),
		.io_in_b_0(b_503_0),
		.io_in_d_0(b_1527_0),
		.io_in_control_0_dataflow(mesh_23_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2551_0),
		.io_in_last_0(r_3575_0),
		.io_in_valid_0(r_1527_0),
		.io_out_a_0(_mesh_23_15_io_out_a_0),
		.io_out_c_0(_mesh_23_15_io_out_c_0),
		.io_out_b_0(_mesh_23_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_15_io_out_id_0),
		.io_out_last_0(_mesh_23_15_io_out_last_0),
		.io_out_valid_0(_mesh_23_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10122 == GlobalFiModInstNr[0]) || (10122 == GlobalFiModInstNr[1]) || (10122 == GlobalFiModInstNr[2]) || (10122 == GlobalFiModInstNr[3]))));
	Tile mesh_23_16(
		.clock(clock),
		.io_in_a_0(r_752_0),
		.io_in_b_0(b_535_0),
		.io_in_d_0(b_1559_0),
		.io_in_control_0_dataflow(mesh_23_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2583_0),
		.io_in_last_0(r_3607_0),
		.io_in_valid_0(r_1559_0),
		.io_out_a_0(_mesh_23_16_io_out_a_0),
		.io_out_c_0(_mesh_23_16_io_out_c_0),
		.io_out_b_0(_mesh_23_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_16_io_out_id_0),
		.io_out_last_0(_mesh_23_16_io_out_last_0),
		.io_out_valid_0(_mesh_23_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10123 == GlobalFiModInstNr[0]) || (10123 == GlobalFiModInstNr[1]) || (10123 == GlobalFiModInstNr[2]) || (10123 == GlobalFiModInstNr[3]))));
	Tile mesh_23_17(
		.clock(clock),
		.io_in_a_0(r_753_0),
		.io_in_b_0(b_567_0),
		.io_in_d_0(b_1591_0),
		.io_in_control_0_dataflow(mesh_23_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2615_0),
		.io_in_last_0(r_3639_0),
		.io_in_valid_0(r_1591_0),
		.io_out_a_0(_mesh_23_17_io_out_a_0),
		.io_out_c_0(_mesh_23_17_io_out_c_0),
		.io_out_b_0(_mesh_23_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_17_io_out_id_0),
		.io_out_last_0(_mesh_23_17_io_out_last_0),
		.io_out_valid_0(_mesh_23_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10124 == GlobalFiModInstNr[0]) || (10124 == GlobalFiModInstNr[1]) || (10124 == GlobalFiModInstNr[2]) || (10124 == GlobalFiModInstNr[3]))));
	Tile mesh_23_18(
		.clock(clock),
		.io_in_a_0(r_754_0),
		.io_in_b_0(b_599_0),
		.io_in_d_0(b_1623_0),
		.io_in_control_0_dataflow(mesh_23_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2647_0),
		.io_in_last_0(r_3671_0),
		.io_in_valid_0(r_1623_0),
		.io_out_a_0(_mesh_23_18_io_out_a_0),
		.io_out_c_0(_mesh_23_18_io_out_c_0),
		.io_out_b_0(_mesh_23_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_18_io_out_id_0),
		.io_out_last_0(_mesh_23_18_io_out_last_0),
		.io_out_valid_0(_mesh_23_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10125 == GlobalFiModInstNr[0]) || (10125 == GlobalFiModInstNr[1]) || (10125 == GlobalFiModInstNr[2]) || (10125 == GlobalFiModInstNr[3]))));
	Tile mesh_23_19(
		.clock(clock),
		.io_in_a_0(r_755_0),
		.io_in_b_0(b_631_0),
		.io_in_d_0(b_1655_0),
		.io_in_control_0_dataflow(mesh_23_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2679_0),
		.io_in_last_0(r_3703_0),
		.io_in_valid_0(r_1655_0),
		.io_out_a_0(_mesh_23_19_io_out_a_0),
		.io_out_c_0(_mesh_23_19_io_out_c_0),
		.io_out_b_0(_mesh_23_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_19_io_out_id_0),
		.io_out_last_0(_mesh_23_19_io_out_last_0),
		.io_out_valid_0(_mesh_23_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10126 == GlobalFiModInstNr[0]) || (10126 == GlobalFiModInstNr[1]) || (10126 == GlobalFiModInstNr[2]) || (10126 == GlobalFiModInstNr[3]))));
	Tile mesh_23_20(
		.clock(clock),
		.io_in_a_0(r_756_0),
		.io_in_b_0(b_663_0),
		.io_in_d_0(b_1687_0),
		.io_in_control_0_dataflow(mesh_23_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2711_0),
		.io_in_last_0(r_3735_0),
		.io_in_valid_0(r_1687_0),
		.io_out_a_0(_mesh_23_20_io_out_a_0),
		.io_out_c_0(_mesh_23_20_io_out_c_0),
		.io_out_b_0(_mesh_23_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_20_io_out_id_0),
		.io_out_last_0(_mesh_23_20_io_out_last_0),
		.io_out_valid_0(_mesh_23_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10127 == GlobalFiModInstNr[0]) || (10127 == GlobalFiModInstNr[1]) || (10127 == GlobalFiModInstNr[2]) || (10127 == GlobalFiModInstNr[3]))));
	Tile mesh_23_21(
		.clock(clock),
		.io_in_a_0(r_757_0),
		.io_in_b_0(b_695_0),
		.io_in_d_0(b_1719_0),
		.io_in_control_0_dataflow(mesh_23_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2743_0),
		.io_in_last_0(r_3767_0),
		.io_in_valid_0(r_1719_0),
		.io_out_a_0(_mesh_23_21_io_out_a_0),
		.io_out_c_0(_mesh_23_21_io_out_c_0),
		.io_out_b_0(_mesh_23_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_21_io_out_id_0),
		.io_out_last_0(_mesh_23_21_io_out_last_0),
		.io_out_valid_0(_mesh_23_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10128 == GlobalFiModInstNr[0]) || (10128 == GlobalFiModInstNr[1]) || (10128 == GlobalFiModInstNr[2]) || (10128 == GlobalFiModInstNr[3]))));
	Tile mesh_23_22(
		.clock(clock),
		.io_in_a_0(r_758_0),
		.io_in_b_0(b_727_0),
		.io_in_d_0(b_1751_0),
		.io_in_control_0_dataflow(mesh_23_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2775_0),
		.io_in_last_0(r_3799_0),
		.io_in_valid_0(r_1751_0),
		.io_out_a_0(_mesh_23_22_io_out_a_0),
		.io_out_c_0(_mesh_23_22_io_out_c_0),
		.io_out_b_0(_mesh_23_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_22_io_out_id_0),
		.io_out_last_0(_mesh_23_22_io_out_last_0),
		.io_out_valid_0(_mesh_23_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10129 == GlobalFiModInstNr[0]) || (10129 == GlobalFiModInstNr[1]) || (10129 == GlobalFiModInstNr[2]) || (10129 == GlobalFiModInstNr[3]))));
	Tile mesh_23_23(
		.clock(clock),
		.io_in_a_0(r_759_0),
		.io_in_b_0(b_759_0),
		.io_in_d_0(b_1783_0),
		.io_in_control_0_dataflow(mesh_23_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2807_0),
		.io_in_last_0(r_3831_0),
		.io_in_valid_0(r_1783_0),
		.io_out_a_0(_mesh_23_23_io_out_a_0),
		.io_out_c_0(_mesh_23_23_io_out_c_0),
		.io_out_b_0(_mesh_23_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_23_io_out_id_0),
		.io_out_last_0(_mesh_23_23_io_out_last_0),
		.io_out_valid_0(_mesh_23_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10130 == GlobalFiModInstNr[0]) || (10130 == GlobalFiModInstNr[1]) || (10130 == GlobalFiModInstNr[2]) || (10130 == GlobalFiModInstNr[3]))));
	Tile mesh_23_24(
		.clock(clock),
		.io_in_a_0(r_760_0),
		.io_in_b_0(b_791_0),
		.io_in_d_0(b_1815_0),
		.io_in_control_0_dataflow(mesh_23_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2839_0),
		.io_in_last_0(r_3863_0),
		.io_in_valid_0(r_1815_0),
		.io_out_a_0(_mesh_23_24_io_out_a_0),
		.io_out_c_0(_mesh_23_24_io_out_c_0),
		.io_out_b_0(_mesh_23_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_24_io_out_id_0),
		.io_out_last_0(_mesh_23_24_io_out_last_0),
		.io_out_valid_0(_mesh_23_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10131 == GlobalFiModInstNr[0]) || (10131 == GlobalFiModInstNr[1]) || (10131 == GlobalFiModInstNr[2]) || (10131 == GlobalFiModInstNr[3]))));
	Tile mesh_23_25(
		.clock(clock),
		.io_in_a_0(r_761_0),
		.io_in_b_0(b_823_0),
		.io_in_d_0(b_1847_0),
		.io_in_control_0_dataflow(mesh_23_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2871_0),
		.io_in_last_0(r_3895_0),
		.io_in_valid_0(r_1847_0),
		.io_out_a_0(_mesh_23_25_io_out_a_0),
		.io_out_c_0(_mesh_23_25_io_out_c_0),
		.io_out_b_0(_mesh_23_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_25_io_out_id_0),
		.io_out_last_0(_mesh_23_25_io_out_last_0),
		.io_out_valid_0(_mesh_23_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10132 == GlobalFiModInstNr[0]) || (10132 == GlobalFiModInstNr[1]) || (10132 == GlobalFiModInstNr[2]) || (10132 == GlobalFiModInstNr[3]))));
	Tile mesh_23_26(
		.clock(clock),
		.io_in_a_0(r_762_0),
		.io_in_b_0(b_855_0),
		.io_in_d_0(b_1879_0),
		.io_in_control_0_dataflow(mesh_23_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2903_0),
		.io_in_last_0(r_3927_0),
		.io_in_valid_0(r_1879_0),
		.io_out_a_0(_mesh_23_26_io_out_a_0),
		.io_out_c_0(_mesh_23_26_io_out_c_0),
		.io_out_b_0(_mesh_23_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_26_io_out_id_0),
		.io_out_last_0(_mesh_23_26_io_out_last_0),
		.io_out_valid_0(_mesh_23_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10133 == GlobalFiModInstNr[0]) || (10133 == GlobalFiModInstNr[1]) || (10133 == GlobalFiModInstNr[2]) || (10133 == GlobalFiModInstNr[3]))));
	Tile mesh_23_27(
		.clock(clock),
		.io_in_a_0(r_763_0),
		.io_in_b_0(b_887_0),
		.io_in_d_0(b_1911_0),
		.io_in_control_0_dataflow(mesh_23_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2935_0),
		.io_in_last_0(r_3959_0),
		.io_in_valid_0(r_1911_0),
		.io_out_a_0(_mesh_23_27_io_out_a_0),
		.io_out_c_0(_mesh_23_27_io_out_c_0),
		.io_out_b_0(_mesh_23_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_27_io_out_id_0),
		.io_out_last_0(_mesh_23_27_io_out_last_0),
		.io_out_valid_0(_mesh_23_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10134 == GlobalFiModInstNr[0]) || (10134 == GlobalFiModInstNr[1]) || (10134 == GlobalFiModInstNr[2]) || (10134 == GlobalFiModInstNr[3]))));
	Tile mesh_23_28(
		.clock(clock),
		.io_in_a_0(r_764_0),
		.io_in_b_0(b_919_0),
		.io_in_d_0(b_1943_0),
		.io_in_control_0_dataflow(mesh_23_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2967_0),
		.io_in_last_0(r_3991_0),
		.io_in_valid_0(r_1943_0),
		.io_out_a_0(_mesh_23_28_io_out_a_0),
		.io_out_c_0(_mesh_23_28_io_out_c_0),
		.io_out_b_0(_mesh_23_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_28_io_out_id_0),
		.io_out_last_0(_mesh_23_28_io_out_last_0),
		.io_out_valid_0(_mesh_23_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10135 == GlobalFiModInstNr[0]) || (10135 == GlobalFiModInstNr[1]) || (10135 == GlobalFiModInstNr[2]) || (10135 == GlobalFiModInstNr[3]))));
	Tile mesh_23_29(
		.clock(clock),
		.io_in_a_0(r_765_0),
		.io_in_b_0(b_951_0),
		.io_in_d_0(b_1975_0),
		.io_in_control_0_dataflow(mesh_23_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_29_io_in_control_0_shift_b),
		.io_in_id_0(r_2999_0),
		.io_in_last_0(r_4023_0),
		.io_in_valid_0(r_1975_0),
		.io_out_a_0(_mesh_23_29_io_out_a_0),
		.io_out_c_0(_mesh_23_29_io_out_c_0),
		.io_out_b_0(_mesh_23_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_29_io_out_id_0),
		.io_out_last_0(_mesh_23_29_io_out_last_0),
		.io_out_valid_0(_mesh_23_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10136 == GlobalFiModInstNr[0]) || (10136 == GlobalFiModInstNr[1]) || (10136 == GlobalFiModInstNr[2]) || (10136 == GlobalFiModInstNr[3]))));
	Tile mesh_23_30(
		.clock(clock),
		.io_in_a_0(r_766_0),
		.io_in_b_0(b_983_0),
		.io_in_d_0(b_2007_0),
		.io_in_control_0_dataflow(mesh_23_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3031_0),
		.io_in_last_0(r_4055_0),
		.io_in_valid_0(r_2007_0),
		.io_out_a_0(_mesh_23_30_io_out_a_0),
		.io_out_c_0(_mesh_23_30_io_out_c_0),
		.io_out_b_0(_mesh_23_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_30_io_out_id_0),
		.io_out_last_0(_mesh_23_30_io_out_last_0),
		.io_out_valid_0(_mesh_23_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10137 == GlobalFiModInstNr[0]) || (10137 == GlobalFiModInstNr[1]) || (10137 == GlobalFiModInstNr[2]) || (10137 == GlobalFiModInstNr[3]))));
	Tile mesh_23_31(
		.clock(clock),
		.io_in_a_0(r_767_0),
		.io_in_b_0(b_1015_0),
		.io_in_d_0(b_2039_0),
		.io_in_control_0_dataflow(mesh_23_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_23_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_23_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3063_0),
		.io_in_last_0(r_4087_0),
		.io_in_valid_0(r_2039_0),
		.io_out_a_0(_mesh_23_31_io_out_a_0),
		.io_out_c_0(_mesh_23_31_io_out_c_0),
		.io_out_b_0(_mesh_23_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_23_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_23_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_23_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_23_31_io_out_id_0),
		.io_out_last_0(_mesh_23_31_io_out_last_0),
		.io_out_valid_0(_mesh_23_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10138 == GlobalFiModInstNr[0]) || (10138 == GlobalFiModInstNr[1]) || (10138 == GlobalFiModInstNr[2]) || (10138 == GlobalFiModInstNr[3]))));
	Tile mesh_24_0(
		.clock(clock),
		.io_in_a_0(r_768_0),
		.io_in_b_0(b_24_0),
		.io_in_d_0(b_1048_0),
		.io_in_control_0_dataflow(mesh_24_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2072_0),
		.io_in_last_0(r_3096_0),
		.io_in_valid_0(r_1048_0),
		.io_out_a_0(_mesh_24_0_io_out_a_0),
		.io_out_c_0(_mesh_24_0_io_out_c_0),
		.io_out_b_0(_mesh_24_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_0_io_out_id_0),
		.io_out_last_0(_mesh_24_0_io_out_last_0),
		.io_out_valid_0(_mesh_24_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10139 == GlobalFiModInstNr[0]) || (10139 == GlobalFiModInstNr[1]) || (10139 == GlobalFiModInstNr[2]) || (10139 == GlobalFiModInstNr[3]))));
	Tile mesh_24_1(
		.clock(clock),
		.io_in_a_0(r_769_0),
		.io_in_b_0(b_56_0),
		.io_in_d_0(b_1080_0),
		.io_in_control_0_dataflow(mesh_24_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2104_0),
		.io_in_last_0(r_3128_0),
		.io_in_valid_0(r_1080_0),
		.io_out_a_0(_mesh_24_1_io_out_a_0),
		.io_out_c_0(_mesh_24_1_io_out_c_0),
		.io_out_b_0(_mesh_24_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_1_io_out_id_0),
		.io_out_last_0(_mesh_24_1_io_out_last_0),
		.io_out_valid_0(_mesh_24_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10140 == GlobalFiModInstNr[0]) || (10140 == GlobalFiModInstNr[1]) || (10140 == GlobalFiModInstNr[2]) || (10140 == GlobalFiModInstNr[3]))));
	Tile mesh_24_2(
		.clock(clock),
		.io_in_a_0(r_770_0),
		.io_in_b_0(b_88_0),
		.io_in_d_0(b_1112_0),
		.io_in_control_0_dataflow(mesh_24_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2136_0),
		.io_in_last_0(r_3160_0),
		.io_in_valid_0(r_1112_0),
		.io_out_a_0(_mesh_24_2_io_out_a_0),
		.io_out_c_0(_mesh_24_2_io_out_c_0),
		.io_out_b_0(_mesh_24_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_2_io_out_id_0),
		.io_out_last_0(_mesh_24_2_io_out_last_0),
		.io_out_valid_0(_mesh_24_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10141 == GlobalFiModInstNr[0]) || (10141 == GlobalFiModInstNr[1]) || (10141 == GlobalFiModInstNr[2]) || (10141 == GlobalFiModInstNr[3]))));
	Tile mesh_24_3(
		.clock(clock),
		.io_in_a_0(r_771_0),
		.io_in_b_0(b_120_0),
		.io_in_d_0(b_1144_0),
		.io_in_control_0_dataflow(mesh_24_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2168_0),
		.io_in_last_0(r_3192_0),
		.io_in_valid_0(r_1144_0),
		.io_out_a_0(_mesh_24_3_io_out_a_0),
		.io_out_c_0(_mesh_24_3_io_out_c_0),
		.io_out_b_0(_mesh_24_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_3_io_out_id_0),
		.io_out_last_0(_mesh_24_3_io_out_last_0),
		.io_out_valid_0(_mesh_24_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10142 == GlobalFiModInstNr[0]) || (10142 == GlobalFiModInstNr[1]) || (10142 == GlobalFiModInstNr[2]) || (10142 == GlobalFiModInstNr[3]))));
	Tile mesh_24_4(
		.clock(clock),
		.io_in_a_0(r_772_0),
		.io_in_b_0(b_152_0),
		.io_in_d_0(b_1176_0),
		.io_in_control_0_dataflow(mesh_24_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2200_0),
		.io_in_last_0(r_3224_0),
		.io_in_valid_0(r_1176_0),
		.io_out_a_0(_mesh_24_4_io_out_a_0),
		.io_out_c_0(_mesh_24_4_io_out_c_0),
		.io_out_b_0(_mesh_24_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_4_io_out_id_0),
		.io_out_last_0(_mesh_24_4_io_out_last_0),
		.io_out_valid_0(_mesh_24_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10143 == GlobalFiModInstNr[0]) || (10143 == GlobalFiModInstNr[1]) || (10143 == GlobalFiModInstNr[2]) || (10143 == GlobalFiModInstNr[3]))));
	Tile mesh_24_5(
		.clock(clock),
		.io_in_a_0(r_773_0),
		.io_in_b_0(b_184_0),
		.io_in_d_0(b_1208_0),
		.io_in_control_0_dataflow(mesh_24_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2232_0),
		.io_in_last_0(r_3256_0),
		.io_in_valid_0(r_1208_0),
		.io_out_a_0(_mesh_24_5_io_out_a_0),
		.io_out_c_0(_mesh_24_5_io_out_c_0),
		.io_out_b_0(_mesh_24_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_5_io_out_id_0),
		.io_out_last_0(_mesh_24_5_io_out_last_0),
		.io_out_valid_0(_mesh_24_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10144 == GlobalFiModInstNr[0]) || (10144 == GlobalFiModInstNr[1]) || (10144 == GlobalFiModInstNr[2]) || (10144 == GlobalFiModInstNr[3]))));
	Tile mesh_24_6(
		.clock(clock),
		.io_in_a_0(r_774_0),
		.io_in_b_0(b_216_0),
		.io_in_d_0(b_1240_0),
		.io_in_control_0_dataflow(mesh_24_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2264_0),
		.io_in_last_0(r_3288_0),
		.io_in_valid_0(r_1240_0),
		.io_out_a_0(_mesh_24_6_io_out_a_0),
		.io_out_c_0(_mesh_24_6_io_out_c_0),
		.io_out_b_0(_mesh_24_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_6_io_out_id_0),
		.io_out_last_0(_mesh_24_6_io_out_last_0),
		.io_out_valid_0(_mesh_24_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10145 == GlobalFiModInstNr[0]) || (10145 == GlobalFiModInstNr[1]) || (10145 == GlobalFiModInstNr[2]) || (10145 == GlobalFiModInstNr[3]))));
	Tile mesh_24_7(
		.clock(clock),
		.io_in_a_0(r_775_0),
		.io_in_b_0(b_248_0),
		.io_in_d_0(b_1272_0),
		.io_in_control_0_dataflow(mesh_24_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2296_0),
		.io_in_last_0(r_3320_0),
		.io_in_valid_0(r_1272_0),
		.io_out_a_0(_mesh_24_7_io_out_a_0),
		.io_out_c_0(_mesh_24_7_io_out_c_0),
		.io_out_b_0(_mesh_24_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_7_io_out_id_0),
		.io_out_last_0(_mesh_24_7_io_out_last_0),
		.io_out_valid_0(_mesh_24_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10146 == GlobalFiModInstNr[0]) || (10146 == GlobalFiModInstNr[1]) || (10146 == GlobalFiModInstNr[2]) || (10146 == GlobalFiModInstNr[3]))));
	Tile mesh_24_8(
		.clock(clock),
		.io_in_a_0(r_776_0),
		.io_in_b_0(b_280_0),
		.io_in_d_0(b_1304_0),
		.io_in_control_0_dataflow(mesh_24_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2328_0),
		.io_in_last_0(r_3352_0),
		.io_in_valid_0(r_1304_0),
		.io_out_a_0(_mesh_24_8_io_out_a_0),
		.io_out_c_0(_mesh_24_8_io_out_c_0),
		.io_out_b_0(_mesh_24_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_8_io_out_id_0),
		.io_out_last_0(_mesh_24_8_io_out_last_0),
		.io_out_valid_0(_mesh_24_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10147 == GlobalFiModInstNr[0]) || (10147 == GlobalFiModInstNr[1]) || (10147 == GlobalFiModInstNr[2]) || (10147 == GlobalFiModInstNr[3]))));
	Tile mesh_24_9(
		.clock(clock),
		.io_in_a_0(r_777_0),
		.io_in_b_0(b_312_0),
		.io_in_d_0(b_1336_0),
		.io_in_control_0_dataflow(mesh_24_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2360_0),
		.io_in_last_0(r_3384_0),
		.io_in_valid_0(r_1336_0),
		.io_out_a_0(_mesh_24_9_io_out_a_0),
		.io_out_c_0(_mesh_24_9_io_out_c_0),
		.io_out_b_0(_mesh_24_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_9_io_out_id_0),
		.io_out_last_0(_mesh_24_9_io_out_last_0),
		.io_out_valid_0(_mesh_24_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10148 == GlobalFiModInstNr[0]) || (10148 == GlobalFiModInstNr[1]) || (10148 == GlobalFiModInstNr[2]) || (10148 == GlobalFiModInstNr[3]))));
	Tile mesh_24_10(
		.clock(clock),
		.io_in_a_0(r_778_0),
		.io_in_b_0(b_344_0),
		.io_in_d_0(b_1368_0),
		.io_in_control_0_dataflow(mesh_24_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2392_0),
		.io_in_last_0(r_3416_0),
		.io_in_valid_0(r_1368_0),
		.io_out_a_0(_mesh_24_10_io_out_a_0),
		.io_out_c_0(_mesh_24_10_io_out_c_0),
		.io_out_b_0(_mesh_24_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_10_io_out_id_0),
		.io_out_last_0(_mesh_24_10_io_out_last_0),
		.io_out_valid_0(_mesh_24_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10149 == GlobalFiModInstNr[0]) || (10149 == GlobalFiModInstNr[1]) || (10149 == GlobalFiModInstNr[2]) || (10149 == GlobalFiModInstNr[3]))));
	Tile mesh_24_11(
		.clock(clock),
		.io_in_a_0(r_779_0),
		.io_in_b_0(b_376_0),
		.io_in_d_0(b_1400_0),
		.io_in_control_0_dataflow(mesh_24_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2424_0),
		.io_in_last_0(r_3448_0),
		.io_in_valid_0(r_1400_0),
		.io_out_a_0(_mesh_24_11_io_out_a_0),
		.io_out_c_0(_mesh_24_11_io_out_c_0),
		.io_out_b_0(_mesh_24_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_11_io_out_id_0),
		.io_out_last_0(_mesh_24_11_io_out_last_0),
		.io_out_valid_0(_mesh_24_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10150 == GlobalFiModInstNr[0]) || (10150 == GlobalFiModInstNr[1]) || (10150 == GlobalFiModInstNr[2]) || (10150 == GlobalFiModInstNr[3]))));
	Tile mesh_24_12(
		.clock(clock),
		.io_in_a_0(r_780_0),
		.io_in_b_0(b_408_0),
		.io_in_d_0(b_1432_0),
		.io_in_control_0_dataflow(mesh_24_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2456_0),
		.io_in_last_0(r_3480_0),
		.io_in_valid_0(r_1432_0),
		.io_out_a_0(_mesh_24_12_io_out_a_0),
		.io_out_c_0(_mesh_24_12_io_out_c_0),
		.io_out_b_0(_mesh_24_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_12_io_out_id_0),
		.io_out_last_0(_mesh_24_12_io_out_last_0),
		.io_out_valid_0(_mesh_24_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10151 == GlobalFiModInstNr[0]) || (10151 == GlobalFiModInstNr[1]) || (10151 == GlobalFiModInstNr[2]) || (10151 == GlobalFiModInstNr[3]))));
	Tile mesh_24_13(
		.clock(clock),
		.io_in_a_0(r_781_0),
		.io_in_b_0(b_440_0),
		.io_in_d_0(b_1464_0),
		.io_in_control_0_dataflow(mesh_24_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2488_0),
		.io_in_last_0(r_3512_0),
		.io_in_valid_0(r_1464_0),
		.io_out_a_0(_mesh_24_13_io_out_a_0),
		.io_out_c_0(_mesh_24_13_io_out_c_0),
		.io_out_b_0(_mesh_24_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_13_io_out_id_0),
		.io_out_last_0(_mesh_24_13_io_out_last_0),
		.io_out_valid_0(_mesh_24_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10152 == GlobalFiModInstNr[0]) || (10152 == GlobalFiModInstNr[1]) || (10152 == GlobalFiModInstNr[2]) || (10152 == GlobalFiModInstNr[3]))));
	Tile mesh_24_14(
		.clock(clock),
		.io_in_a_0(r_782_0),
		.io_in_b_0(b_472_0),
		.io_in_d_0(b_1496_0),
		.io_in_control_0_dataflow(mesh_24_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2520_0),
		.io_in_last_0(r_3544_0),
		.io_in_valid_0(r_1496_0),
		.io_out_a_0(_mesh_24_14_io_out_a_0),
		.io_out_c_0(_mesh_24_14_io_out_c_0),
		.io_out_b_0(_mesh_24_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_14_io_out_id_0),
		.io_out_last_0(_mesh_24_14_io_out_last_0),
		.io_out_valid_0(_mesh_24_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10153 == GlobalFiModInstNr[0]) || (10153 == GlobalFiModInstNr[1]) || (10153 == GlobalFiModInstNr[2]) || (10153 == GlobalFiModInstNr[3]))));
	Tile mesh_24_15(
		.clock(clock),
		.io_in_a_0(r_783_0),
		.io_in_b_0(b_504_0),
		.io_in_d_0(b_1528_0),
		.io_in_control_0_dataflow(mesh_24_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2552_0),
		.io_in_last_0(r_3576_0),
		.io_in_valid_0(r_1528_0),
		.io_out_a_0(_mesh_24_15_io_out_a_0),
		.io_out_c_0(_mesh_24_15_io_out_c_0),
		.io_out_b_0(_mesh_24_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_15_io_out_id_0),
		.io_out_last_0(_mesh_24_15_io_out_last_0),
		.io_out_valid_0(_mesh_24_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10154 == GlobalFiModInstNr[0]) || (10154 == GlobalFiModInstNr[1]) || (10154 == GlobalFiModInstNr[2]) || (10154 == GlobalFiModInstNr[3]))));
	Tile mesh_24_16(
		.clock(clock),
		.io_in_a_0(r_784_0),
		.io_in_b_0(b_536_0),
		.io_in_d_0(b_1560_0),
		.io_in_control_0_dataflow(mesh_24_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2584_0),
		.io_in_last_0(r_3608_0),
		.io_in_valid_0(r_1560_0),
		.io_out_a_0(_mesh_24_16_io_out_a_0),
		.io_out_c_0(_mesh_24_16_io_out_c_0),
		.io_out_b_0(_mesh_24_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_16_io_out_id_0),
		.io_out_last_0(_mesh_24_16_io_out_last_0),
		.io_out_valid_0(_mesh_24_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10155 == GlobalFiModInstNr[0]) || (10155 == GlobalFiModInstNr[1]) || (10155 == GlobalFiModInstNr[2]) || (10155 == GlobalFiModInstNr[3]))));
	Tile mesh_24_17(
		.clock(clock),
		.io_in_a_0(r_785_0),
		.io_in_b_0(b_568_0),
		.io_in_d_0(b_1592_0),
		.io_in_control_0_dataflow(mesh_24_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2616_0),
		.io_in_last_0(r_3640_0),
		.io_in_valid_0(r_1592_0),
		.io_out_a_0(_mesh_24_17_io_out_a_0),
		.io_out_c_0(_mesh_24_17_io_out_c_0),
		.io_out_b_0(_mesh_24_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_17_io_out_id_0),
		.io_out_last_0(_mesh_24_17_io_out_last_0),
		.io_out_valid_0(_mesh_24_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10156 == GlobalFiModInstNr[0]) || (10156 == GlobalFiModInstNr[1]) || (10156 == GlobalFiModInstNr[2]) || (10156 == GlobalFiModInstNr[3]))));
	Tile mesh_24_18(
		.clock(clock),
		.io_in_a_0(r_786_0),
		.io_in_b_0(b_600_0),
		.io_in_d_0(b_1624_0),
		.io_in_control_0_dataflow(mesh_24_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2648_0),
		.io_in_last_0(r_3672_0),
		.io_in_valid_0(r_1624_0),
		.io_out_a_0(_mesh_24_18_io_out_a_0),
		.io_out_c_0(_mesh_24_18_io_out_c_0),
		.io_out_b_0(_mesh_24_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_18_io_out_id_0),
		.io_out_last_0(_mesh_24_18_io_out_last_0),
		.io_out_valid_0(_mesh_24_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10157 == GlobalFiModInstNr[0]) || (10157 == GlobalFiModInstNr[1]) || (10157 == GlobalFiModInstNr[2]) || (10157 == GlobalFiModInstNr[3]))));
	Tile mesh_24_19(
		.clock(clock),
		.io_in_a_0(r_787_0),
		.io_in_b_0(b_632_0),
		.io_in_d_0(b_1656_0),
		.io_in_control_0_dataflow(mesh_24_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2680_0),
		.io_in_last_0(r_3704_0),
		.io_in_valid_0(r_1656_0),
		.io_out_a_0(_mesh_24_19_io_out_a_0),
		.io_out_c_0(_mesh_24_19_io_out_c_0),
		.io_out_b_0(_mesh_24_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_19_io_out_id_0),
		.io_out_last_0(_mesh_24_19_io_out_last_0),
		.io_out_valid_0(_mesh_24_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10158 == GlobalFiModInstNr[0]) || (10158 == GlobalFiModInstNr[1]) || (10158 == GlobalFiModInstNr[2]) || (10158 == GlobalFiModInstNr[3]))));
	Tile mesh_24_20(
		.clock(clock),
		.io_in_a_0(r_788_0),
		.io_in_b_0(b_664_0),
		.io_in_d_0(b_1688_0),
		.io_in_control_0_dataflow(mesh_24_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2712_0),
		.io_in_last_0(r_3736_0),
		.io_in_valid_0(r_1688_0),
		.io_out_a_0(_mesh_24_20_io_out_a_0),
		.io_out_c_0(_mesh_24_20_io_out_c_0),
		.io_out_b_0(_mesh_24_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_20_io_out_id_0),
		.io_out_last_0(_mesh_24_20_io_out_last_0),
		.io_out_valid_0(_mesh_24_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10159 == GlobalFiModInstNr[0]) || (10159 == GlobalFiModInstNr[1]) || (10159 == GlobalFiModInstNr[2]) || (10159 == GlobalFiModInstNr[3]))));
	Tile mesh_24_21(
		.clock(clock),
		.io_in_a_0(r_789_0),
		.io_in_b_0(b_696_0),
		.io_in_d_0(b_1720_0),
		.io_in_control_0_dataflow(mesh_24_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2744_0),
		.io_in_last_0(r_3768_0),
		.io_in_valid_0(r_1720_0),
		.io_out_a_0(_mesh_24_21_io_out_a_0),
		.io_out_c_0(_mesh_24_21_io_out_c_0),
		.io_out_b_0(_mesh_24_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_21_io_out_id_0),
		.io_out_last_0(_mesh_24_21_io_out_last_0),
		.io_out_valid_0(_mesh_24_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10160 == GlobalFiModInstNr[0]) || (10160 == GlobalFiModInstNr[1]) || (10160 == GlobalFiModInstNr[2]) || (10160 == GlobalFiModInstNr[3]))));
	Tile mesh_24_22(
		.clock(clock),
		.io_in_a_0(r_790_0),
		.io_in_b_0(b_728_0),
		.io_in_d_0(b_1752_0),
		.io_in_control_0_dataflow(mesh_24_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2776_0),
		.io_in_last_0(r_3800_0),
		.io_in_valid_0(r_1752_0),
		.io_out_a_0(_mesh_24_22_io_out_a_0),
		.io_out_c_0(_mesh_24_22_io_out_c_0),
		.io_out_b_0(_mesh_24_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_22_io_out_id_0),
		.io_out_last_0(_mesh_24_22_io_out_last_0),
		.io_out_valid_0(_mesh_24_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10161 == GlobalFiModInstNr[0]) || (10161 == GlobalFiModInstNr[1]) || (10161 == GlobalFiModInstNr[2]) || (10161 == GlobalFiModInstNr[3]))));
	Tile mesh_24_23(
		.clock(clock),
		.io_in_a_0(r_791_0),
		.io_in_b_0(b_760_0),
		.io_in_d_0(b_1784_0),
		.io_in_control_0_dataflow(mesh_24_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2808_0),
		.io_in_last_0(r_3832_0),
		.io_in_valid_0(r_1784_0),
		.io_out_a_0(_mesh_24_23_io_out_a_0),
		.io_out_c_0(_mesh_24_23_io_out_c_0),
		.io_out_b_0(_mesh_24_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_23_io_out_id_0),
		.io_out_last_0(_mesh_24_23_io_out_last_0),
		.io_out_valid_0(_mesh_24_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10162 == GlobalFiModInstNr[0]) || (10162 == GlobalFiModInstNr[1]) || (10162 == GlobalFiModInstNr[2]) || (10162 == GlobalFiModInstNr[3]))));
	Tile mesh_24_24(
		.clock(clock),
		.io_in_a_0(r_792_0),
		.io_in_b_0(b_792_0),
		.io_in_d_0(b_1816_0),
		.io_in_control_0_dataflow(mesh_24_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2840_0),
		.io_in_last_0(r_3864_0),
		.io_in_valid_0(r_1816_0),
		.io_out_a_0(_mesh_24_24_io_out_a_0),
		.io_out_c_0(_mesh_24_24_io_out_c_0),
		.io_out_b_0(_mesh_24_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_24_io_out_id_0),
		.io_out_last_0(_mesh_24_24_io_out_last_0),
		.io_out_valid_0(_mesh_24_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10163 == GlobalFiModInstNr[0]) || (10163 == GlobalFiModInstNr[1]) || (10163 == GlobalFiModInstNr[2]) || (10163 == GlobalFiModInstNr[3]))));
	Tile mesh_24_25(
		.clock(clock),
		.io_in_a_0(r_793_0),
		.io_in_b_0(b_824_0),
		.io_in_d_0(b_1848_0),
		.io_in_control_0_dataflow(mesh_24_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2872_0),
		.io_in_last_0(r_3896_0),
		.io_in_valid_0(r_1848_0),
		.io_out_a_0(_mesh_24_25_io_out_a_0),
		.io_out_c_0(_mesh_24_25_io_out_c_0),
		.io_out_b_0(_mesh_24_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_25_io_out_id_0),
		.io_out_last_0(_mesh_24_25_io_out_last_0),
		.io_out_valid_0(_mesh_24_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10164 == GlobalFiModInstNr[0]) || (10164 == GlobalFiModInstNr[1]) || (10164 == GlobalFiModInstNr[2]) || (10164 == GlobalFiModInstNr[3]))));
	Tile mesh_24_26(
		.clock(clock),
		.io_in_a_0(r_794_0),
		.io_in_b_0(b_856_0),
		.io_in_d_0(b_1880_0),
		.io_in_control_0_dataflow(mesh_24_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2904_0),
		.io_in_last_0(r_3928_0),
		.io_in_valid_0(r_1880_0),
		.io_out_a_0(_mesh_24_26_io_out_a_0),
		.io_out_c_0(_mesh_24_26_io_out_c_0),
		.io_out_b_0(_mesh_24_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_26_io_out_id_0),
		.io_out_last_0(_mesh_24_26_io_out_last_0),
		.io_out_valid_0(_mesh_24_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10165 == GlobalFiModInstNr[0]) || (10165 == GlobalFiModInstNr[1]) || (10165 == GlobalFiModInstNr[2]) || (10165 == GlobalFiModInstNr[3]))));
	Tile mesh_24_27(
		.clock(clock),
		.io_in_a_0(r_795_0),
		.io_in_b_0(b_888_0),
		.io_in_d_0(b_1912_0),
		.io_in_control_0_dataflow(mesh_24_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2936_0),
		.io_in_last_0(r_3960_0),
		.io_in_valid_0(r_1912_0),
		.io_out_a_0(_mesh_24_27_io_out_a_0),
		.io_out_c_0(_mesh_24_27_io_out_c_0),
		.io_out_b_0(_mesh_24_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_27_io_out_id_0),
		.io_out_last_0(_mesh_24_27_io_out_last_0),
		.io_out_valid_0(_mesh_24_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10166 == GlobalFiModInstNr[0]) || (10166 == GlobalFiModInstNr[1]) || (10166 == GlobalFiModInstNr[2]) || (10166 == GlobalFiModInstNr[3]))));
	Tile mesh_24_28(
		.clock(clock),
		.io_in_a_0(r_796_0),
		.io_in_b_0(b_920_0),
		.io_in_d_0(b_1944_0),
		.io_in_control_0_dataflow(mesh_24_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2968_0),
		.io_in_last_0(r_3992_0),
		.io_in_valid_0(r_1944_0),
		.io_out_a_0(_mesh_24_28_io_out_a_0),
		.io_out_c_0(_mesh_24_28_io_out_c_0),
		.io_out_b_0(_mesh_24_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_28_io_out_id_0),
		.io_out_last_0(_mesh_24_28_io_out_last_0),
		.io_out_valid_0(_mesh_24_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10167 == GlobalFiModInstNr[0]) || (10167 == GlobalFiModInstNr[1]) || (10167 == GlobalFiModInstNr[2]) || (10167 == GlobalFiModInstNr[3]))));
	Tile mesh_24_29(
		.clock(clock),
		.io_in_a_0(r_797_0),
		.io_in_b_0(b_952_0),
		.io_in_d_0(b_1976_0),
		.io_in_control_0_dataflow(mesh_24_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3000_0),
		.io_in_last_0(r_4024_0),
		.io_in_valid_0(r_1976_0),
		.io_out_a_0(_mesh_24_29_io_out_a_0),
		.io_out_c_0(_mesh_24_29_io_out_c_0),
		.io_out_b_0(_mesh_24_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_29_io_out_id_0),
		.io_out_last_0(_mesh_24_29_io_out_last_0),
		.io_out_valid_0(_mesh_24_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10168 == GlobalFiModInstNr[0]) || (10168 == GlobalFiModInstNr[1]) || (10168 == GlobalFiModInstNr[2]) || (10168 == GlobalFiModInstNr[3]))));
	Tile mesh_24_30(
		.clock(clock),
		.io_in_a_0(r_798_0),
		.io_in_b_0(b_984_0),
		.io_in_d_0(b_2008_0),
		.io_in_control_0_dataflow(mesh_24_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3032_0),
		.io_in_last_0(r_4056_0),
		.io_in_valid_0(r_2008_0),
		.io_out_a_0(_mesh_24_30_io_out_a_0),
		.io_out_c_0(_mesh_24_30_io_out_c_0),
		.io_out_b_0(_mesh_24_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_30_io_out_id_0),
		.io_out_last_0(_mesh_24_30_io_out_last_0),
		.io_out_valid_0(_mesh_24_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10169 == GlobalFiModInstNr[0]) || (10169 == GlobalFiModInstNr[1]) || (10169 == GlobalFiModInstNr[2]) || (10169 == GlobalFiModInstNr[3]))));
	Tile mesh_24_31(
		.clock(clock),
		.io_in_a_0(r_799_0),
		.io_in_b_0(b_1016_0),
		.io_in_d_0(b_2040_0),
		.io_in_control_0_dataflow(mesh_24_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_24_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_24_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3064_0),
		.io_in_last_0(r_4088_0),
		.io_in_valid_0(r_2040_0),
		.io_out_a_0(_mesh_24_31_io_out_a_0),
		.io_out_c_0(_mesh_24_31_io_out_c_0),
		.io_out_b_0(_mesh_24_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_24_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_24_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_24_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_24_31_io_out_id_0),
		.io_out_last_0(_mesh_24_31_io_out_last_0),
		.io_out_valid_0(_mesh_24_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10170 == GlobalFiModInstNr[0]) || (10170 == GlobalFiModInstNr[1]) || (10170 == GlobalFiModInstNr[2]) || (10170 == GlobalFiModInstNr[3]))));
	Tile mesh_25_0(
		.clock(clock),
		.io_in_a_0(r_800_0),
		.io_in_b_0(b_25_0),
		.io_in_d_0(b_1049_0),
		.io_in_control_0_dataflow(mesh_25_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2073_0),
		.io_in_last_0(r_3097_0),
		.io_in_valid_0(r_1049_0),
		.io_out_a_0(_mesh_25_0_io_out_a_0),
		.io_out_c_0(_mesh_25_0_io_out_c_0),
		.io_out_b_0(_mesh_25_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_0_io_out_id_0),
		.io_out_last_0(_mesh_25_0_io_out_last_0),
		.io_out_valid_0(_mesh_25_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10171 == GlobalFiModInstNr[0]) || (10171 == GlobalFiModInstNr[1]) || (10171 == GlobalFiModInstNr[2]) || (10171 == GlobalFiModInstNr[3]))));
	Tile mesh_25_1(
		.clock(clock),
		.io_in_a_0(r_801_0),
		.io_in_b_0(b_57_0),
		.io_in_d_0(b_1081_0),
		.io_in_control_0_dataflow(mesh_25_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2105_0),
		.io_in_last_0(r_3129_0),
		.io_in_valid_0(r_1081_0),
		.io_out_a_0(_mesh_25_1_io_out_a_0),
		.io_out_c_0(_mesh_25_1_io_out_c_0),
		.io_out_b_0(_mesh_25_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_1_io_out_id_0),
		.io_out_last_0(_mesh_25_1_io_out_last_0),
		.io_out_valid_0(_mesh_25_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10172 == GlobalFiModInstNr[0]) || (10172 == GlobalFiModInstNr[1]) || (10172 == GlobalFiModInstNr[2]) || (10172 == GlobalFiModInstNr[3]))));
	Tile mesh_25_2(
		.clock(clock),
		.io_in_a_0(r_802_0),
		.io_in_b_0(b_89_0),
		.io_in_d_0(b_1113_0),
		.io_in_control_0_dataflow(mesh_25_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2137_0),
		.io_in_last_0(r_3161_0),
		.io_in_valid_0(r_1113_0),
		.io_out_a_0(_mesh_25_2_io_out_a_0),
		.io_out_c_0(_mesh_25_2_io_out_c_0),
		.io_out_b_0(_mesh_25_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_2_io_out_id_0),
		.io_out_last_0(_mesh_25_2_io_out_last_0),
		.io_out_valid_0(_mesh_25_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10173 == GlobalFiModInstNr[0]) || (10173 == GlobalFiModInstNr[1]) || (10173 == GlobalFiModInstNr[2]) || (10173 == GlobalFiModInstNr[3]))));
	Tile mesh_25_3(
		.clock(clock),
		.io_in_a_0(r_803_0),
		.io_in_b_0(b_121_0),
		.io_in_d_0(b_1145_0),
		.io_in_control_0_dataflow(mesh_25_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2169_0),
		.io_in_last_0(r_3193_0),
		.io_in_valid_0(r_1145_0),
		.io_out_a_0(_mesh_25_3_io_out_a_0),
		.io_out_c_0(_mesh_25_3_io_out_c_0),
		.io_out_b_0(_mesh_25_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_3_io_out_id_0),
		.io_out_last_0(_mesh_25_3_io_out_last_0),
		.io_out_valid_0(_mesh_25_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10174 == GlobalFiModInstNr[0]) || (10174 == GlobalFiModInstNr[1]) || (10174 == GlobalFiModInstNr[2]) || (10174 == GlobalFiModInstNr[3]))));
	Tile mesh_25_4(
		.clock(clock),
		.io_in_a_0(r_804_0),
		.io_in_b_0(b_153_0),
		.io_in_d_0(b_1177_0),
		.io_in_control_0_dataflow(mesh_25_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2201_0),
		.io_in_last_0(r_3225_0),
		.io_in_valid_0(r_1177_0),
		.io_out_a_0(_mesh_25_4_io_out_a_0),
		.io_out_c_0(_mesh_25_4_io_out_c_0),
		.io_out_b_0(_mesh_25_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_4_io_out_id_0),
		.io_out_last_0(_mesh_25_4_io_out_last_0),
		.io_out_valid_0(_mesh_25_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10175 == GlobalFiModInstNr[0]) || (10175 == GlobalFiModInstNr[1]) || (10175 == GlobalFiModInstNr[2]) || (10175 == GlobalFiModInstNr[3]))));
	Tile mesh_25_5(
		.clock(clock),
		.io_in_a_0(r_805_0),
		.io_in_b_0(b_185_0),
		.io_in_d_0(b_1209_0),
		.io_in_control_0_dataflow(mesh_25_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2233_0),
		.io_in_last_0(r_3257_0),
		.io_in_valid_0(r_1209_0),
		.io_out_a_0(_mesh_25_5_io_out_a_0),
		.io_out_c_0(_mesh_25_5_io_out_c_0),
		.io_out_b_0(_mesh_25_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_5_io_out_id_0),
		.io_out_last_0(_mesh_25_5_io_out_last_0),
		.io_out_valid_0(_mesh_25_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10176 == GlobalFiModInstNr[0]) || (10176 == GlobalFiModInstNr[1]) || (10176 == GlobalFiModInstNr[2]) || (10176 == GlobalFiModInstNr[3]))));
	Tile mesh_25_6(
		.clock(clock),
		.io_in_a_0(r_806_0),
		.io_in_b_0(b_217_0),
		.io_in_d_0(b_1241_0),
		.io_in_control_0_dataflow(mesh_25_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2265_0),
		.io_in_last_0(r_3289_0),
		.io_in_valid_0(r_1241_0),
		.io_out_a_0(_mesh_25_6_io_out_a_0),
		.io_out_c_0(_mesh_25_6_io_out_c_0),
		.io_out_b_0(_mesh_25_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_6_io_out_id_0),
		.io_out_last_0(_mesh_25_6_io_out_last_0),
		.io_out_valid_0(_mesh_25_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10177 == GlobalFiModInstNr[0]) || (10177 == GlobalFiModInstNr[1]) || (10177 == GlobalFiModInstNr[2]) || (10177 == GlobalFiModInstNr[3]))));
	Tile mesh_25_7(
		.clock(clock),
		.io_in_a_0(r_807_0),
		.io_in_b_0(b_249_0),
		.io_in_d_0(b_1273_0),
		.io_in_control_0_dataflow(mesh_25_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2297_0),
		.io_in_last_0(r_3321_0),
		.io_in_valid_0(r_1273_0),
		.io_out_a_0(_mesh_25_7_io_out_a_0),
		.io_out_c_0(_mesh_25_7_io_out_c_0),
		.io_out_b_0(_mesh_25_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_7_io_out_id_0),
		.io_out_last_0(_mesh_25_7_io_out_last_0),
		.io_out_valid_0(_mesh_25_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10178 == GlobalFiModInstNr[0]) || (10178 == GlobalFiModInstNr[1]) || (10178 == GlobalFiModInstNr[2]) || (10178 == GlobalFiModInstNr[3]))));
	Tile mesh_25_8(
		.clock(clock),
		.io_in_a_0(r_808_0),
		.io_in_b_0(b_281_0),
		.io_in_d_0(b_1305_0),
		.io_in_control_0_dataflow(mesh_25_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2329_0),
		.io_in_last_0(r_3353_0),
		.io_in_valid_0(r_1305_0),
		.io_out_a_0(_mesh_25_8_io_out_a_0),
		.io_out_c_0(_mesh_25_8_io_out_c_0),
		.io_out_b_0(_mesh_25_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_8_io_out_id_0),
		.io_out_last_0(_mesh_25_8_io_out_last_0),
		.io_out_valid_0(_mesh_25_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10179 == GlobalFiModInstNr[0]) || (10179 == GlobalFiModInstNr[1]) || (10179 == GlobalFiModInstNr[2]) || (10179 == GlobalFiModInstNr[3]))));
	Tile mesh_25_9(
		.clock(clock),
		.io_in_a_0(r_809_0),
		.io_in_b_0(b_313_0),
		.io_in_d_0(b_1337_0),
		.io_in_control_0_dataflow(mesh_25_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2361_0),
		.io_in_last_0(r_3385_0),
		.io_in_valid_0(r_1337_0),
		.io_out_a_0(_mesh_25_9_io_out_a_0),
		.io_out_c_0(_mesh_25_9_io_out_c_0),
		.io_out_b_0(_mesh_25_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_9_io_out_id_0),
		.io_out_last_0(_mesh_25_9_io_out_last_0),
		.io_out_valid_0(_mesh_25_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10180 == GlobalFiModInstNr[0]) || (10180 == GlobalFiModInstNr[1]) || (10180 == GlobalFiModInstNr[2]) || (10180 == GlobalFiModInstNr[3]))));
	Tile mesh_25_10(
		.clock(clock),
		.io_in_a_0(r_810_0),
		.io_in_b_0(b_345_0),
		.io_in_d_0(b_1369_0),
		.io_in_control_0_dataflow(mesh_25_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2393_0),
		.io_in_last_0(r_3417_0),
		.io_in_valid_0(r_1369_0),
		.io_out_a_0(_mesh_25_10_io_out_a_0),
		.io_out_c_0(_mesh_25_10_io_out_c_0),
		.io_out_b_0(_mesh_25_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_10_io_out_id_0),
		.io_out_last_0(_mesh_25_10_io_out_last_0),
		.io_out_valid_0(_mesh_25_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10181 == GlobalFiModInstNr[0]) || (10181 == GlobalFiModInstNr[1]) || (10181 == GlobalFiModInstNr[2]) || (10181 == GlobalFiModInstNr[3]))));
	Tile mesh_25_11(
		.clock(clock),
		.io_in_a_0(r_811_0),
		.io_in_b_0(b_377_0),
		.io_in_d_0(b_1401_0),
		.io_in_control_0_dataflow(mesh_25_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2425_0),
		.io_in_last_0(r_3449_0),
		.io_in_valid_0(r_1401_0),
		.io_out_a_0(_mesh_25_11_io_out_a_0),
		.io_out_c_0(_mesh_25_11_io_out_c_0),
		.io_out_b_0(_mesh_25_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_11_io_out_id_0),
		.io_out_last_0(_mesh_25_11_io_out_last_0),
		.io_out_valid_0(_mesh_25_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10182 == GlobalFiModInstNr[0]) || (10182 == GlobalFiModInstNr[1]) || (10182 == GlobalFiModInstNr[2]) || (10182 == GlobalFiModInstNr[3]))));
	Tile mesh_25_12(
		.clock(clock),
		.io_in_a_0(r_812_0),
		.io_in_b_0(b_409_0),
		.io_in_d_0(b_1433_0),
		.io_in_control_0_dataflow(mesh_25_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2457_0),
		.io_in_last_0(r_3481_0),
		.io_in_valid_0(r_1433_0),
		.io_out_a_0(_mesh_25_12_io_out_a_0),
		.io_out_c_0(_mesh_25_12_io_out_c_0),
		.io_out_b_0(_mesh_25_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_12_io_out_id_0),
		.io_out_last_0(_mesh_25_12_io_out_last_0),
		.io_out_valid_0(_mesh_25_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10183 == GlobalFiModInstNr[0]) || (10183 == GlobalFiModInstNr[1]) || (10183 == GlobalFiModInstNr[2]) || (10183 == GlobalFiModInstNr[3]))));
	Tile mesh_25_13(
		.clock(clock),
		.io_in_a_0(r_813_0),
		.io_in_b_0(b_441_0),
		.io_in_d_0(b_1465_0),
		.io_in_control_0_dataflow(mesh_25_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2489_0),
		.io_in_last_0(r_3513_0),
		.io_in_valid_0(r_1465_0),
		.io_out_a_0(_mesh_25_13_io_out_a_0),
		.io_out_c_0(_mesh_25_13_io_out_c_0),
		.io_out_b_0(_mesh_25_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_13_io_out_id_0),
		.io_out_last_0(_mesh_25_13_io_out_last_0),
		.io_out_valid_0(_mesh_25_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10184 == GlobalFiModInstNr[0]) || (10184 == GlobalFiModInstNr[1]) || (10184 == GlobalFiModInstNr[2]) || (10184 == GlobalFiModInstNr[3]))));
	Tile mesh_25_14(
		.clock(clock),
		.io_in_a_0(r_814_0),
		.io_in_b_0(b_473_0),
		.io_in_d_0(b_1497_0),
		.io_in_control_0_dataflow(mesh_25_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2521_0),
		.io_in_last_0(r_3545_0),
		.io_in_valid_0(r_1497_0),
		.io_out_a_0(_mesh_25_14_io_out_a_0),
		.io_out_c_0(_mesh_25_14_io_out_c_0),
		.io_out_b_0(_mesh_25_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_14_io_out_id_0),
		.io_out_last_0(_mesh_25_14_io_out_last_0),
		.io_out_valid_0(_mesh_25_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10185 == GlobalFiModInstNr[0]) || (10185 == GlobalFiModInstNr[1]) || (10185 == GlobalFiModInstNr[2]) || (10185 == GlobalFiModInstNr[3]))));
	Tile mesh_25_15(
		.clock(clock),
		.io_in_a_0(r_815_0),
		.io_in_b_0(b_505_0),
		.io_in_d_0(b_1529_0),
		.io_in_control_0_dataflow(mesh_25_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2553_0),
		.io_in_last_0(r_3577_0),
		.io_in_valid_0(r_1529_0),
		.io_out_a_0(_mesh_25_15_io_out_a_0),
		.io_out_c_0(_mesh_25_15_io_out_c_0),
		.io_out_b_0(_mesh_25_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_15_io_out_id_0),
		.io_out_last_0(_mesh_25_15_io_out_last_0),
		.io_out_valid_0(_mesh_25_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10186 == GlobalFiModInstNr[0]) || (10186 == GlobalFiModInstNr[1]) || (10186 == GlobalFiModInstNr[2]) || (10186 == GlobalFiModInstNr[3]))));
	Tile mesh_25_16(
		.clock(clock),
		.io_in_a_0(r_816_0),
		.io_in_b_0(b_537_0),
		.io_in_d_0(b_1561_0),
		.io_in_control_0_dataflow(mesh_25_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2585_0),
		.io_in_last_0(r_3609_0),
		.io_in_valid_0(r_1561_0),
		.io_out_a_0(_mesh_25_16_io_out_a_0),
		.io_out_c_0(_mesh_25_16_io_out_c_0),
		.io_out_b_0(_mesh_25_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_16_io_out_id_0),
		.io_out_last_0(_mesh_25_16_io_out_last_0),
		.io_out_valid_0(_mesh_25_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10187 == GlobalFiModInstNr[0]) || (10187 == GlobalFiModInstNr[1]) || (10187 == GlobalFiModInstNr[2]) || (10187 == GlobalFiModInstNr[3]))));
	Tile mesh_25_17(
		.clock(clock),
		.io_in_a_0(r_817_0),
		.io_in_b_0(b_569_0),
		.io_in_d_0(b_1593_0),
		.io_in_control_0_dataflow(mesh_25_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2617_0),
		.io_in_last_0(r_3641_0),
		.io_in_valid_0(r_1593_0),
		.io_out_a_0(_mesh_25_17_io_out_a_0),
		.io_out_c_0(_mesh_25_17_io_out_c_0),
		.io_out_b_0(_mesh_25_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_17_io_out_id_0),
		.io_out_last_0(_mesh_25_17_io_out_last_0),
		.io_out_valid_0(_mesh_25_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10188 == GlobalFiModInstNr[0]) || (10188 == GlobalFiModInstNr[1]) || (10188 == GlobalFiModInstNr[2]) || (10188 == GlobalFiModInstNr[3]))));
	Tile mesh_25_18(
		.clock(clock),
		.io_in_a_0(r_818_0),
		.io_in_b_0(b_601_0),
		.io_in_d_0(b_1625_0),
		.io_in_control_0_dataflow(mesh_25_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2649_0),
		.io_in_last_0(r_3673_0),
		.io_in_valid_0(r_1625_0),
		.io_out_a_0(_mesh_25_18_io_out_a_0),
		.io_out_c_0(_mesh_25_18_io_out_c_0),
		.io_out_b_0(_mesh_25_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_18_io_out_id_0),
		.io_out_last_0(_mesh_25_18_io_out_last_0),
		.io_out_valid_0(_mesh_25_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10189 == GlobalFiModInstNr[0]) || (10189 == GlobalFiModInstNr[1]) || (10189 == GlobalFiModInstNr[2]) || (10189 == GlobalFiModInstNr[3]))));
	Tile mesh_25_19(
		.clock(clock),
		.io_in_a_0(r_819_0),
		.io_in_b_0(b_633_0),
		.io_in_d_0(b_1657_0),
		.io_in_control_0_dataflow(mesh_25_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2681_0),
		.io_in_last_0(r_3705_0),
		.io_in_valid_0(r_1657_0),
		.io_out_a_0(_mesh_25_19_io_out_a_0),
		.io_out_c_0(_mesh_25_19_io_out_c_0),
		.io_out_b_0(_mesh_25_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_19_io_out_id_0),
		.io_out_last_0(_mesh_25_19_io_out_last_0),
		.io_out_valid_0(_mesh_25_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10190 == GlobalFiModInstNr[0]) || (10190 == GlobalFiModInstNr[1]) || (10190 == GlobalFiModInstNr[2]) || (10190 == GlobalFiModInstNr[3]))));
	Tile mesh_25_20(
		.clock(clock),
		.io_in_a_0(r_820_0),
		.io_in_b_0(b_665_0),
		.io_in_d_0(b_1689_0),
		.io_in_control_0_dataflow(mesh_25_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2713_0),
		.io_in_last_0(r_3737_0),
		.io_in_valid_0(r_1689_0),
		.io_out_a_0(_mesh_25_20_io_out_a_0),
		.io_out_c_0(_mesh_25_20_io_out_c_0),
		.io_out_b_0(_mesh_25_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_20_io_out_id_0),
		.io_out_last_0(_mesh_25_20_io_out_last_0),
		.io_out_valid_0(_mesh_25_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10191 == GlobalFiModInstNr[0]) || (10191 == GlobalFiModInstNr[1]) || (10191 == GlobalFiModInstNr[2]) || (10191 == GlobalFiModInstNr[3]))));
	Tile mesh_25_21(
		.clock(clock),
		.io_in_a_0(r_821_0),
		.io_in_b_0(b_697_0),
		.io_in_d_0(b_1721_0),
		.io_in_control_0_dataflow(mesh_25_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2745_0),
		.io_in_last_0(r_3769_0),
		.io_in_valid_0(r_1721_0),
		.io_out_a_0(_mesh_25_21_io_out_a_0),
		.io_out_c_0(_mesh_25_21_io_out_c_0),
		.io_out_b_0(_mesh_25_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_21_io_out_id_0),
		.io_out_last_0(_mesh_25_21_io_out_last_0),
		.io_out_valid_0(_mesh_25_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10192 == GlobalFiModInstNr[0]) || (10192 == GlobalFiModInstNr[1]) || (10192 == GlobalFiModInstNr[2]) || (10192 == GlobalFiModInstNr[3]))));
	Tile mesh_25_22(
		.clock(clock),
		.io_in_a_0(r_822_0),
		.io_in_b_0(b_729_0),
		.io_in_d_0(b_1753_0),
		.io_in_control_0_dataflow(mesh_25_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2777_0),
		.io_in_last_0(r_3801_0),
		.io_in_valid_0(r_1753_0),
		.io_out_a_0(_mesh_25_22_io_out_a_0),
		.io_out_c_0(_mesh_25_22_io_out_c_0),
		.io_out_b_0(_mesh_25_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_22_io_out_id_0),
		.io_out_last_0(_mesh_25_22_io_out_last_0),
		.io_out_valid_0(_mesh_25_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10193 == GlobalFiModInstNr[0]) || (10193 == GlobalFiModInstNr[1]) || (10193 == GlobalFiModInstNr[2]) || (10193 == GlobalFiModInstNr[3]))));
	Tile mesh_25_23(
		.clock(clock),
		.io_in_a_0(r_823_0),
		.io_in_b_0(b_761_0),
		.io_in_d_0(b_1785_0),
		.io_in_control_0_dataflow(mesh_25_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2809_0),
		.io_in_last_0(r_3833_0),
		.io_in_valid_0(r_1785_0),
		.io_out_a_0(_mesh_25_23_io_out_a_0),
		.io_out_c_0(_mesh_25_23_io_out_c_0),
		.io_out_b_0(_mesh_25_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_23_io_out_id_0),
		.io_out_last_0(_mesh_25_23_io_out_last_0),
		.io_out_valid_0(_mesh_25_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10194 == GlobalFiModInstNr[0]) || (10194 == GlobalFiModInstNr[1]) || (10194 == GlobalFiModInstNr[2]) || (10194 == GlobalFiModInstNr[3]))));
	Tile mesh_25_24(
		.clock(clock),
		.io_in_a_0(r_824_0),
		.io_in_b_0(b_793_0),
		.io_in_d_0(b_1817_0),
		.io_in_control_0_dataflow(mesh_25_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2841_0),
		.io_in_last_0(r_3865_0),
		.io_in_valid_0(r_1817_0),
		.io_out_a_0(_mesh_25_24_io_out_a_0),
		.io_out_c_0(_mesh_25_24_io_out_c_0),
		.io_out_b_0(_mesh_25_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_24_io_out_id_0),
		.io_out_last_0(_mesh_25_24_io_out_last_0),
		.io_out_valid_0(_mesh_25_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10195 == GlobalFiModInstNr[0]) || (10195 == GlobalFiModInstNr[1]) || (10195 == GlobalFiModInstNr[2]) || (10195 == GlobalFiModInstNr[3]))));
	Tile mesh_25_25(
		.clock(clock),
		.io_in_a_0(r_825_0),
		.io_in_b_0(b_825_0),
		.io_in_d_0(b_1849_0),
		.io_in_control_0_dataflow(mesh_25_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2873_0),
		.io_in_last_0(r_3897_0),
		.io_in_valid_0(r_1849_0),
		.io_out_a_0(_mesh_25_25_io_out_a_0),
		.io_out_c_0(_mesh_25_25_io_out_c_0),
		.io_out_b_0(_mesh_25_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_25_io_out_id_0),
		.io_out_last_0(_mesh_25_25_io_out_last_0),
		.io_out_valid_0(_mesh_25_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10196 == GlobalFiModInstNr[0]) || (10196 == GlobalFiModInstNr[1]) || (10196 == GlobalFiModInstNr[2]) || (10196 == GlobalFiModInstNr[3]))));
	Tile mesh_25_26(
		.clock(clock),
		.io_in_a_0(r_826_0),
		.io_in_b_0(b_857_0),
		.io_in_d_0(b_1881_0),
		.io_in_control_0_dataflow(mesh_25_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2905_0),
		.io_in_last_0(r_3929_0),
		.io_in_valid_0(r_1881_0),
		.io_out_a_0(_mesh_25_26_io_out_a_0),
		.io_out_c_0(_mesh_25_26_io_out_c_0),
		.io_out_b_0(_mesh_25_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_26_io_out_id_0),
		.io_out_last_0(_mesh_25_26_io_out_last_0),
		.io_out_valid_0(_mesh_25_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10197 == GlobalFiModInstNr[0]) || (10197 == GlobalFiModInstNr[1]) || (10197 == GlobalFiModInstNr[2]) || (10197 == GlobalFiModInstNr[3]))));
	Tile mesh_25_27(
		.clock(clock),
		.io_in_a_0(r_827_0),
		.io_in_b_0(b_889_0),
		.io_in_d_0(b_1913_0),
		.io_in_control_0_dataflow(mesh_25_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2937_0),
		.io_in_last_0(r_3961_0),
		.io_in_valid_0(r_1913_0),
		.io_out_a_0(_mesh_25_27_io_out_a_0),
		.io_out_c_0(_mesh_25_27_io_out_c_0),
		.io_out_b_0(_mesh_25_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_27_io_out_id_0),
		.io_out_last_0(_mesh_25_27_io_out_last_0),
		.io_out_valid_0(_mesh_25_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10198 == GlobalFiModInstNr[0]) || (10198 == GlobalFiModInstNr[1]) || (10198 == GlobalFiModInstNr[2]) || (10198 == GlobalFiModInstNr[3]))));
	Tile mesh_25_28(
		.clock(clock),
		.io_in_a_0(r_828_0),
		.io_in_b_0(b_921_0),
		.io_in_d_0(b_1945_0),
		.io_in_control_0_dataflow(mesh_25_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2969_0),
		.io_in_last_0(r_3993_0),
		.io_in_valid_0(r_1945_0),
		.io_out_a_0(_mesh_25_28_io_out_a_0),
		.io_out_c_0(_mesh_25_28_io_out_c_0),
		.io_out_b_0(_mesh_25_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_28_io_out_id_0),
		.io_out_last_0(_mesh_25_28_io_out_last_0),
		.io_out_valid_0(_mesh_25_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10199 == GlobalFiModInstNr[0]) || (10199 == GlobalFiModInstNr[1]) || (10199 == GlobalFiModInstNr[2]) || (10199 == GlobalFiModInstNr[3]))));
	Tile mesh_25_29(
		.clock(clock),
		.io_in_a_0(r_829_0),
		.io_in_b_0(b_953_0),
		.io_in_d_0(b_1977_0),
		.io_in_control_0_dataflow(mesh_25_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3001_0),
		.io_in_last_0(r_4025_0),
		.io_in_valid_0(r_1977_0),
		.io_out_a_0(_mesh_25_29_io_out_a_0),
		.io_out_c_0(_mesh_25_29_io_out_c_0),
		.io_out_b_0(_mesh_25_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_29_io_out_id_0),
		.io_out_last_0(_mesh_25_29_io_out_last_0),
		.io_out_valid_0(_mesh_25_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10200 == GlobalFiModInstNr[0]) || (10200 == GlobalFiModInstNr[1]) || (10200 == GlobalFiModInstNr[2]) || (10200 == GlobalFiModInstNr[3]))));
	Tile mesh_25_30(
		.clock(clock),
		.io_in_a_0(r_830_0),
		.io_in_b_0(b_985_0),
		.io_in_d_0(b_2009_0),
		.io_in_control_0_dataflow(mesh_25_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3033_0),
		.io_in_last_0(r_4057_0),
		.io_in_valid_0(r_2009_0),
		.io_out_a_0(_mesh_25_30_io_out_a_0),
		.io_out_c_0(_mesh_25_30_io_out_c_0),
		.io_out_b_0(_mesh_25_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_30_io_out_id_0),
		.io_out_last_0(_mesh_25_30_io_out_last_0),
		.io_out_valid_0(_mesh_25_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10201 == GlobalFiModInstNr[0]) || (10201 == GlobalFiModInstNr[1]) || (10201 == GlobalFiModInstNr[2]) || (10201 == GlobalFiModInstNr[3]))));
	Tile mesh_25_31(
		.clock(clock),
		.io_in_a_0(r_831_0),
		.io_in_b_0(b_1017_0),
		.io_in_d_0(b_2041_0),
		.io_in_control_0_dataflow(mesh_25_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_25_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_25_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3065_0),
		.io_in_last_0(r_4089_0),
		.io_in_valid_0(r_2041_0),
		.io_out_a_0(_mesh_25_31_io_out_a_0),
		.io_out_c_0(_mesh_25_31_io_out_c_0),
		.io_out_b_0(_mesh_25_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_25_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_25_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_25_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_25_31_io_out_id_0),
		.io_out_last_0(_mesh_25_31_io_out_last_0),
		.io_out_valid_0(_mesh_25_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10202 == GlobalFiModInstNr[0]) || (10202 == GlobalFiModInstNr[1]) || (10202 == GlobalFiModInstNr[2]) || (10202 == GlobalFiModInstNr[3]))));
	Tile mesh_26_0(
		.clock(clock),
		.io_in_a_0(r_832_0),
		.io_in_b_0(b_26_0),
		.io_in_d_0(b_1050_0),
		.io_in_control_0_dataflow(mesh_26_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2074_0),
		.io_in_last_0(r_3098_0),
		.io_in_valid_0(r_1050_0),
		.io_out_a_0(_mesh_26_0_io_out_a_0),
		.io_out_c_0(_mesh_26_0_io_out_c_0),
		.io_out_b_0(_mesh_26_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_0_io_out_id_0),
		.io_out_last_0(_mesh_26_0_io_out_last_0),
		.io_out_valid_0(_mesh_26_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10203 == GlobalFiModInstNr[0]) || (10203 == GlobalFiModInstNr[1]) || (10203 == GlobalFiModInstNr[2]) || (10203 == GlobalFiModInstNr[3]))));
	Tile mesh_26_1(
		.clock(clock),
		.io_in_a_0(r_833_0),
		.io_in_b_0(b_58_0),
		.io_in_d_0(b_1082_0),
		.io_in_control_0_dataflow(mesh_26_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2106_0),
		.io_in_last_0(r_3130_0),
		.io_in_valid_0(r_1082_0),
		.io_out_a_0(_mesh_26_1_io_out_a_0),
		.io_out_c_0(_mesh_26_1_io_out_c_0),
		.io_out_b_0(_mesh_26_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_1_io_out_id_0),
		.io_out_last_0(_mesh_26_1_io_out_last_0),
		.io_out_valid_0(_mesh_26_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10204 == GlobalFiModInstNr[0]) || (10204 == GlobalFiModInstNr[1]) || (10204 == GlobalFiModInstNr[2]) || (10204 == GlobalFiModInstNr[3]))));
	Tile mesh_26_2(
		.clock(clock),
		.io_in_a_0(r_834_0),
		.io_in_b_0(b_90_0),
		.io_in_d_0(b_1114_0),
		.io_in_control_0_dataflow(mesh_26_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2138_0),
		.io_in_last_0(r_3162_0),
		.io_in_valid_0(r_1114_0),
		.io_out_a_0(_mesh_26_2_io_out_a_0),
		.io_out_c_0(_mesh_26_2_io_out_c_0),
		.io_out_b_0(_mesh_26_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_2_io_out_id_0),
		.io_out_last_0(_mesh_26_2_io_out_last_0),
		.io_out_valid_0(_mesh_26_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10205 == GlobalFiModInstNr[0]) || (10205 == GlobalFiModInstNr[1]) || (10205 == GlobalFiModInstNr[2]) || (10205 == GlobalFiModInstNr[3]))));
	Tile mesh_26_3(
		.clock(clock),
		.io_in_a_0(r_835_0),
		.io_in_b_0(b_122_0),
		.io_in_d_0(b_1146_0),
		.io_in_control_0_dataflow(mesh_26_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2170_0),
		.io_in_last_0(r_3194_0),
		.io_in_valid_0(r_1146_0),
		.io_out_a_0(_mesh_26_3_io_out_a_0),
		.io_out_c_0(_mesh_26_3_io_out_c_0),
		.io_out_b_0(_mesh_26_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_3_io_out_id_0),
		.io_out_last_0(_mesh_26_3_io_out_last_0),
		.io_out_valid_0(_mesh_26_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10206 == GlobalFiModInstNr[0]) || (10206 == GlobalFiModInstNr[1]) || (10206 == GlobalFiModInstNr[2]) || (10206 == GlobalFiModInstNr[3]))));
	Tile mesh_26_4(
		.clock(clock),
		.io_in_a_0(r_836_0),
		.io_in_b_0(b_154_0),
		.io_in_d_0(b_1178_0),
		.io_in_control_0_dataflow(mesh_26_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2202_0),
		.io_in_last_0(r_3226_0),
		.io_in_valid_0(r_1178_0),
		.io_out_a_0(_mesh_26_4_io_out_a_0),
		.io_out_c_0(_mesh_26_4_io_out_c_0),
		.io_out_b_0(_mesh_26_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_4_io_out_id_0),
		.io_out_last_0(_mesh_26_4_io_out_last_0),
		.io_out_valid_0(_mesh_26_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10207 == GlobalFiModInstNr[0]) || (10207 == GlobalFiModInstNr[1]) || (10207 == GlobalFiModInstNr[2]) || (10207 == GlobalFiModInstNr[3]))));
	Tile mesh_26_5(
		.clock(clock),
		.io_in_a_0(r_837_0),
		.io_in_b_0(b_186_0),
		.io_in_d_0(b_1210_0),
		.io_in_control_0_dataflow(mesh_26_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2234_0),
		.io_in_last_0(r_3258_0),
		.io_in_valid_0(r_1210_0),
		.io_out_a_0(_mesh_26_5_io_out_a_0),
		.io_out_c_0(_mesh_26_5_io_out_c_0),
		.io_out_b_0(_mesh_26_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_5_io_out_id_0),
		.io_out_last_0(_mesh_26_5_io_out_last_0),
		.io_out_valid_0(_mesh_26_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10208 == GlobalFiModInstNr[0]) || (10208 == GlobalFiModInstNr[1]) || (10208 == GlobalFiModInstNr[2]) || (10208 == GlobalFiModInstNr[3]))));
	Tile mesh_26_6(
		.clock(clock),
		.io_in_a_0(r_838_0),
		.io_in_b_0(b_218_0),
		.io_in_d_0(b_1242_0),
		.io_in_control_0_dataflow(mesh_26_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2266_0),
		.io_in_last_0(r_3290_0),
		.io_in_valid_0(r_1242_0),
		.io_out_a_0(_mesh_26_6_io_out_a_0),
		.io_out_c_0(_mesh_26_6_io_out_c_0),
		.io_out_b_0(_mesh_26_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_6_io_out_id_0),
		.io_out_last_0(_mesh_26_6_io_out_last_0),
		.io_out_valid_0(_mesh_26_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10209 == GlobalFiModInstNr[0]) || (10209 == GlobalFiModInstNr[1]) || (10209 == GlobalFiModInstNr[2]) || (10209 == GlobalFiModInstNr[3]))));
	Tile mesh_26_7(
		.clock(clock),
		.io_in_a_0(r_839_0),
		.io_in_b_0(b_250_0),
		.io_in_d_0(b_1274_0),
		.io_in_control_0_dataflow(mesh_26_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2298_0),
		.io_in_last_0(r_3322_0),
		.io_in_valid_0(r_1274_0),
		.io_out_a_0(_mesh_26_7_io_out_a_0),
		.io_out_c_0(_mesh_26_7_io_out_c_0),
		.io_out_b_0(_mesh_26_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_7_io_out_id_0),
		.io_out_last_0(_mesh_26_7_io_out_last_0),
		.io_out_valid_0(_mesh_26_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10210 == GlobalFiModInstNr[0]) || (10210 == GlobalFiModInstNr[1]) || (10210 == GlobalFiModInstNr[2]) || (10210 == GlobalFiModInstNr[3]))));
	Tile mesh_26_8(
		.clock(clock),
		.io_in_a_0(r_840_0),
		.io_in_b_0(b_282_0),
		.io_in_d_0(b_1306_0),
		.io_in_control_0_dataflow(mesh_26_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2330_0),
		.io_in_last_0(r_3354_0),
		.io_in_valid_0(r_1306_0),
		.io_out_a_0(_mesh_26_8_io_out_a_0),
		.io_out_c_0(_mesh_26_8_io_out_c_0),
		.io_out_b_0(_mesh_26_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_8_io_out_id_0),
		.io_out_last_0(_mesh_26_8_io_out_last_0),
		.io_out_valid_0(_mesh_26_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10211 == GlobalFiModInstNr[0]) || (10211 == GlobalFiModInstNr[1]) || (10211 == GlobalFiModInstNr[2]) || (10211 == GlobalFiModInstNr[3]))));
	Tile mesh_26_9(
		.clock(clock),
		.io_in_a_0(r_841_0),
		.io_in_b_0(b_314_0),
		.io_in_d_0(b_1338_0),
		.io_in_control_0_dataflow(mesh_26_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2362_0),
		.io_in_last_0(r_3386_0),
		.io_in_valid_0(r_1338_0),
		.io_out_a_0(_mesh_26_9_io_out_a_0),
		.io_out_c_0(_mesh_26_9_io_out_c_0),
		.io_out_b_0(_mesh_26_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_9_io_out_id_0),
		.io_out_last_0(_mesh_26_9_io_out_last_0),
		.io_out_valid_0(_mesh_26_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10212 == GlobalFiModInstNr[0]) || (10212 == GlobalFiModInstNr[1]) || (10212 == GlobalFiModInstNr[2]) || (10212 == GlobalFiModInstNr[3]))));
	Tile mesh_26_10(
		.clock(clock),
		.io_in_a_0(r_842_0),
		.io_in_b_0(b_346_0),
		.io_in_d_0(b_1370_0),
		.io_in_control_0_dataflow(mesh_26_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2394_0),
		.io_in_last_0(r_3418_0),
		.io_in_valid_0(r_1370_0),
		.io_out_a_0(_mesh_26_10_io_out_a_0),
		.io_out_c_0(_mesh_26_10_io_out_c_0),
		.io_out_b_0(_mesh_26_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_10_io_out_id_0),
		.io_out_last_0(_mesh_26_10_io_out_last_0),
		.io_out_valid_0(_mesh_26_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10213 == GlobalFiModInstNr[0]) || (10213 == GlobalFiModInstNr[1]) || (10213 == GlobalFiModInstNr[2]) || (10213 == GlobalFiModInstNr[3]))));
	Tile mesh_26_11(
		.clock(clock),
		.io_in_a_0(r_843_0),
		.io_in_b_0(b_378_0),
		.io_in_d_0(b_1402_0),
		.io_in_control_0_dataflow(mesh_26_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2426_0),
		.io_in_last_0(r_3450_0),
		.io_in_valid_0(r_1402_0),
		.io_out_a_0(_mesh_26_11_io_out_a_0),
		.io_out_c_0(_mesh_26_11_io_out_c_0),
		.io_out_b_0(_mesh_26_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_11_io_out_id_0),
		.io_out_last_0(_mesh_26_11_io_out_last_0),
		.io_out_valid_0(_mesh_26_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10214 == GlobalFiModInstNr[0]) || (10214 == GlobalFiModInstNr[1]) || (10214 == GlobalFiModInstNr[2]) || (10214 == GlobalFiModInstNr[3]))));
	Tile mesh_26_12(
		.clock(clock),
		.io_in_a_0(r_844_0),
		.io_in_b_0(b_410_0),
		.io_in_d_0(b_1434_0),
		.io_in_control_0_dataflow(mesh_26_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2458_0),
		.io_in_last_0(r_3482_0),
		.io_in_valid_0(r_1434_0),
		.io_out_a_0(_mesh_26_12_io_out_a_0),
		.io_out_c_0(_mesh_26_12_io_out_c_0),
		.io_out_b_0(_mesh_26_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_12_io_out_id_0),
		.io_out_last_0(_mesh_26_12_io_out_last_0),
		.io_out_valid_0(_mesh_26_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10215 == GlobalFiModInstNr[0]) || (10215 == GlobalFiModInstNr[1]) || (10215 == GlobalFiModInstNr[2]) || (10215 == GlobalFiModInstNr[3]))));
	Tile mesh_26_13(
		.clock(clock),
		.io_in_a_0(r_845_0),
		.io_in_b_0(b_442_0),
		.io_in_d_0(b_1466_0),
		.io_in_control_0_dataflow(mesh_26_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2490_0),
		.io_in_last_0(r_3514_0),
		.io_in_valid_0(r_1466_0),
		.io_out_a_0(_mesh_26_13_io_out_a_0),
		.io_out_c_0(_mesh_26_13_io_out_c_0),
		.io_out_b_0(_mesh_26_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_13_io_out_id_0),
		.io_out_last_0(_mesh_26_13_io_out_last_0),
		.io_out_valid_0(_mesh_26_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10216 == GlobalFiModInstNr[0]) || (10216 == GlobalFiModInstNr[1]) || (10216 == GlobalFiModInstNr[2]) || (10216 == GlobalFiModInstNr[3]))));
	Tile mesh_26_14(
		.clock(clock),
		.io_in_a_0(r_846_0),
		.io_in_b_0(b_474_0),
		.io_in_d_0(b_1498_0),
		.io_in_control_0_dataflow(mesh_26_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2522_0),
		.io_in_last_0(r_3546_0),
		.io_in_valid_0(r_1498_0),
		.io_out_a_0(_mesh_26_14_io_out_a_0),
		.io_out_c_0(_mesh_26_14_io_out_c_0),
		.io_out_b_0(_mesh_26_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_14_io_out_id_0),
		.io_out_last_0(_mesh_26_14_io_out_last_0),
		.io_out_valid_0(_mesh_26_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10217 == GlobalFiModInstNr[0]) || (10217 == GlobalFiModInstNr[1]) || (10217 == GlobalFiModInstNr[2]) || (10217 == GlobalFiModInstNr[3]))));
	Tile mesh_26_15(
		.clock(clock),
		.io_in_a_0(r_847_0),
		.io_in_b_0(b_506_0),
		.io_in_d_0(b_1530_0),
		.io_in_control_0_dataflow(mesh_26_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2554_0),
		.io_in_last_0(r_3578_0),
		.io_in_valid_0(r_1530_0),
		.io_out_a_0(_mesh_26_15_io_out_a_0),
		.io_out_c_0(_mesh_26_15_io_out_c_0),
		.io_out_b_0(_mesh_26_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_15_io_out_id_0),
		.io_out_last_0(_mesh_26_15_io_out_last_0),
		.io_out_valid_0(_mesh_26_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10218 == GlobalFiModInstNr[0]) || (10218 == GlobalFiModInstNr[1]) || (10218 == GlobalFiModInstNr[2]) || (10218 == GlobalFiModInstNr[3]))));
	Tile mesh_26_16(
		.clock(clock),
		.io_in_a_0(r_848_0),
		.io_in_b_0(b_538_0),
		.io_in_d_0(b_1562_0),
		.io_in_control_0_dataflow(mesh_26_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2586_0),
		.io_in_last_0(r_3610_0),
		.io_in_valid_0(r_1562_0),
		.io_out_a_0(_mesh_26_16_io_out_a_0),
		.io_out_c_0(_mesh_26_16_io_out_c_0),
		.io_out_b_0(_mesh_26_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_16_io_out_id_0),
		.io_out_last_0(_mesh_26_16_io_out_last_0),
		.io_out_valid_0(_mesh_26_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10219 == GlobalFiModInstNr[0]) || (10219 == GlobalFiModInstNr[1]) || (10219 == GlobalFiModInstNr[2]) || (10219 == GlobalFiModInstNr[3]))));
	Tile mesh_26_17(
		.clock(clock),
		.io_in_a_0(r_849_0),
		.io_in_b_0(b_570_0),
		.io_in_d_0(b_1594_0),
		.io_in_control_0_dataflow(mesh_26_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2618_0),
		.io_in_last_0(r_3642_0),
		.io_in_valid_0(r_1594_0),
		.io_out_a_0(_mesh_26_17_io_out_a_0),
		.io_out_c_0(_mesh_26_17_io_out_c_0),
		.io_out_b_0(_mesh_26_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_17_io_out_id_0),
		.io_out_last_0(_mesh_26_17_io_out_last_0),
		.io_out_valid_0(_mesh_26_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10220 == GlobalFiModInstNr[0]) || (10220 == GlobalFiModInstNr[1]) || (10220 == GlobalFiModInstNr[2]) || (10220 == GlobalFiModInstNr[3]))));
	Tile mesh_26_18(
		.clock(clock),
		.io_in_a_0(r_850_0),
		.io_in_b_0(b_602_0),
		.io_in_d_0(b_1626_0),
		.io_in_control_0_dataflow(mesh_26_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2650_0),
		.io_in_last_0(r_3674_0),
		.io_in_valid_0(r_1626_0),
		.io_out_a_0(_mesh_26_18_io_out_a_0),
		.io_out_c_0(_mesh_26_18_io_out_c_0),
		.io_out_b_0(_mesh_26_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_18_io_out_id_0),
		.io_out_last_0(_mesh_26_18_io_out_last_0),
		.io_out_valid_0(_mesh_26_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10221 == GlobalFiModInstNr[0]) || (10221 == GlobalFiModInstNr[1]) || (10221 == GlobalFiModInstNr[2]) || (10221 == GlobalFiModInstNr[3]))));
	Tile mesh_26_19(
		.clock(clock),
		.io_in_a_0(r_851_0),
		.io_in_b_0(b_634_0),
		.io_in_d_0(b_1658_0),
		.io_in_control_0_dataflow(mesh_26_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2682_0),
		.io_in_last_0(r_3706_0),
		.io_in_valid_0(r_1658_0),
		.io_out_a_0(_mesh_26_19_io_out_a_0),
		.io_out_c_0(_mesh_26_19_io_out_c_0),
		.io_out_b_0(_mesh_26_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_19_io_out_id_0),
		.io_out_last_0(_mesh_26_19_io_out_last_0),
		.io_out_valid_0(_mesh_26_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10222 == GlobalFiModInstNr[0]) || (10222 == GlobalFiModInstNr[1]) || (10222 == GlobalFiModInstNr[2]) || (10222 == GlobalFiModInstNr[3]))));
	Tile mesh_26_20(
		.clock(clock),
		.io_in_a_0(r_852_0),
		.io_in_b_0(b_666_0),
		.io_in_d_0(b_1690_0),
		.io_in_control_0_dataflow(mesh_26_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2714_0),
		.io_in_last_0(r_3738_0),
		.io_in_valid_0(r_1690_0),
		.io_out_a_0(_mesh_26_20_io_out_a_0),
		.io_out_c_0(_mesh_26_20_io_out_c_0),
		.io_out_b_0(_mesh_26_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_20_io_out_id_0),
		.io_out_last_0(_mesh_26_20_io_out_last_0),
		.io_out_valid_0(_mesh_26_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10223 == GlobalFiModInstNr[0]) || (10223 == GlobalFiModInstNr[1]) || (10223 == GlobalFiModInstNr[2]) || (10223 == GlobalFiModInstNr[3]))));
	Tile mesh_26_21(
		.clock(clock),
		.io_in_a_0(r_853_0),
		.io_in_b_0(b_698_0),
		.io_in_d_0(b_1722_0),
		.io_in_control_0_dataflow(mesh_26_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2746_0),
		.io_in_last_0(r_3770_0),
		.io_in_valid_0(r_1722_0),
		.io_out_a_0(_mesh_26_21_io_out_a_0),
		.io_out_c_0(_mesh_26_21_io_out_c_0),
		.io_out_b_0(_mesh_26_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_21_io_out_id_0),
		.io_out_last_0(_mesh_26_21_io_out_last_0),
		.io_out_valid_0(_mesh_26_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10224 == GlobalFiModInstNr[0]) || (10224 == GlobalFiModInstNr[1]) || (10224 == GlobalFiModInstNr[2]) || (10224 == GlobalFiModInstNr[3]))));
	Tile mesh_26_22(
		.clock(clock),
		.io_in_a_0(r_854_0),
		.io_in_b_0(b_730_0),
		.io_in_d_0(b_1754_0),
		.io_in_control_0_dataflow(mesh_26_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2778_0),
		.io_in_last_0(r_3802_0),
		.io_in_valid_0(r_1754_0),
		.io_out_a_0(_mesh_26_22_io_out_a_0),
		.io_out_c_0(_mesh_26_22_io_out_c_0),
		.io_out_b_0(_mesh_26_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_22_io_out_id_0),
		.io_out_last_0(_mesh_26_22_io_out_last_0),
		.io_out_valid_0(_mesh_26_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10225 == GlobalFiModInstNr[0]) || (10225 == GlobalFiModInstNr[1]) || (10225 == GlobalFiModInstNr[2]) || (10225 == GlobalFiModInstNr[3]))));
	Tile mesh_26_23(
		.clock(clock),
		.io_in_a_0(r_855_0),
		.io_in_b_0(b_762_0),
		.io_in_d_0(b_1786_0),
		.io_in_control_0_dataflow(mesh_26_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2810_0),
		.io_in_last_0(r_3834_0),
		.io_in_valid_0(r_1786_0),
		.io_out_a_0(_mesh_26_23_io_out_a_0),
		.io_out_c_0(_mesh_26_23_io_out_c_0),
		.io_out_b_0(_mesh_26_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_23_io_out_id_0),
		.io_out_last_0(_mesh_26_23_io_out_last_0),
		.io_out_valid_0(_mesh_26_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10226 == GlobalFiModInstNr[0]) || (10226 == GlobalFiModInstNr[1]) || (10226 == GlobalFiModInstNr[2]) || (10226 == GlobalFiModInstNr[3]))));
	Tile mesh_26_24(
		.clock(clock),
		.io_in_a_0(r_856_0),
		.io_in_b_0(b_794_0),
		.io_in_d_0(b_1818_0),
		.io_in_control_0_dataflow(mesh_26_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2842_0),
		.io_in_last_0(r_3866_0),
		.io_in_valid_0(r_1818_0),
		.io_out_a_0(_mesh_26_24_io_out_a_0),
		.io_out_c_0(_mesh_26_24_io_out_c_0),
		.io_out_b_0(_mesh_26_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_24_io_out_id_0),
		.io_out_last_0(_mesh_26_24_io_out_last_0),
		.io_out_valid_0(_mesh_26_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10227 == GlobalFiModInstNr[0]) || (10227 == GlobalFiModInstNr[1]) || (10227 == GlobalFiModInstNr[2]) || (10227 == GlobalFiModInstNr[3]))));
	Tile mesh_26_25(
		.clock(clock),
		.io_in_a_0(r_857_0),
		.io_in_b_0(b_826_0),
		.io_in_d_0(b_1850_0),
		.io_in_control_0_dataflow(mesh_26_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2874_0),
		.io_in_last_0(r_3898_0),
		.io_in_valid_0(r_1850_0),
		.io_out_a_0(_mesh_26_25_io_out_a_0),
		.io_out_c_0(_mesh_26_25_io_out_c_0),
		.io_out_b_0(_mesh_26_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_25_io_out_id_0),
		.io_out_last_0(_mesh_26_25_io_out_last_0),
		.io_out_valid_0(_mesh_26_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10228 == GlobalFiModInstNr[0]) || (10228 == GlobalFiModInstNr[1]) || (10228 == GlobalFiModInstNr[2]) || (10228 == GlobalFiModInstNr[3]))));
	Tile mesh_26_26(
		.clock(clock),
		.io_in_a_0(r_858_0),
		.io_in_b_0(b_858_0),
		.io_in_d_0(b_1882_0),
		.io_in_control_0_dataflow(mesh_26_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2906_0),
		.io_in_last_0(r_3930_0),
		.io_in_valid_0(r_1882_0),
		.io_out_a_0(_mesh_26_26_io_out_a_0),
		.io_out_c_0(_mesh_26_26_io_out_c_0),
		.io_out_b_0(_mesh_26_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_26_io_out_id_0),
		.io_out_last_0(_mesh_26_26_io_out_last_0),
		.io_out_valid_0(_mesh_26_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10229 == GlobalFiModInstNr[0]) || (10229 == GlobalFiModInstNr[1]) || (10229 == GlobalFiModInstNr[2]) || (10229 == GlobalFiModInstNr[3]))));
	Tile mesh_26_27(
		.clock(clock),
		.io_in_a_0(r_859_0),
		.io_in_b_0(b_890_0),
		.io_in_d_0(b_1914_0),
		.io_in_control_0_dataflow(mesh_26_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2938_0),
		.io_in_last_0(r_3962_0),
		.io_in_valid_0(r_1914_0),
		.io_out_a_0(_mesh_26_27_io_out_a_0),
		.io_out_c_0(_mesh_26_27_io_out_c_0),
		.io_out_b_0(_mesh_26_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_27_io_out_id_0),
		.io_out_last_0(_mesh_26_27_io_out_last_0),
		.io_out_valid_0(_mesh_26_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10230 == GlobalFiModInstNr[0]) || (10230 == GlobalFiModInstNr[1]) || (10230 == GlobalFiModInstNr[2]) || (10230 == GlobalFiModInstNr[3]))));
	Tile mesh_26_28(
		.clock(clock),
		.io_in_a_0(r_860_0),
		.io_in_b_0(b_922_0),
		.io_in_d_0(b_1946_0),
		.io_in_control_0_dataflow(mesh_26_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2970_0),
		.io_in_last_0(r_3994_0),
		.io_in_valid_0(r_1946_0),
		.io_out_a_0(_mesh_26_28_io_out_a_0),
		.io_out_c_0(_mesh_26_28_io_out_c_0),
		.io_out_b_0(_mesh_26_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_28_io_out_id_0),
		.io_out_last_0(_mesh_26_28_io_out_last_0),
		.io_out_valid_0(_mesh_26_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10231 == GlobalFiModInstNr[0]) || (10231 == GlobalFiModInstNr[1]) || (10231 == GlobalFiModInstNr[2]) || (10231 == GlobalFiModInstNr[3]))));
	Tile mesh_26_29(
		.clock(clock),
		.io_in_a_0(r_861_0),
		.io_in_b_0(b_954_0),
		.io_in_d_0(b_1978_0),
		.io_in_control_0_dataflow(mesh_26_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3002_0),
		.io_in_last_0(r_4026_0),
		.io_in_valid_0(r_1978_0),
		.io_out_a_0(_mesh_26_29_io_out_a_0),
		.io_out_c_0(_mesh_26_29_io_out_c_0),
		.io_out_b_0(_mesh_26_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_29_io_out_id_0),
		.io_out_last_0(_mesh_26_29_io_out_last_0),
		.io_out_valid_0(_mesh_26_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10232 == GlobalFiModInstNr[0]) || (10232 == GlobalFiModInstNr[1]) || (10232 == GlobalFiModInstNr[2]) || (10232 == GlobalFiModInstNr[3]))));
	Tile mesh_26_30(
		.clock(clock),
		.io_in_a_0(r_862_0),
		.io_in_b_0(b_986_0),
		.io_in_d_0(b_2010_0),
		.io_in_control_0_dataflow(mesh_26_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3034_0),
		.io_in_last_0(r_4058_0),
		.io_in_valid_0(r_2010_0),
		.io_out_a_0(_mesh_26_30_io_out_a_0),
		.io_out_c_0(_mesh_26_30_io_out_c_0),
		.io_out_b_0(_mesh_26_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_30_io_out_id_0),
		.io_out_last_0(_mesh_26_30_io_out_last_0),
		.io_out_valid_0(_mesh_26_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10233 == GlobalFiModInstNr[0]) || (10233 == GlobalFiModInstNr[1]) || (10233 == GlobalFiModInstNr[2]) || (10233 == GlobalFiModInstNr[3]))));
	Tile mesh_26_31(
		.clock(clock),
		.io_in_a_0(r_863_0),
		.io_in_b_0(b_1018_0),
		.io_in_d_0(b_2042_0),
		.io_in_control_0_dataflow(mesh_26_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_26_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_26_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3066_0),
		.io_in_last_0(r_4090_0),
		.io_in_valid_0(r_2042_0),
		.io_out_a_0(_mesh_26_31_io_out_a_0),
		.io_out_c_0(_mesh_26_31_io_out_c_0),
		.io_out_b_0(_mesh_26_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_26_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_26_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_26_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_26_31_io_out_id_0),
		.io_out_last_0(_mesh_26_31_io_out_last_0),
		.io_out_valid_0(_mesh_26_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10234 == GlobalFiModInstNr[0]) || (10234 == GlobalFiModInstNr[1]) || (10234 == GlobalFiModInstNr[2]) || (10234 == GlobalFiModInstNr[3]))));
	Tile mesh_27_0(
		.clock(clock),
		.io_in_a_0(r_864_0),
		.io_in_b_0(b_27_0),
		.io_in_d_0(b_1051_0),
		.io_in_control_0_dataflow(mesh_27_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2075_0),
		.io_in_last_0(r_3099_0),
		.io_in_valid_0(r_1051_0),
		.io_out_a_0(_mesh_27_0_io_out_a_0),
		.io_out_c_0(_mesh_27_0_io_out_c_0),
		.io_out_b_0(_mesh_27_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_0_io_out_id_0),
		.io_out_last_0(_mesh_27_0_io_out_last_0),
		.io_out_valid_0(_mesh_27_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10235 == GlobalFiModInstNr[0]) || (10235 == GlobalFiModInstNr[1]) || (10235 == GlobalFiModInstNr[2]) || (10235 == GlobalFiModInstNr[3]))));
	Tile mesh_27_1(
		.clock(clock),
		.io_in_a_0(r_865_0),
		.io_in_b_0(b_59_0),
		.io_in_d_0(b_1083_0),
		.io_in_control_0_dataflow(mesh_27_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2107_0),
		.io_in_last_0(r_3131_0),
		.io_in_valid_0(r_1083_0),
		.io_out_a_0(_mesh_27_1_io_out_a_0),
		.io_out_c_0(_mesh_27_1_io_out_c_0),
		.io_out_b_0(_mesh_27_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_1_io_out_id_0),
		.io_out_last_0(_mesh_27_1_io_out_last_0),
		.io_out_valid_0(_mesh_27_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10236 == GlobalFiModInstNr[0]) || (10236 == GlobalFiModInstNr[1]) || (10236 == GlobalFiModInstNr[2]) || (10236 == GlobalFiModInstNr[3]))));
	Tile mesh_27_2(
		.clock(clock),
		.io_in_a_0(r_866_0),
		.io_in_b_0(b_91_0),
		.io_in_d_0(b_1115_0),
		.io_in_control_0_dataflow(mesh_27_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2139_0),
		.io_in_last_0(r_3163_0),
		.io_in_valid_0(r_1115_0),
		.io_out_a_0(_mesh_27_2_io_out_a_0),
		.io_out_c_0(_mesh_27_2_io_out_c_0),
		.io_out_b_0(_mesh_27_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_2_io_out_id_0),
		.io_out_last_0(_mesh_27_2_io_out_last_0),
		.io_out_valid_0(_mesh_27_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10237 == GlobalFiModInstNr[0]) || (10237 == GlobalFiModInstNr[1]) || (10237 == GlobalFiModInstNr[2]) || (10237 == GlobalFiModInstNr[3]))));
	Tile mesh_27_3(
		.clock(clock),
		.io_in_a_0(r_867_0),
		.io_in_b_0(b_123_0),
		.io_in_d_0(b_1147_0),
		.io_in_control_0_dataflow(mesh_27_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2171_0),
		.io_in_last_0(r_3195_0),
		.io_in_valid_0(r_1147_0),
		.io_out_a_0(_mesh_27_3_io_out_a_0),
		.io_out_c_0(_mesh_27_3_io_out_c_0),
		.io_out_b_0(_mesh_27_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_3_io_out_id_0),
		.io_out_last_0(_mesh_27_3_io_out_last_0),
		.io_out_valid_0(_mesh_27_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10238 == GlobalFiModInstNr[0]) || (10238 == GlobalFiModInstNr[1]) || (10238 == GlobalFiModInstNr[2]) || (10238 == GlobalFiModInstNr[3]))));
	Tile mesh_27_4(
		.clock(clock),
		.io_in_a_0(r_868_0),
		.io_in_b_0(b_155_0),
		.io_in_d_0(b_1179_0),
		.io_in_control_0_dataflow(mesh_27_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2203_0),
		.io_in_last_0(r_3227_0),
		.io_in_valid_0(r_1179_0),
		.io_out_a_0(_mesh_27_4_io_out_a_0),
		.io_out_c_0(_mesh_27_4_io_out_c_0),
		.io_out_b_0(_mesh_27_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_4_io_out_id_0),
		.io_out_last_0(_mesh_27_4_io_out_last_0),
		.io_out_valid_0(_mesh_27_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10239 == GlobalFiModInstNr[0]) || (10239 == GlobalFiModInstNr[1]) || (10239 == GlobalFiModInstNr[2]) || (10239 == GlobalFiModInstNr[3]))));
	Tile mesh_27_5(
		.clock(clock),
		.io_in_a_0(r_869_0),
		.io_in_b_0(b_187_0),
		.io_in_d_0(b_1211_0),
		.io_in_control_0_dataflow(mesh_27_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2235_0),
		.io_in_last_0(r_3259_0),
		.io_in_valid_0(r_1211_0),
		.io_out_a_0(_mesh_27_5_io_out_a_0),
		.io_out_c_0(_mesh_27_5_io_out_c_0),
		.io_out_b_0(_mesh_27_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_5_io_out_id_0),
		.io_out_last_0(_mesh_27_5_io_out_last_0),
		.io_out_valid_0(_mesh_27_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10240 == GlobalFiModInstNr[0]) || (10240 == GlobalFiModInstNr[1]) || (10240 == GlobalFiModInstNr[2]) || (10240 == GlobalFiModInstNr[3]))));
	Tile mesh_27_6(
		.clock(clock),
		.io_in_a_0(r_870_0),
		.io_in_b_0(b_219_0),
		.io_in_d_0(b_1243_0),
		.io_in_control_0_dataflow(mesh_27_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2267_0),
		.io_in_last_0(r_3291_0),
		.io_in_valid_0(r_1243_0),
		.io_out_a_0(_mesh_27_6_io_out_a_0),
		.io_out_c_0(_mesh_27_6_io_out_c_0),
		.io_out_b_0(_mesh_27_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_6_io_out_id_0),
		.io_out_last_0(_mesh_27_6_io_out_last_0),
		.io_out_valid_0(_mesh_27_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10241 == GlobalFiModInstNr[0]) || (10241 == GlobalFiModInstNr[1]) || (10241 == GlobalFiModInstNr[2]) || (10241 == GlobalFiModInstNr[3]))));
	Tile mesh_27_7(
		.clock(clock),
		.io_in_a_0(r_871_0),
		.io_in_b_0(b_251_0),
		.io_in_d_0(b_1275_0),
		.io_in_control_0_dataflow(mesh_27_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2299_0),
		.io_in_last_0(r_3323_0),
		.io_in_valid_0(r_1275_0),
		.io_out_a_0(_mesh_27_7_io_out_a_0),
		.io_out_c_0(_mesh_27_7_io_out_c_0),
		.io_out_b_0(_mesh_27_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_7_io_out_id_0),
		.io_out_last_0(_mesh_27_7_io_out_last_0),
		.io_out_valid_0(_mesh_27_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10242 == GlobalFiModInstNr[0]) || (10242 == GlobalFiModInstNr[1]) || (10242 == GlobalFiModInstNr[2]) || (10242 == GlobalFiModInstNr[3]))));
	Tile mesh_27_8(
		.clock(clock),
		.io_in_a_0(r_872_0),
		.io_in_b_0(b_283_0),
		.io_in_d_0(b_1307_0),
		.io_in_control_0_dataflow(mesh_27_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2331_0),
		.io_in_last_0(r_3355_0),
		.io_in_valid_0(r_1307_0),
		.io_out_a_0(_mesh_27_8_io_out_a_0),
		.io_out_c_0(_mesh_27_8_io_out_c_0),
		.io_out_b_0(_mesh_27_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_8_io_out_id_0),
		.io_out_last_0(_mesh_27_8_io_out_last_0),
		.io_out_valid_0(_mesh_27_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10243 == GlobalFiModInstNr[0]) || (10243 == GlobalFiModInstNr[1]) || (10243 == GlobalFiModInstNr[2]) || (10243 == GlobalFiModInstNr[3]))));
	Tile mesh_27_9(
		.clock(clock),
		.io_in_a_0(r_873_0),
		.io_in_b_0(b_315_0),
		.io_in_d_0(b_1339_0),
		.io_in_control_0_dataflow(mesh_27_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2363_0),
		.io_in_last_0(r_3387_0),
		.io_in_valid_0(r_1339_0),
		.io_out_a_0(_mesh_27_9_io_out_a_0),
		.io_out_c_0(_mesh_27_9_io_out_c_0),
		.io_out_b_0(_mesh_27_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_9_io_out_id_0),
		.io_out_last_0(_mesh_27_9_io_out_last_0),
		.io_out_valid_0(_mesh_27_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10244 == GlobalFiModInstNr[0]) || (10244 == GlobalFiModInstNr[1]) || (10244 == GlobalFiModInstNr[2]) || (10244 == GlobalFiModInstNr[3]))));
	Tile mesh_27_10(
		.clock(clock),
		.io_in_a_0(r_874_0),
		.io_in_b_0(b_347_0),
		.io_in_d_0(b_1371_0),
		.io_in_control_0_dataflow(mesh_27_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2395_0),
		.io_in_last_0(r_3419_0),
		.io_in_valid_0(r_1371_0),
		.io_out_a_0(_mesh_27_10_io_out_a_0),
		.io_out_c_0(_mesh_27_10_io_out_c_0),
		.io_out_b_0(_mesh_27_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_10_io_out_id_0),
		.io_out_last_0(_mesh_27_10_io_out_last_0),
		.io_out_valid_0(_mesh_27_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10245 == GlobalFiModInstNr[0]) || (10245 == GlobalFiModInstNr[1]) || (10245 == GlobalFiModInstNr[2]) || (10245 == GlobalFiModInstNr[3]))));
	Tile mesh_27_11(
		.clock(clock),
		.io_in_a_0(r_875_0),
		.io_in_b_0(b_379_0),
		.io_in_d_0(b_1403_0),
		.io_in_control_0_dataflow(mesh_27_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2427_0),
		.io_in_last_0(r_3451_0),
		.io_in_valid_0(r_1403_0),
		.io_out_a_0(_mesh_27_11_io_out_a_0),
		.io_out_c_0(_mesh_27_11_io_out_c_0),
		.io_out_b_0(_mesh_27_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_11_io_out_id_0),
		.io_out_last_0(_mesh_27_11_io_out_last_0),
		.io_out_valid_0(_mesh_27_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10246 == GlobalFiModInstNr[0]) || (10246 == GlobalFiModInstNr[1]) || (10246 == GlobalFiModInstNr[2]) || (10246 == GlobalFiModInstNr[3]))));
	Tile mesh_27_12(
		.clock(clock),
		.io_in_a_0(r_876_0),
		.io_in_b_0(b_411_0),
		.io_in_d_0(b_1435_0),
		.io_in_control_0_dataflow(mesh_27_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2459_0),
		.io_in_last_0(r_3483_0),
		.io_in_valid_0(r_1435_0),
		.io_out_a_0(_mesh_27_12_io_out_a_0),
		.io_out_c_0(_mesh_27_12_io_out_c_0),
		.io_out_b_0(_mesh_27_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_12_io_out_id_0),
		.io_out_last_0(_mesh_27_12_io_out_last_0),
		.io_out_valid_0(_mesh_27_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10247 == GlobalFiModInstNr[0]) || (10247 == GlobalFiModInstNr[1]) || (10247 == GlobalFiModInstNr[2]) || (10247 == GlobalFiModInstNr[3]))));
	Tile mesh_27_13(
		.clock(clock),
		.io_in_a_0(r_877_0),
		.io_in_b_0(b_443_0),
		.io_in_d_0(b_1467_0),
		.io_in_control_0_dataflow(mesh_27_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2491_0),
		.io_in_last_0(r_3515_0),
		.io_in_valid_0(r_1467_0),
		.io_out_a_0(_mesh_27_13_io_out_a_0),
		.io_out_c_0(_mesh_27_13_io_out_c_0),
		.io_out_b_0(_mesh_27_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_13_io_out_id_0),
		.io_out_last_0(_mesh_27_13_io_out_last_0),
		.io_out_valid_0(_mesh_27_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10248 == GlobalFiModInstNr[0]) || (10248 == GlobalFiModInstNr[1]) || (10248 == GlobalFiModInstNr[2]) || (10248 == GlobalFiModInstNr[3]))));
	Tile mesh_27_14(
		.clock(clock),
		.io_in_a_0(r_878_0),
		.io_in_b_0(b_475_0),
		.io_in_d_0(b_1499_0),
		.io_in_control_0_dataflow(mesh_27_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2523_0),
		.io_in_last_0(r_3547_0),
		.io_in_valid_0(r_1499_0),
		.io_out_a_0(_mesh_27_14_io_out_a_0),
		.io_out_c_0(_mesh_27_14_io_out_c_0),
		.io_out_b_0(_mesh_27_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_14_io_out_id_0),
		.io_out_last_0(_mesh_27_14_io_out_last_0),
		.io_out_valid_0(_mesh_27_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10249 == GlobalFiModInstNr[0]) || (10249 == GlobalFiModInstNr[1]) || (10249 == GlobalFiModInstNr[2]) || (10249 == GlobalFiModInstNr[3]))));
	Tile mesh_27_15(
		.clock(clock),
		.io_in_a_0(r_879_0),
		.io_in_b_0(b_507_0),
		.io_in_d_0(b_1531_0),
		.io_in_control_0_dataflow(mesh_27_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2555_0),
		.io_in_last_0(r_3579_0),
		.io_in_valid_0(r_1531_0),
		.io_out_a_0(_mesh_27_15_io_out_a_0),
		.io_out_c_0(_mesh_27_15_io_out_c_0),
		.io_out_b_0(_mesh_27_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_15_io_out_id_0),
		.io_out_last_0(_mesh_27_15_io_out_last_0),
		.io_out_valid_0(_mesh_27_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10250 == GlobalFiModInstNr[0]) || (10250 == GlobalFiModInstNr[1]) || (10250 == GlobalFiModInstNr[2]) || (10250 == GlobalFiModInstNr[3]))));
	Tile mesh_27_16(
		.clock(clock),
		.io_in_a_0(r_880_0),
		.io_in_b_0(b_539_0),
		.io_in_d_0(b_1563_0),
		.io_in_control_0_dataflow(mesh_27_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2587_0),
		.io_in_last_0(r_3611_0),
		.io_in_valid_0(r_1563_0),
		.io_out_a_0(_mesh_27_16_io_out_a_0),
		.io_out_c_0(_mesh_27_16_io_out_c_0),
		.io_out_b_0(_mesh_27_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_16_io_out_id_0),
		.io_out_last_0(_mesh_27_16_io_out_last_0),
		.io_out_valid_0(_mesh_27_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10251 == GlobalFiModInstNr[0]) || (10251 == GlobalFiModInstNr[1]) || (10251 == GlobalFiModInstNr[2]) || (10251 == GlobalFiModInstNr[3]))));
	Tile mesh_27_17(
		.clock(clock),
		.io_in_a_0(r_881_0),
		.io_in_b_0(b_571_0),
		.io_in_d_0(b_1595_0),
		.io_in_control_0_dataflow(mesh_27_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2619_0),
		.io_in_last_0(r_3643_0),
		.io_in_valid_0(r_1595_0),
		.io_out_a_0(_mesh_27_17_io_out_a_0),
		.io_out_c_0(_mesh_27_17_io_out_c_0),
		.io_out_b_0(_mesh_27_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_17_io_out_id_0),
		.io_out_last_0(_mesh_27_17_io_out_last_0),
		.io_out_valid_0(_mesh_27_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10252 == GlobalFiModInstNr[0]) || (10252 == GlobalFiModInstNr[1]) || (10252 == GlobalFiModInstNr[2]) || (10252 == GlobalFiModInstNr[3]))));
	Tile mesh_27_18(
		.clock(clock),
		.io_in_a_0(r_882_0),
		.io_in_b_0(b_603_0),
		.io_in_d_0(b_1627_0),
		.io_in_control_0_dataflow(mesh_27_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2651_0),
		.io_in_last_0(r_3675_0),
		.io_in_valid_0(r_1627_0),
		.io_out_a_0(_mesh_27_18_io_out_a_0),
		.io_out_c_0(_mesh_27_18_io_out_c_0),
		.io_out_b_0(_mesh_27_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_18_io_out_id_0),
		.io_out_last_0(_mesh_27_18_io_out_last_0),
		.io_out_valid_0(_mesh_27_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10253 == GlobalFiModInstNr[0]) || (10253 == GlobalFiModInstNr[1]) || (10253 == GlobalFiModInstNr[2]) || (10253 == GlobalFiModInstNr[3]))));
	Tile mesh_27_19(
		.clock(clock),
		.io_in_a_0(r_883_0),
		.io_in_b_0(b_635_0),
		.io_in_d_0(b_1659_0),
		.io_in_control_0_dataflow(mesh_27_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2683_0),
		.io_in_last_0(r_3707_0),
		.io_in_valid_0(r_1659_0),
		.io_out_a_0(_mesh_27_19_io_out_a_0),
		.io_out_c_0(_mesh_27_19_io_out_c_0),
		.io_out_b_0(_mesh_27_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_19_io_out_id_0),
		.io_out_last_0(_mesh_27_19_io_out_last_0),
		.io_out_valid_0(_mesh_27_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10254 == GlobalFiModInstNr[0]) || (10254 == GlobalFiModInstNr[1]) || (10254 == GlobalFiModInstNr[2]) || (10254 == GlobalFiModInstNr[3]))));
	Tile mesh_27_20(
		.clock(clock),
		.io_in_a_0(r_884_0),
		.io_in_b_0(b_667_0),
		.io_in_d_0(b_1691_0),
		.io_in_control_0_dataflow(mesh_27_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2715_0),
		.io_in_last_0(r_3739_0),
		.io_in_valid_0(r_1691_0),
		.io_out_a_0(_mesh_27_20_io_out_a_0),
		.io_out_c_0(_mesh_27_20_io_out_c_0),
		.io_out_b_0(_mesh_27_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_20_io_out_id_0),
		.io_out_last_0(_mesh_27_20_io_out_last_0),
		.io_out_valid_0(_mesh_27_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10255 == GlobalFiModInstNr[0]) || (10255 == GlobalFiModInstNr[1]) || (10255 == GlobalFiModInstNr[2]) || (10255 == GlobalFiModInstNr[3]))));
	Tile mesh_27_21(
		.clock(clock),
		.io_in_a_0(r_885_0),
		.io_in_b_0(b_699_0),
		.io_in_d_0(b_1723_0),
		.io_in_control_0_dataflow(mesh_27_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2747_0),
		.io_in_last_0(r_3771_0),
		.io_in_valid_0(r_1723_0),
		.io_out_a_0(_mesh_27_21_io_out_a_0),
		.io_out_c_0(_mesh_27_21_io_out_c_0),
		.io_out_b_0(_mesh_27_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_21_io_out_id_0),
		.io_out_last_0(_mesh_27_21_io_out_last_0),
		.io_out_valid_0(_mesh_27_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10256 == GlobalFiModInstNr[0]) || (10256 == GlobalFiModInstNr[1]) || (10256 == GlobalFiModInstNr[2]) || (10256 == GlobalFiModInstNr[3]))));
	Tile mesh_27_22(
		.clock(clock),
		.io_in_a_0(r_886_0),
		.io_in_b_0(b_731_0),
		.io_in_d_0(b_1755_0),
		.io_in_control_0_dataflow(mesh_27_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2779_0),
		.io_in_last_0(r_3803_0),
		.io_in_valid_0(r_1755_0),
		.io_out_a_0(_mesh_27_22_io_out_a_0),
		.io_out_c_0(_mesh_27_22_io_out_c_0),
		.io_out_b_0(_mesh_27_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_22_io_out_id_0),
		.io_out_last_0(_mesh_27_22_io_out_last_0),
		.io_out_valid_0(_mesh_27_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10257 == GlobalFiModInstNr[0]) || (10257 == GlobalFiModInstNr[1]) || (10257 == GlobalFiModInstNr[2]) || (10257 == GlobalFiModInstNr[3]))));
	Tile mesh_27_23(
		.clock(clock),
		.io_in_a_0(r_887_0),
		.io_in_b_0(b_763_0),
		.io_in_d_0(b_1787_0),
		.io_in_control_0_dataflow(mesh_27_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2811_0),
		.io_in_last_0(r_3835_0),
		.io_in_valid_0(r_1787_0),
		.io_out_a_0(_mesh_27_23_io_out_a_0),
		.io_out_c_0(_mesh_27_23_io_out_c_0),
		.io_out_b_0(_mesh_27_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_23_io_out_id_0),
		.io_out_last_0(_mesh_27_23_io_out_last_0),
		.io_out_valid_0(_mesh_27_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10258 == GlobalFiModInstNr[0]) || (10258 == GlobalFiModInstNr[1]) || (10258 == GlobalFiModInstNr[2]) || (10258 == GlobalFiModInstNr[3]))));
	Tile mesh_27_24(
		.clock(clock),
		.io_in_a_0(r_888_0),
		.io_in_b_0(b_795_0),
		.io_in_d_0(b_1819_0),
		.io_in_control_0_dataflow(mesh_27_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2843_0),
		.io_in_last_0(r_3867_0),
		.io_in_valid_0(r_1819_0),
		.io_out_a_0(_mesh_27_24_io_out_a_0),
		.io_out_c_0(_mesh_27_24_io_out_c_0),
		.io_out_b_0(_mesh_27_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_24_io_out_id_0),
		.io_out_last_0(_mesh_27_24_io_out_last_0),
		.io_out_valid_0(_mesh_27_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10259 == GlobalFiModInstNr[0]) || (10259 == GlobalFiModInstNr[1]) || (10259 == GlobalFiModInstNr[2]) || (10259 == GlobalFiModInstNr[3]))));
	Tile mesh_27_25(
		.clock(clock),
		.io_in_a_0(r_889_0),
		.io_in_b_0(b_827_0),
		.io_in_d_0(b_1851_0),
		.io_in_control_0_dataflow(mesh_27_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2875_0),
		.io_in_last_0(r_3899_0),
		.io_in_valid_0(r_1851_0),
		.io_out_a_0(_mesh_27_25_io_out_a_0),
		.io_out_c_0(_mesh_27_25_io_out_c_0),
		.io_out_b_0(_mesh_27_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_25_io_out_id_0),
		.io_out_last_0(_mesh_27_25_io_out_last_0),
		.io_out_valid_0(_mesh_27_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10260 == GlobalFiModInstNr[0]) || (10260 == GlobalFiModInstNr[1]) || (10260 == GlobalFiModInstNr[2]) || (10260 == GlobalFiModInstNr[3]))));
	Tile mesh_27_26(
		.clock(clock),
		.io_in_a_0(r_890_0),
		.io_in_b_0(b_859_0),
		.io_in_d_0(b_1883_0),
		.io_in_control_0_dataflow(mesh_27_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2907_0),
		.io_in_last_0(r_3931_0),
		.io_in_valid_0(r_1883_0),
		.io_out_a_0(_mesh_27_26_io_out_a_0),
		.io_out_c_0(_mesh_27_26_io_out_c_0),
		.io_out_b_0(_mesh_27_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_26_io_out_id_0),
		.io_out_last_0(_mesh_27_26_io_out_last_0),
		.io_out_valid_0(_mesh_27_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10261 == GlobalFiModInstNr[0]) || (10261 == GlobalFiModInstNr[1]) || (10261 == GlobalFiModInstNr[2]) || (10261 == GlobalFiModInstNr[3]))));
	Tile mesh_27_27(
		.clock(clock),
		.io_in_a_0(r_891_0),
		.io_in_b_0(b_891_0),
		.io_in_d_0(b_1915_0),
		.io_in_control_0_dataflow(mesh_27_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2939_0),
		.io_in_last_0(r_3963_0),
		.io_in_valid_0(r_1915_0),
		.io_out_a_0(_mesh_27_27_io_out_a_0),
		.io_out_c_0(_mesh_27_27_io_out_c_0),
		.io_out_b_0(_mesh_27_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_27_io_out_id_0),
		.io_out_last_0(_mesh_27_27_io_out_last_0),
		.io_out_valid_0(_mesh_27_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10262 == GlobalFiModInstNr[0]) || (10262 == GlobalFiModInstNr[1]) || (10262 == GlobalFiModInstNr[2]) || (10262 == GlobalFiModInstNr[3]))));
	Tile mesh_27_28(
		.clock(clock),
		.io_in_a_0(r_892_0),
		.io_in_b_0(b_923_0),
		.io_in_d_0(b_1947_0),
		.io_in_control_0_dataflow(mesh_27_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2971_0),
		.io_in_last_0(r_3995_0),
		.io_in_valid_0(r_1947_0),
		.io_out_a_0(_mesh_27_28_io_out_a_0),
		.io_out_c_0(_mesh_27_28_io_out_c_0),
		.io_out_b_0(_mesh_27_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_28_io_out_id_0),
		.io_out_last_0(_mesh_27_28_io_out_last_0),
		.io_out_valid_0(_mesh_27_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10263 == GlobalFiModInstNr[0]) || (10263 == GlobalFiModInstNr[1]) || (10263 == GlobalFiModInstNr[2]) || (10263 == GlobalFiModInstNr[3]))));
	Tile mesh_27_29(
		.clock(clock),
		.io_in_a_0(r_893_0),
		.io_in_b_0(b_955_0),
		.io_in_d_0(b_1979_0),
		.io_in_control_0_dataflow(mesh_27_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3003_0),
		.io_in_last_0(r_4027_0),
		.io_in_valid_0(r_1979_0),
		.io_out_a_0(_mesh_27_29_io_out_a_0),
		.io_out_c_0(_mesh_27_29_io_out_c_0),
		.io_out_b_0(_mesh_27_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_29_io_out_id_0),
		.io_out_last_0(_mesh_27_29_io_out_last_0),
		.io_out_valid_0(_mesh_27_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10264 == GlobalFiModInstNr[0]) || (10264 == GlobalFiModInstNr[1]) || (10264 == GlobalFiModInstNr[2]) || (10264 == GlobalFiModInstNr[3]))));
	Tile mesh_27_30(
		.clock(clock),
		.io_in_a_0(r_894_0),
		.io_in_b_0(b_987_0),
		.io_in_d_0(b_2011_0),
		.io_in_control_0_dataflow(mesh_27_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3035_0),
		.io_in_last_0(r_4059_0),
		.io_in_valid_0(r_2011_0),
		.io_out_a_0(_mesh_27_30_io_out_a_0),
		.io_out_c_0(_mesh_27_30_io_out_c_0),
		.io_out_b_0(_mesh_27_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_30_io_out_id_0),
		.io_out_last_0(_mesh_27_30_io_out_last_0),
		.io_out_valid_0(_mesh_27_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10265 == GlobalFiModInstNr[0]) || (10265 == GlobalFiModInstNr[1]) || (10265 == GlobalFiModInstNr[2]) || (10265 == GlobalFiModInstNr[3]))));
	Tile mesh_27_31(
		.clock(clock),
		.io_in_a_0(r_895_0),
		.io_in_b_0(b_1019_0),
		.io_in_d_0(b_2043_0),
		.io_in_control_0_dataflow(mesh_27_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_27_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_27_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3067_0),
		.io_in_last_0(r_4091_0),
		.io_in_valid_0(r_2043_0),
		.io_out_a_0(_mesh_27_31_io_out_a_0),
		.io_out_c_0(_mesh_27_31_io_out_c_0),
		.io_out_b_0(_mesh_27_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_27_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_27_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_27_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_27_31_io_out_id_0),
		.io_out_last_0(_mesh_27_31_io_out_last_0),
		.io_out_valid_0(_mesh_27_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10266 == GlobalFiModInstNr[0]) || (10266 == GlobalFiModInstNr[1]) || (10266 == GlobalFiModInstNr[2]) || (10266 == GlobalFiModInstNr[3]))));
	Tile mesh_28_0(
		.clock(clock),
		.io_in_a_0(r_896_0),
		.io_in_b_0(b_28_0),
		.io_in_d_0(b_1052_0),
		.io_in_control_0_dataflow(mesh_28_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2076_0),
		.io_in_last_0(r_3100_0),
		.io_in_valid_0(r_1052_0),
		.io_out_a_0(_mesh_28_0_io_out_a_0),
		.io_out_c_0(_mesh_28_0_io_out_c_0),
		.io_out_b_0(_mesh_28_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_0_io_out_id_0),
		.io_out_last_0(_mesh_28_0_io_out_last_0),
		.io_out_valid_0(_mesh_28_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10267 == GlobalFiModInstNr[0]) || (10267 == GlobalFiModInstNr[1]) || (10267 == GlobalFiModInstNr[2]) || (10267 == GlobalFiModInstNr[3]))));
	Tile mesh_28_1(
		.clock(clock),
		.io_in_a_0(r_897_0),
		.io_in_b_0(b_60_0),
		.io_in_d_0(b_1084_0),
		.io_in_control_0_dataflow(mesh_28_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2108_0),
		.io_in_last_0(r_3132_0),
		.io_in_valid_0(r_1084_0),
		.io_out_a_0(_mesh_28_1_io_out_a_0),
		.io_out_c_0(_mesh_28_1_io_out_c_0),
		.io_out_b_0(_mesh_28_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_1_io_out_id_0),
		.io_out_last_0(_mesh_28_1_io_out_last_0),
		.io_out_valid_0(_mesh_28_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10268 == GlobalFiModInstNr[0]) || (10268 == GlobalFiModInstNr[1]) || (10268 == GlobalFiModInstNr[2]) || (10268 == GlobalFiModInstNr[3]))));
	Tile mesh_28_2(
		.clock(clock),
		.io_in_a_0(r_898_0),
		.io_in_b_0(b_92_0),
		.io_in_d_0(b_1116_0),
		.io_in_control_0_dataflow(mesh_28_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2140_0),
		.io_in_last_0(r_3164_0),
		.io_in_valid_0(r_1116_0),
		.io_out_a_0(_mesh_28_2_io_out_a_0),
		.io_out_c_0(_mesh_28_2_io_out_c_0),
		.io_out_b_0(_mesh_28_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_2_io_out_id_0),
		.io_out_last_0(_mesh_28_2_io_out_last_0),
		.io_out_valid_0(_mesh_28_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10269 == GlobalFiModInstNr[0]) || (10269 == GlobalFiModInstNr[1]) || (10269 == GlobalFiModInstNr[2]) || (10269 == GlobalFiModInstNr[3]))));
	Tile mesh_28_3(
		.clock(clock),
		.io_in_a_0(r_899_0),
		.io_in_b_0(b_124_0),
		.io_in_d_0(b_1148_0),
		.io_in_control_0_dataflow(mesh_28_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2172_0),
		.io_in_last_0(r_3196_0),
		.io_in_valid_0(r_1148_0),
		.io_out_a_0(_mesh_28_3_io_out_a_0),
		.io_out_c_0(_mesh_28_3_io_out_c_0),
		.io_out_b_0(_mesh_28_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_3_io_out_id_0),
		.io_out_last_0(_mesh_28_3_io_out_last_0),
		.io_out_valid_0(_mesh_28_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10270 == GlobalFiModInstNr[0]) || (10270 == GlobalFiModInstNr[1]) || (10270 == GlobalFiModInstNr[2]) || (10270 == GlobalFiModInstNr[3]))));
	Tile mesh_28_4(
		.clock(clock),
		.io_in_a_0(r_900_0),
		.io_in_b_0(b_156_0),
		.io_in_d_0(b_1180_0),
		.io_in_control_0_dataflow(mesh_28_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2204_0),
		.io_in_last_0(r_3228_0),
		.io_in_valid_0(r_1180_0),
		.io_out_a_0(_mesh_28_4_io_out_a_0),
		.io_out_c_0(_mesh_28_4_io_out_c_0),
		.io_out_b_0(_mesh_28_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_4_io_out_id_0),
		.io_out_last_0(_mesh_28_4_io_out_last_0),
		.io_out_valid_0(_mesh_28_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10271 == GlobalFiModInstNr[0]) || (10271 == GlobalFiModInstNr[1]) || (10271 == GlobalFiModInstNr[2]) || (10271 == GlobalFiModInstNr[3]))));
	Tile mesh_28_5(
		.clock(clock),
		.io_in_a_0(r_901_0),
		.io_in_b_0(b_188_0),
		.io_in_d_0(b_1212_0),
		.io_in_control_0_dataflow(mesh_28_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2236_0),
		.io_in_last_0(r_3260_0),
		.io_in_valid_0(r_1212_0),
		.io_out_a_0(_mesh_28_5_io_out_a_0),
		.io_out_c_0(_mesh_28_5_io_out_c_0),
		.io_out_b_0(_mesh_28_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_5_io_out_id_0),
		.io_out_last_0(_mesh_28_5_io_out_last_0),
		.io_out_valid_0(_mesh_28_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10272 == GlobalFiModInstNr[0]) || (10272 == GlobalFiModInstNr[1]) || (10272 == GlobalFiModInstNr[2]) || (10272 == GlobalFiModInstNr[3]))));
	Tile mesh_28_6(
		.clock(clock),
		.io_in_a_0(r_902_0),
		.io_in_b_0(b_220_0),
		.io_in_d_0(b_1244_0),
		.io_in_control_0_dataflow(mesh_28_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2268_0),
		.io_in_last_0(r_3292_0),
		.io_in_valid_0(r_1244_0),
		.io_out_a_0(_mesh_28_6_io_out_a_0),
		.io_out_c_0(_mesh_28_6_io_out_c_0),
		.io_out_b_0(_mesh_28_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_6_io_out_id_0),
		.io_out_last_0(_mesh_28_6_io_out_last_0),
		.io_out_valid_0(_mesh_28_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10273 == GlobalFiModInstNr[0]) || (10273 == GlobalFiModInstNr[1]) || (10273 == GlobalFiModInstNr[2]) || (10273 == GlobalFiModInstNr[3]))));
	Tile mesh_28_7(
		.clock(clock),
		.io_in_a_0(r_903_0),
		.io_in_b_0(b_252_0),
		.io_in_d_0(b_1276_0),
		.io_in_control_0_dataflow(mesh_28_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2300_0),
		.io_in_last_0(r_3324_0),
		.io_in_valid_0(r_1276_0),
		.io_out_a_0(_mesh_28_7_io_out_a_0),
		.io_out_c_0(_mesh_28_7_io_out_c_0),
		.io_out_b_0(_mesh_28_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_7_io_out_id_0),
		.io_out_last_0(_mesh_28_7_io_out_last_0),
		.io_out_valid_0(_mesh_28_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10274 == GlobalFiModInstNr[0]) || (10274 == GlobalFiModInstNr[1]) || (10274 == GlobalFiModInstNr[2]) || (10274 == GlobalFiModInstNr[3]))));
	Tile mesh_28_8(
		.clock(clock),
		.io_in_a_0(r_904_0),
		.io_in_b_0(b_284_0),
		.io_in_d_0(b_1308_0),
		.io_in_control_0_dataflow(mesh_28_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2332_0),
		.io_in_last_0(r_3356_0),
		.io_in_valid_0(r_1308_0),
		.io_out_a_0(_mesh_28_8_io_out_a_0),
		.io_out_c_0(_mesh_28_8_io_out_c_0),
		.io_out_b_0(_mesh_28_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_8_io_out_id_0),
		.io_out_last_0(_mesh_28_8_io_out_last_0),
		.io_out_valid_0(_mesh_28_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10275 == GlobalFiModInstNr[0]) || (10275 == GlobalFiModInstNr[1]) || (10275 == GlobalFiModInstNr[2]) || (10275 == GlobalFiModInstNr[3]))));
	Tile mesh_28_9(
		.clock(clock),
		.io_in_a_0(r_905_0),
		.io_in_b_0(b_316_0),
		.io_in_d_0(b_1340_0),
		.io_in_control_0_dataflow(mesh_28_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2364_0),
		.io_in_last_0(r_3388_0),
		.io_in_valid_0(r_1340_0),
		.io_out_a_0(_mesh_28_9_io_out_a_0),
		.io_out_c_0(_mesh_28_9_io_out_c_0),
		.io_out_b_0(_mesh_28_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_9_io_out_id_0),
		.io_out_last_0(_mesh_28_9_io_out_last_0),
		.io_out_valid_0(_mesh_28_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10276 == GlobalFiModInstNr[0]) || (10276 == GlobalFiModInstNr[1]) || (10276 == GlobalFiModInstNr[2]) || (10276 == GlobalFiModInstNr[3]))));
	Tile mesh_28_10(
		.clock(clock),
		.io_in_a_0(r_906_0),
		.io_in_b_0(b_348_0),
		.io_in_d_0(b_1372_0),
		.io_in_control_0_dataflow(mesh_28_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2396_0),
		.io_in_last_0(r_3420_0),
		.io_in_valid_0(r_1372_0),
		.io_out_a_0(_mesh_28_10_io_out_a_0),
		.io_out_c_0(_mesh_28_10_io_out_c_0),
		.io_out_b_0(_mesh_28_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_10_io_out_id_0),
		.io_out_last_0(_mesh_28_10_io_out_last_0),
		.io_out_valid_0(_mesh_28_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10277 == GlobalFiModInstNr[0]) || (10277 == GlobalFiModInstNr[1]) || (10277 == GlobalFiModInstNr[2]) || (10277 == GlobalFiModInstNr[3]))));
	Tile mesh_28_11(
		.clock(clock),
		.io_in_a_0(r_907_0),
		.io_in_b_0(b_380_0),
		.io_in_d_0(b_1404_0),
		.io_in_control_0_dataflow(mesh_28_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2428_0),
		.io_in_last_0(r_3452_0),
		.io_in_valid_0(r_1404_0),
		.io_out_a_0(_mesh_28_11_io_out_a_0),
		.io_out_c_0(_mesh_28_11_io_out_c_0),
		.io_out_b_0(_mesh_28_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_11_io_out_id_0),
		.io_out_last_0(_mesh_28_11_io_out_last_0),
		.io_out_valid_0(_mesh_28_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10278 == GlobalFiModInstNr[0]) || (10278 == GlobalFiModInstNr[1]) || (10278 == GlobalFiModInstNr[2]) || (10278 == GlobalFiModInstNr[3]))));
	Tile mesh_28_12(
		.clock(clock),
		.io_in_a_0(r_908_0),
		.io_in_b_0(b_412_0),
		.io_in_d_0(b_1436_0),
		.io_in_control_0_dataflow(mesh_28_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2460_0),
		.io_in_last_0(r_3484_0),
		.io_in_valid_0(r_1436_0),
		.io_out_a_0(_mesh_28_12_io_out_a_0),
		.io_out_c_0(_mesh_28_12_io_out_c_0),
		.io_out_b_0(_mesh_28_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_12_io_out_id_0),
		.io_out_last_0(_mesh_28_12_io_out_last_0),
		.io_out_valid_0(_mesh_28_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10279 == GlobalFiModInstNr[0]) || (10279 == GlobalFiModInstNr[1]) || (10279 == GlobalFiModInstNr[2]) || (10279 == GlobalFiModInstNr[3]))));
	Tile mesh_28_13(
		.clock(clock),
		.io_in_a_0(r_909_0),
		.io_in_b_0(b_444_0),
		.io_in_d_0(b_1468_0),
		.io_in_control_0_dataflow(mesh_28_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2492_0),
		.io_in_last_0(r_3516_0),
		.io_in_valid_0(r_1468_0),
		.io_out_a_0(_mesh_28_13_io_out_a_0),
		.io_out_c_0(_mesh_28_13_io_out_c_0),
		.io_out_b_0(_mesh_28_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_13_io_out_id_0),
		.io_out_last_0(_mesh_28_13_io_out_last_0),
		.io_out_valid_0(_mesh_28_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10280 == GlobalFiModInstNr[0]) || (10280 == GlobalFiModInstNr[1]) || (10280 == GlobalFiModInstNr[2]) || (10280 == GlobalFiModInstNr[3]))));
	Tile mesh_28_14(
		.clock(clock),
		.io_in_a_0(r_910_0),
		.io_in_b_0(b_476_0),
		.io_in_d_0(b_1500_0),
		.io_in_control_0_dataflow(mesh_28_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2524_0),
		.io_in_last_0(r_3548_0),
		.io_in_valid_0(r_1500_0),
		.io_out_a_0(_mesh_28_14_io_out_a_0),
		.io_out_c_0(_mesh_28_14_io_out_c_0),
		.io_out_b_0(_mesh_28_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_14_io_out_id_0),
		.io_out_last_0(_mesh_28_14_io_out_last_0),
		.io_out_valid_0(_mesh_28_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10281 == GlobalFiModInstNr[0]) || (10281 == GlobalFiModInstNr[1]) || (10281 == GlobalFiModInstNr[2]) || (10281 == GlobalFiModInstNr[3]))));
	Tile mesh_28_15(
		.clock(clock),
		.io_in_a_0(r_911_0),
		.io_in_b_0(b_508_0),
		.io_in_d_0(b_1532_0),
		.io_in_control_0_dataflow(mesh_28_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2556_0),
		.io_in_last_0(r_3580_0),
		.io_in_valid_0(r_1532_0),
		.io_out_a_0(_mesh_28_15_io_out_a_0),
		.io_out_c_0(_mesh_28_15_io_out_c_0),
		.io_out_b_0(_mesh_28_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_15_io_out_id_0),
		.io_out_last_0(_mesh_28_15_io_out_last_0),
		.io_out_valid_0(_mesh_28_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10282 == GlobalFiModInstNr[0]) || (10282 == GlobalFiModInstNr[1]) || (10282 == GlobalFiModInstNr[2]) || (10282 == GlobalFiModInstNr[3]))));
	Tile mesh_28_16(
		.clock(clock),
		.io_in_a_0(r_912_0),
		.io_in_b_0(b_540_0),
		.io_in_d_0(b_1564_0),
		.io_in_control_0_dataflow(mesh_28_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2588_0),
		.io_in_last_0(r_3612_0),
		.io_in_valid_0(r_1564_0),
		.io_out_a_0(_mesh_28_16_io_out_a_0),
		.io_out_c_0(_mesh_28_16_io_out_c_0),
		.io_out_b_0(_mesh_28_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_16_io_out_id_0),
		.io_out_last_0(_mesh_28_16_io_out_last_0),
		.io_out_valid_0(_mesh_28_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10283 == GlobalFiModInstNr[0]) || (10283 == GlobalFiModInstNr[1]) || (10283 == GlobalFiModInstNr[2]) || (10283 == GlobalFiModInstNr[3]))));
	Tile mesh_28_17(
		.clock(clock),
		.io_in_a_0(r_913_0),
		.io_in_b_0(b_572_0),
		.io_in_d_0(b_1596_0),
		.io_in_control_0_dataflow(mesh_28_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2620_0),
		.io_in_last_0(r_3644_0),
		.io_in_valid_0(r_1596_0),
		.io_out_a_0(_mesh_28_17_io_out_a_0),
		.io_out_c_0(_mesh_28_17_io_out_c_0),
		.io_out_b_0(_mesh_28_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_17_io_out_id_0),
		.io_out_last_0(_mesh_28_17_io_out_last_0),
		.io_out_valid_0(_mesh_28_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10284 == GlobalFiModInstNr[0]) || (10284 == GlobalFiModInstNr[1]) || (10284 == GlobalFiModInstNr[2]) || (10284 == GlobalFiModInstNr[3]))));
	Tile mesh_28_18(
		.clock(clock),
		.io_in_a_0(r_914_0),
		.io_in_b_0(b_604_0),
		.io_in_d_0(b_1628_0),
		.io_in_control_0_dataflow(mesh_28_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2652_0),
		.io_in_last_0(r_3676_0),
		.io_in_valid_0(r_1628_0),
		.io_out_a_0(_mesh_28_18_io_out_a_0),
		.io_out_c_0(_mesh_28_18_io_out_c_0),
		.io_out_b_0(_mesh_28_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_18_io_out_id_0),
		.io_out_last_0(_mesh_28_18_io_out_last_0),
		.io_out_valid_0(_mesh_28_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10285 == GlobalFiModInstNr[0]) || (10285 == GlobalFiModInstNr[1]) || (10285 == GlobalFiModInstNr[2]) || (10285 == GlobalFiModInstNr[3]))));
	Tile mesh_28_19(
		.clock(clock),
		.io_in_a_0(r_915_0),
		.io_in_b_0(b_636_0),
		.io_in_d_0(b_1660_0),
		.io_in_control_0_dataflow(mesh_28_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2684_0),
		.io_in_last_0(r_3708_0),
		.io_in_valid_0(r_1660_0),
		.io_out_a_0(_mesh_28_19_io_out_a_0),
		.io_out_c_0(_mesh_28_19_io_out_c_0),
		.io_out_b_0(_mesh_28_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_19_io_out_id_0),
		.io_out_last_0(_mesh_28_19_io_out_last_0),
		.io_out_valid_0(_mesh_28_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10286 == GlobalFiModInstNr[0]) || (10286 == GlobalFiModInstNr[1]) || (10286 == GlobalFiModInstNr[2]) || (10286 == GlobalFiModInstNr[3]))));
	Tile mesh_28_20(
		.clock(clock),
		.io_in_a_0(r_916_0),
		.io_in_b_0(b_668_0),
		.io_in_d_0(b_1692_0),
		.io_in_control_0_dataflow(mesh_28_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2716_0),
		.io_in_last_0(r_3740_0),
		.io_in_valid_0(r_1692_0),
		.io_out_a_0(_mesh_28_20_io_out_a_0),
		.io_out_c_0(_mesh_28_20_io_out_c_0),
		.io_out_b_0(_mesh_28_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_20_io_out_id_0),
		.io_out_last_0(_mesh_28_20_io_out_last_0),
		.io_out_valid_0(_mesh_28_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10287 == GlobalFiModInstNr[0]) || (10287 == GlobalFiModInstNr[1]) || (10287 == GlobalFiModInstNr[2]) || (10287 == GlobalFiModInstNr[3]))));
	Tile mesh_28_21(
		.clock(clock),
		.io_in_a_0(r_917_0),
		.io_in_b_0(b_700_0),
		.io_in_d_0(b_1724_0),
		.io_in_control_0_dataflow(mesh_28_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2748_0),
		.io_in_last_0(r_3772_0),
		.io_in_valid_0(r_1724_0),
		.io_out_a_0(_mesh_28_21_io_out_a_0),
		.io_out_c_0(_mesh_28_21_io_out_c_0),
		.io_out_b_0(_mesh_28_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_21_io_out_id_0),
		.io_out_last_0(_mesh_28_21_io_out_last_0),
		.io_out_valid_0(_mesh_28_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10288 == GlobalFiModInstNr[0]) || (10288 == GlobalFiModInstNr[1]) || (10288 == GlobalFiModInstNr[2]) || (10288 == GlobalFiModInstNr[3]))));
	Tile mesh_28_22(
		.clock(clock),
		.io_in_a_0(r_918_0),
		.io_in_b_0(b_732_0),
		.io_in_d_0(b_1756_0),
		.io_in_control_0_dataflow(mesh_28_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2780_0),
		.io_in_last_0(r_3804_0),
		.io_in_valid_0(r_1756_0),
		.io_out_a_0(_mesh_28_22_io_out_a_0),
		.io_out_c_0(_mesh_28_22_io_out_c_0),
		.io_out_b_0(_mesh_28_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_22_io_out_id_0),
		.io_out_last_0(_mesh_28_22_io_out_last_0),
		.io_out_valid_0(_mesh_28_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10289 == GlobalFiModInstNr[0]) || (10289 == GlobalFiModInstNr[1]) || (10289 == GlobalFiModInstNr[2]) || (10289 == GlobalFiModInstNr[3]))));
	Tile mesh_28_23(
		.clock(clock),
		.io_in_a_0(r_919_0),
		.io_in_b_0(b_764_0),
		.io_in_d_0(b_1788_0),
		.io_in_control_0_dataflow(mesh_28_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2812_0),
		.io_in_last_0(r_3836_0),
		.io_in_valid_0(r_1788_0),
		.io_out_a_0(_mesh_28_23_io_out_a_0),
		.io_out_c_0(_mesh_28_23_io_out_c_0),
		.io_out_b_0(_mesh_28_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_23_io_out_id_0),
		.io_out_last_0(_mesh_28_23_io_out_last_0),
		.io_out_valid_0(_mesh_28_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10290 == GlobalFiModInstNr[0]) || (10290 == GlobalFiModInstNr[1]) || (10290 == GlobalFiModInstNr[2]) || (10290 == GlobalFiModInstNr[3]))));
	Tile mesh_28_24(
		.clock(clock),
		.io_in_a_0(r_920_0),
		.io_in_b_0(b_796_0),
		.io_in_d_0(b_1820_0),
		.io_in_control_0_dataflow(mesh_28_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2844_0),
		.io_in_last_0(r_3868_0),
		.io_in_valid_0(r_1820_0),
		.io_out_a_0(_mesh_28_24_io_out_a_0),
		.io_out_c_0(_mesh_28_24_io_out_c_0),
		.io_out_b_0(_mesh_28_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_24_io_out_id_0),
		.io_out_last_0(_mesh_28_24_io_out_last_0),
		.io_out_valid_0(_mesh_28_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10291 == GlobalFiModInstNr[0]) || (10291 == GlobalFiModInstNr[1]) || (10291 == GlobalFiModInstNr[2]) || (10291 == GlobalFiModInstNr[3]))));
	Tile mesh_28_25(
		.clock(clock),
		.io_in_a_0(r_921_0),
		.io_in_b_0(b_828_0),
		.io_in_d_0(b_1852_0),
		.io_in_control_0_dataflow(mesh_28_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2876_0),
		.io_in_last_0(r_3900_0),
		.io_in_valid_0(r_1852_0),
		.io_out_a_0(_mesh_28_25_io_out_a_0),
		.io_out_c_0(_mesh_28_25_io_out_c_0),
		.io_out_b_0(_mesh_28_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_25_io_out_id_0),
		.io_out_last_0(_mesh_28_25_io_out_last_0),
		.io_out_valid_0(_mesh_28_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10292 == GlobalFiModInstNr[0]) || (10292 == GlobalFiModInstNr[1]) || (10292 == GlobalFiModInstNr[2]) || (10292 == GlobalFiModInstNr[3]))));
	Tile mesh_28_26(
		.clock(clock),
		.io_in_a_0(r_922_0),
		.io_in_b_0(b_860_0),
		.io_in_d_0(b_1884_0),
		.io_in_control_0_dataflow(mesh_28_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2908_0),
		.io_in_last_0(r_3932_0),
		.io_in_valid_0(r_1884_0),
		.io_out_a_0(_mesh_28_26_io_out_a_0),
		.io_out_c_0(_mesh_28_26_io_out_c_0),
		.io_out_b_0(_mesh_28_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_26_io_out_id_0),
		.io_out_last_0(_mesh_28_26_io_out_last_0),
		.io_out_valid_0(_mesh_28_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10293 == GlobalFiModInstNr[0]) || (10293 == GlobalFiModInstNr[1]) || (10293 == GlobalFiModInstNr[2]) || (10293 == GlobalFiModInstNr[3]))));
	Tile mesh_28_27(
		.clock(clock),
		.io_in_a_0(r_923_0),
		.io_in_b_0(b_892_0),
		.io_in_d_0(b_1916_0),
		.io_in_control_0_dataflow(mesh_28_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2940_0),
		.io_in_last_0(r_3964_0),
		.io_in_valid_0(r_1916_0),
		.io_out_a_0(_mesh_28_27_io_out_a_0),
		.io_out_c_0(_mesh_28_27_io_out_c_0),
		.io_out_b_0(_mesh_28_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_27_io_out_id_0),
		.io_out_last_0(_mesh_28_27_io_out_last_0),
		.io_out_valid_0(_mesh_28_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10294 == GlobalFiModInstNr[0]) || (10294 == GlobalFiModInstNr[1]) || (10294 == GlobalFiModInstNr[2]) || (10294 == GlobalFiModInstNr[3]))));
	Tile mesh_28_28(
		.clock(clock),
		.io_in_a_0(r_924_0),
		.io_in_b_0(b_924_0),
		.io_in_d_0(b_1948_0),
		.io_in_control_0_dataflow(mesh_28_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2972_0),
		.io_in_last_0(r_3996_0),
		.io_in_valid_0(r_1948_0),
		.io_out_a_0(_mesh_28_28_io_out_a_0),
		.io_out_c_0(_mesh_28_28_io_out_c_0),
		.io_out_b_0(_mesh_28_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_28_io_out_id_0),
		.io_out_last_0(_mesh_28_28_io_out_last_0),
		.io_out_valid_0(_mesh_28_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10295 == GlobalFiModInstNr[0]) || (10295 == GlobalFiModInstNr[1]) || (10295 == GlobalFiModInstNr[2]) || (10295 == GlobalFiModInstNr[3]))));
	Tile mesh_28_29(
		.clock(clock),
		.io_in_a_0(r_925_0),
		.io_in_b_0(b_956_0),
		.io_in_d_0(b_1980_0),
		.io_in_control_0_dataflow(mesh_28_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3004_0),
		.io_in_last_0(r_4028_0),
		.io_in_valid_0(r_1980_0),
		.io_out_a_0(_mesh_28_29_io_out_a_0),
		.io_out_c_0(_mesh_28_29_io_out_c_0),
		.io_out_b_0(_mesh_28_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_29_io_out_id_0),
		.io_out_last_0(_mesh_28_29_io_out_last_0),
		.io_out_valid_0(_mesh_28_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10296 == GlobalFiModInstNr[0]) || (10296 == GlobalFiModInstNr[1]) || (10296 == GlobalFiModInstNr[2]) || (10296 == GlobalFiModInstNr[3]))));
	Tile mesh_28_30(
		.clock(clock),
		.io_in_a_0(r_926_0),
		.io_in_b_0(b_988_0),
		.io_in_d_0(b_2012_0),
		.io_in_control_0_dataflow(mesh_28_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3036_0),
		.io_in_last_0(r_4060_0),
		.io_in_valid_0(r_2012_0),
		.io_out_a_0(_mesh_28_30_io_out_a_0),
		.io_out_c_0(_mesh_28_30_io_out_c_0),
		.io_out_b_0(_mesh_28_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_30_io_out_id_0),
		.io_out_last_0(_mesh_28_30_io_out_last_0),
		.io_out_valid_0(_mesh_28_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10297 == GlobalFiModInstNr[0]) || (10297 == GlobalFiModInstNr[1]) || (10297 == GlobalFiModInstNr[2]) || (10297 == GlobalFiModInstNr[3]))));
	Tile mesh_28_31(
		.clock(clock),
		.io_in_a_0(r_927_0),
		.io_in_b_0(b_1020_0),
		.io_in_d_0(b_2044_0),
		.io_in_control_0_dataflow(mesh_28_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_28_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_28_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3068_0),
		.io_in_last_0(r_4092_0),
		.io_in_valid_0(r_2044_0),
		.io_out_a_0(_mesh_28_31_io_out_a_0),
		.io_out_c_0(_mesh_28_31_io_out_c_0),
		.io_out_b_0(_mesh_28_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_28_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_28_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_28_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_28_31_io_out_id_0),
		.io_out_last_0(_mesh_28_31_io_out_last_0),
		.io_out_valid_0(_mesh_28_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10298 == GlobalFiModInstNr[0]) || (10298 == GlobalFiModInstNr[1]) || (10298 == GlobalFiModInstNr[2]) || (10298 == GlobalFiModInstNr[3]))));
	Tile mesh_29_0(
		.clock(clock),
		.io_in_a_0(r_928_0),
		.io_in_b_0(b_29_0),
		.io_in_d_0(b_1053_0),
		.io_in_control_0_dataflow(mesh_29_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2077_0),
		.io_in_last_0(r_3101_0),
		.io_in_valid_0(r_1053_0),
		.io_out_a_0(_mesh_29_0_io_out_a_0),
		.io_out_c_0(_mesh_29_0_io_out_c_0),
		.io_out_b_0(_mesh_29_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_0_io_out_id_0),
		.io_out_last_0(_mesh_29_0_io_out_last_0),
		.io_out_valid_0(_mesh_29_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10299 == GlobalFiModInstNr[0]) || (10299 == GlobalFiModInstNr[1]) || (10299 == GlobalFiModInstNr[2]) || (10299 == GlobalFiModInstNr[3]))));
	Tile mesh_29_1(
		.clock(clock),
		.io_in_a_0(r_929_0),
		.io_in_b_0(b_61_0),
		.io_in_d_0(b_1085_0),
		.io_in_control_0_dataflow(mesh_29_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2109_0),
		.io_in_last_0(r_3133_0),
		.io_in_valid_0(r_1085_0),
		.io_out_a_0(_mesh_29_1_io_out_a_0),
		.io_out_c_0(_mesh_29_1_io_out_c_0),
		.io_out_b_0(_mesh_29_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_1_io_out_id_0),
		.io_out_last_0(_mesh_29_1_io_out_last_0),
		.io_out_valid_0(_mesh_29_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10300 == GlobalFiModInstNr[0]) || (10300 == GlobalFiModInstNr[1]) || (10300 == GlobalFiModInstNr[2]) || (10300 == GlobalFiModInstNr[3]))));
	Tile mesh_29_2(
		.clock(clock),
		.io_in_a_0(r_930_0),
		.io_in_b_0(b_93_0),
		.io_in_d_0(b_1117_0),
		.io_in_control_0_dataflow(mesh_29_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2141_0),
		.io_in_last_0(r_3165_0),
		.io_in_valid_0(r_1117_0),
		.io_out_a_0(_mesh_29_2_io_out_a_0),
		.io_out_c_0(_mesh_29_2_io_out_c_0),
		.io_out_b_0(_mesh_29_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_2_io_out_id_0),
		.io_out_last_0(_mesh_29_2_io_out_last_0),
		.io_out_valid_0(_mesh_29_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10301 == GlobalFiModInstNr[0]) || (10301 == GlobalFiModInstNr[1]) || (10301 == GlobalFiModInstNr[2]) || (10301 == GlobalFiModInstNr[3]))));
	Tile mesh_29_3(
		.clock(clock),
		.io_in_a_0(r_931_0),
		.io_in_b_0(b_125_0),
		.io_in_d_0(b_1149_0),
		.io_in_control_0_dataflow(mesh_29_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2173_0),
		.io_in_last_0(r_3197_0),
		.io_in_valid_0(r_1149_0),
		.io_out_a_0(_mesh_29_3_io_out_a_0),
		.io_out_c_0(_mesh_29_3_io_out_c_0),
		.io_out_b_0(_mesh_29_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_3_io_out_id_0),
		.io_out_last_0(_mesh_29_3_io_out_last_0),
		.io_out_valid_0(_mesh_29_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10302 == GlobalFiModInstNr[0]) || (10302 == GlobalFiModInstNr[1]) || (10302 == GlobalFiModInstNr[2]) || (10302 == GlobalFiModInstNr[3]))));
	Tile mesh_29_4(
		.clock(clock),
		.io_in_a_0(r_932_0),
		.io_in_b_0(b_157_0),
		.io_in_d_0(b_1181_0),
		.io_in_control_0_dataflow(mesh_29_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2205_0),
		.io_in_last_0(r_3229_0),
		.io_in_valid_0(r_1181_0),
		.io_out_a_0(_mesh_29_4_io_out_a_0),
		.io_out_c_0(_mesh_29_4_io_out_c_0),
		.io_out_b_0(_mesh_29_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_4_io_out_id_0),
		.io_out_last_0(_mesh_29_4_io_out_last_0),
		.io_out_valid_0(_mesh_29_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10303 == GlobalFiModInstNr[0]) || (10303 == GlobalFiModInstNr[1]) || (10303 == GlobalFiModInstNr[2]) || (10303 == GlobalFiModInstNr[3]))));
	Tile mesh_29_5(
		.clock(clock),
		.io_in_a_0(r_933_0),
		.io_in_b_0(b_189_0),
		.io_in_d_0(b_1213_0),
		.io_in_control_0_dataflow(mesh_29_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2237_0),
		.io_in_last_0(r_3261_0),
		.io_in_valid_0(r_1213_0),
		.io_out_a_0(_mesh_29_5_io_out_a_0),
		.io_out_c_0(_mesh_29_5_io_out_c_0),
		.io_out_b_0(_mesh_29_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_5_io_out_id_0),
		.io_out_last_0(_mesh_29_5_io_out_last_0),
		.io_out_valid_0(_mesh_29_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10304 == GlobalFiModInstNr[0]) || (10304 == GlobalFiModInstNr[1]) || (10304 == GlobalFiModInstNr[2]) || (10304 == GlobalFiModInstNr[3]))));
	Tile mesh_29_6(
		.clock(clock),
		.io_in_a_0(r_934_0),
		.io_in_b_0(b_221_0),
		.io_in_d_0(b_1245_0),
		.io_in_control_0_dataflow(mesh_29_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2269_0),
		.io_in_last_0(r_3293_0),
		.io_in_valid_0(r_1245_0),
		.io_out_a_0(_mesh_29_6_io_out_a_0),
		.io_out_c_0(_mesh_29_6_io_out_c_0),
		.io_out_b_0(_mesh_29_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_6_io_out_id_0),
		.io_out_last_0(_mesh_29_6_io_out_last_0),
		.io_out_valid_0(_mesh_29_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10305 == GlobalFiModInstNr[0]) || (10305 == GlobalFiModInstNr[1]) || (10305 == GlobalFiModInstNr[2]) || (10305 == GlobalFiModInstNr[3]))));
	Tile mesh_29_7(
		.clock(clock),
		.io_in_a_0(r_935_0),
		.io_in_b_0(b_253_0),
		.io_in_d_0(b_1277_0),
		.io_in_control_0_dataflow(mesh_29_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2301_0),
		.io_in_last_0(r_3325_0),
		.io_in_valid_0(r_1277_0),
		.io_out_a_0(_mesh_29_7_io_out_a_0),
		.io_out_c_0(_mesh_29_7_io_out_c_0),
		.io_out_b_0(_mesh_29_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_7_io_out_id_0),
		.io_out_last_0(_mesh_29_7_io_out_last_0),
		.io_out_valid_0(_mesh_29_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10306 == GlobalFiModInstNr[0]) || (10306 == GlobalFiModInstNr[1]) || (10306 == GlobalFiModInstNr[2]) || (10306 == GlobalFiModInstNr[3]))));
	Tile mesh_29_8(
		.clock(clock),
		.io_in_a_0(r_936_0),
		.io_in_b_0(b_285_0),
		.io_in_d_0(b_1309_0),
		.io_in_control_0_dataflow(mesh_29_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2333_0),
		.io_in_last_0(r_3357_0),
		.io_in_valid_0(r_1309_0),
		.io_out_a_0(_mesh_29_8_io_out_a_0),
		.io_out_c_0(_mesh_29_8_io_out_c_0),
		.io_out_b_0(_mesh_29_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_8_io_out_id_0),
		.io_out_last_0(_mesh_29_8_io_out_last_0),
		.io_out_valid_0(_mesh_29_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10307 == GlobalFiModInstNr[0]) || (10307 == GlobalFiModInstNr[1]) || (10307 == GlobalFiModInstNr[2]) || (10307 == GlobalFiModInstNr[3]))));
	Tile mesh_29_9(
		.clock(clock),
		.io_in_a_0(r_937_0),
		.io_in_b_0(b_317_0),
		.io_in_d_0(b_1341_0),
		.io_in_control_0_dataflow(mesh_29_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2365_0),
		.io_in_last_0(r_3389_0),
		.io_in_valid_0(r_1341_0),
		.io_out_a_0(_mesh_29_9_io_out_a_0),
		.io_out_c_0(_mesh_29_9_io_out_c_0),
		.io_out_b_0(_mesh_29_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_9_io_out_id_0),
		.io_out_last_0(_mesh_29_9_io_out_last_0),
		.io_out_valid_0(_mesh_29_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10308 == GlobalFiModInstNr[0]) || (10308 == GlobalFiModInstNr[1]) || (10308 == GlobalFiModInstNr[2]) || (10308 == GlobalFiModInstNr[3]))));
	Tile mesh_29_10(
		.clock(clock),
		.io_in_a_0(r_938_0),
		.io_in_b_0(b_349_0),
		.io_in_d_0(b_1373_0),
		.io_in_control_0_dataflow(mesh_29_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2397_0),
		.io_in_last_0(r_3421_0),
		.io_in_valid_0(r_1373_0),
		.io_out_a_0(_mesh_29_10_io_out_a_0),
		.io_out_c_0(_mesh_29_10_io_out_c_0),
		.io_out_b_0(_mesh_29_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_10_io_out_id_0),
		.io_out_last_0(_mesh_29_10_io_out_last_0),
		.io_out_valid_0(_mesh_29_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10309 == GlobalFiModInstNr[0]) || (10309 == GlobalFiModInstNr[1]) || (10309 == GlobalFiModInstNr[2]) || (10309 == GlobalFiModInstNr[3]))));
	Tile mesh_29_11(
		.clock(clock),
		.io_in_a_0(r_939_0),
		.io_in_b_0(b_381_0),
		.io_in_d_0(b_1405_0),
		.io_in_control_0_dataflow(mesh_29_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2429_0),
		.io_in_last_0(r_3453_0),
		.io_in_valid_0(r_1405_0),
		.io_out_a_0(_mesh_29_11_io_out_a_0),
		.io_out_c_0(_mesh_29_11_io_out_c_0),
		.io_out_b_0(_mesh_29_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_11_io_out_id_0),
		.io_out_last_0(_mesh_29_11_io_out_last_0),
		.io_out_valid_0(_mesh_29_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10310 == GlobalFiModInstNr[0]) || (10310 == GlobalFiModInstNr[1]) || (10310 == GlobalFiModInstNr[2]) || (10310 == GlobalFiModInstNr[3]))));
	Tile mesh_29_12(
		.clock(clock),
		.io_in_a_0(r_940_0),
		.io_in_b_0(b_413_0),
		.io_in_d_0(b_1437_0),
		.io_in_control_0_dataflow(mesh_29_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2461_0),
		.io_in_last_0(r_3485_0),
		.io_in_valid_0(r_1437_0),
		.io_out_a_0(_mesh_29_12_io_out_a_0),
		.io_out_c_0(_mesh_29_12_io_out_c_0),
		.io_out_b_0(_mesh_29_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_12_io_out_id_0),
		.io_out_last_0(_mesh_29_12_io_out_last_0),
		.io_out_valid_0(_mesh_29_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10311 == GlobalFiModInstNr[0]) || (10311 == GlobalFiModInstNr[1]) || (10311 == GlobalFiModInstNr[2]) || (10311 == GlobalFiModInstNr[3]))));
	Tile mesh_29_13(
		.clock(clock),
		.io_in_a_0(r_941_0),
		.io_in_b_0(b_445_0),
		.io_in_d_0(b_1469_0),
		.io_in_control_0_dataflow(mesh_29_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2493_0),
		.io_in_last_0(r_3517_0),
		.io_in_valid_0(r_1469_0),
		.io_out_a_0(_mesh_29_13_io_out_a_0),
		.io_out_c_0(_mesh_29_13_io_out_c_0),
		.io_out_b_0(_mesh_29_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_13_io_out_id_0),
		.io_out_last_0(_mesh_29_13_io_out_last_0),
		.io_out_valid_0(_mesh_29_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10312 == GlobalFiModInstNr[0]) || (10312 == GlobalFiModInstNr[1]) || (10312 == GlobalFiModInstNr[2]) || (10312 == GlobalFiModInstNr[3]))));
	Tile mesh_29_14(
		.clock(clock),
		.io_in_a_0(r_942_0),
		.io_in_b_0(b_477_0),
		.io_in_d_0(b_1501_0),
		.io_in_control_0_dataflow(mesh_29_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2525_0),
		.io_in_last_0(r_3549_0),
		.io_in_valid_0(r_1501_0),
		.io_out_a_0(_mesh_29_14_io_out_a_0),
		.io_out_c_0(_mesh_29_14_io_out_c_0),
		.io_out_b_0(_mesh_29_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_14_io_out_id_0),
		.io_out_last_0(_mesh_29_14_io_out_last_0),
		.io_out_valid_0(_mesh_29_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10313 == GlobalFiModInstNr[0]) || (10313 == GlobalFiModInstNr[1]) || (10313 == GlobalFiModInstNr[2]) || (10313 == GlobalFiModInstNr[3]))));
	Tile mesh_29_15(
		.clock(clock),
		.io_in_a_0(r_943_0),
		.io_in_b_0(b_509_0),
		.io_in_d_0(b_1533_0),
		.io_in_control_0_dataflow(mesh_29_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2557_0),
		.io_in_last_0(r_3581_0),
		.io_in_valid_0(r_1533_0),
		.io_out_a_0(_mesh_29_15_io_out_a_0),
		.io_out_c_0(_mesh_29_15_io_out_c_0),
		.io_out_b_0(_mesh_29_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_15_io_out_id_0),
		.io_out_last_0(_mesh_29_15_io_out_last_0),
		.io_out_valid_0(_mesh_29_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10314 == GlobalFiModInstNr[0]) || (10314 == GlobalFiModInstNr[1]) || (10314 == GlobalFiModInstNr[2]) || (10314 == GlobalFiModInstNr[3]))));
	Tile mesh_29_16(
		.clock(clock),
		.io_in_a_0(r_944_0),
		.io_in_b_0(b_541_0),
		.io_in_d_0(b_1565_0),
		.io_in_control_0_dataflow(mesh_29_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2589_0),
		.io_in_last_0(r_3613_0),
		.io_in_valid_0(r_1565_0),
		.io_out_a_0(_mesh_29_16_io_out_a_0),
		.io_out_c_0(_mesh_29_16_io_out_c_0),
		.io_out_b_0(_mesh_29_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_16_io_out_id_0),
		.io_out_last_0(_mesh_29_16_io_out_last_0),
		.io_out_valid_0(_mesh_29_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10315 == GlobalFiModInstNr[0]) || (10315 == GlobalFiModInstNr[1]) || (10315 == GlobalFiModInstNr[2]) || (10315 == GlobalFiModInstNr[3]))));
	Tile mesh_29_17(
		.clock(clock),
		.io_in_a_0(r_945_0),
		.io_in_b_0(b_573_0),
		.io_in_d_0(b_1597_0),
		.io_in_control_0_dataflow(mesh_29_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2621_0),
		.io_in_last_0(r_3645_0),
		.io_in_valid_0(r_1597_0),
		.io_out_a_0(_mesh_29_17_io_out_a_0),
		.io_out_c_0(_mesh_29_17_io_out_c_0),
		.io_out_b_0(_mesh_29_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_17_io_out_id_0),
		.io_out_last_0(_mesh_29_17_io_out_last_0),
		.io_out_valid_0(_mesh_29_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10316 == GlobalFiModInstNr[0]) || (10316 == GlobalFiModInstNr[1]) || (10316 == GlobalFiModInstNr[2]) || (10316 == GlobalFiModInstNr[3]))));
	Tile mesh_29_18(
		.clock(clock),
		.io_in_a_0(r_946_0),
		.io_in_b_0(b_605_0),
		.io_in_d_0(b_1629_0),
		.io_in_control_0_dataflow(mesh_29_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2653_0),
		.io_in_last_0(r_3677_0),
		.io_in_valid_0(r_1629_0),
		.io_out_a_0(_mesh_29_18_io_out_a_0),
		.io_out_c_0(_mesh_29_18_io_out_c_0),
		.io_out_b_0(_mesh_29_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_18_io_out_id_0),
		.io_out_last_0(_mesh_29_18_io_out_last_0),
		.io_out_valid_0(_mesh_29_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10317 == GlobalFiModInstNr[0]) || (10317 == GlobalFiModInstNr[1]) || (10317 == GlobalFiModInstNr[2]) || (10317 == GlobalFiModInstNr[3]))));
	Tile mesh_29_19(
		.clock(clock),
		.io_in_a_0(r_947_0),
		.io_in_b_0(b_637_0),
		.io_in_d_0(b_1661_0),
		.io_in_control_0_dataflow(mesh_29_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2685_0),
		.io_in_last_0(r_3709_0),
		.io_in_valid_0(r_1661_0),
		.io_out_a_0(_mesh_29_19_io_out_a_0),
		.io_out_c_0(_mesh_29_19_io_out_c_0),
		.io_out_b_0(_mesh_29_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_19_io_out_id_0),
		.io_out_last_0(_mesh_29_19_io_out_last_0),
		.io_out_valid_0(_mesh_29_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10318 == GlobalFiModInstNr[0]) || (10318 == GlobalFiModInstNr[1]) || (10318 == GlobalFiModInstNr[2]) || (10318 == GlobalFiModInstNr[3]))));
	Tile mesh_29_20(
		.clock(clock),
		.io_in_a_0(r_948_0),
		.io_in_b_0(b_669_0),
		.io_in_d_0(b_1693_0),
		.io_in_control_0_dataflow(mesh_29_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2717_0),
		.io_in_last_0(r_3741_0),
		.io_in_valid_0(r_1693_0),
		.io_out_a_0(_mesh_29_20_io_out_a_0),
		.io_out_c_0(_mesh_29_20_io_out_c_0),
		.io_out_b_0(_mesh_29_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_20_io_out_id_0),
		.io_out_last_0(_mesh_29_20_io_out_last_0),
		.io_out_valid_0(_mesh_29_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10319 == GlobalFiModInstNr[0]) || (10319 == GlobalFiModInstNr[1]) || (10319 == GlobalFiModInstNr[2]) || (10319 == GlobalFiModInstNr[3]))));
	Tile mesh_29_21(
		.clock(clock),
		.io_in_a_0(r_949_0),
		.io_in_b_0(b_701_0),
		.io_in_d_0(b_1725_0),
		.io_in_control_0_dataflow(mesh_29_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2749_0),
		.io_in_last_0(r_3773_0),
		.io_in_valid_0(r_1725_0),
		.io_out_a_0(_mesh_29_21_io_out_a_0),
		.io_out_c_0(_mesh_29_21_io_out_c_0),
		.io_out_b_0(_mesh_29_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_21_io_out_id_0),
		.io_out_last_0(_mesh_29_21_io_out_last_0),
		.io_out_valid_0(_mesh_29_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10320 == GlobalFiModInstNr[0]) || (10320 == GlobalFiModInstNr[1]) || (10320 == GlobalFiModInstNr[2]) || (10320 == GlobalFiModInstNr[3]))));
	Tile mesh_29_22(
		.clock(clock),
		.io_in_a_0(r_950_0),
		.io_in_b_0(b_733_0),
		.io_in_d_0(b_1757_0),
		.io_in_control_0_dataflow(mesh_29_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2781_0),
		.io_in_last_0(r_3805_0),
		.io_in_valid_0(r_1757_0),
		.io_out_a_0(_mesh_29_22_io_out_a_0),
		.io_out_c_0(_mesh_29_22_io_out_c_0),
		.io_out_b_0(_mesh_29_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_22_io_out_id_0),
		.io_out_last_0(_mesh_29_22_io_out_last_0),
		.io_out_valid_0(_mesh_29_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10321 == GlobalFiModInstNr[0]) || (10321 == GlobalFiModInstNr[1]) || (10321 == GlobalFiModInstNr[2]) || (10321 == GlobalFiModInstNr[3]))));
	Tile mesh_29_23(
		.clock(clock),
		.io_in_a_0(r_951_0),
		.io_in_b_0(b_765_0),
		.io_in_d_0(b_1789_0),
		.io_in_control_0_dataflow(mesh_29_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2813_0),
		.io_in_last_0(r_3837_0),
		.io_in_valid_0(r_1789_0),
		.io_out_a_0(_mesh_29_23_io_out_a_0),
		.io_out_c_0(_mesh_29_23_io_out_c_0),
		.io_out_b_0(_mesh_29_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_23_io_out_id_0),
		.io_out_last_0(_mesh_29_23_io_out_last_0),
		.io_out_valid_0(_mesh_29_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10322 == GlobalFiModInstNr[0]) || (10322 == GlobalFiModInstNr[1]) || (10322 == GlobalFiModInstNr[2]) || (10322 == GlobalFiModInstNr[3]))));
	Tile mesh_29_24(
		.clock(clock),
		.io_in_a_0(r_952_0),
		.io_in_b_0(b_797_0),
		.io_in_d_0(b_1821_0),
		.io_in_control_0_dataflow(mesh_29_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2845_0),
		.io_in_last_0(r_3869_0),
		.io_in_valid_0(r_1821_0),
		.io_out_a_0(_mesh_29_24_io_out_a_0),
		.io_out_c_0(_mesh_29_24_io_out_c_0),
		.io_out_b_0(_mesh_29_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_24_io_out_id_0),
		.io_out_last_0(_mesh_29_24_io_out_last_0),
		.io_out_valid_0(_mesh_29_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10323 == GlobalFiModInstNr[0]) || (10323 == GlobalFiModInstNr[1]) || (10323 == GlobalFiModInstNr[2]) || (10323 == GlobalFiModInstNr[3]))));
	Tile mesh_29_25(
		.clock(clock),
		.io_in_a_0(r_953_0),
		.io_in_b_0(b_829_0),
		.io_in_d_0(b_1853_0),
		.io_in_control_0_dataflow(mesh_29_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2877_0),
		.io_in_last_0(r_3901_0),
		.io_in_valid_0(r_1853_0),
		.io_out_a_0(_mesh_29_25_io_out_a_0),
		.io_out_c_0(_mesh_29_25_io_out_c_0),
		.io_out_b_0(_mesh_29_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_25_io_out_id_0),
		.io_out_last_0(_mesh_29_25_io_out_last_0),
		.io_out_valid_0(_mesh_29_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10324 == GlobalFiModInstNr[0]) || (10324 == GlobalFiModInstNr[1]) || (10324 == GlobalFiModInstNr[2]) || (10324 == GlobalFiModInstNr[3]))));
	Tile mesh_29_26(
		.clock(clock),
		.io_in_a_0(r_954_0),
		.io_in_b_0(b_861_0),
		.io_in_d_0(b_1885_0),
		.io_in_control_0_dataflow(mesh_29_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2909_0),
		.io_in_last_0(r_3933_0),
		.io_in_valid_0(r_1885_0),
		.io_out_a_0(_mesh_29_26_io_out_a_0),
		.io_out_c_0(_mesh_29_26_io_out_c_0),
		.io_out_b_0(_mesh_29_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_26_io_out_id_0),
		.io_out_last_0(_mesh_29_26_io_out_last_0),
		.io_out_valid_0(_mesh_29_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10325 == GlobalFiModInstNr[0]) || (10325 == GlobalFiModInstNr[1]) || (10325 == GlobalFiModInstNr[2]) || (10325 == GlobalFiModInstNr[3]))));
	Tile mesh_29_27(
		.clock(clock),
		.io_in_a_0(r_955_0),
		.io_in_b_0(b_893_0),
		.io_in_d_0(b_1917_0),
		.io_in_control_0_dataflow(mesh_29_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2941_0),
		.io_in_last_0(r_3965_0),
		.io_in_valid_0(r_1917_0),
		.io_out_a_0(_mesh_29_27_io_out_a_0),
		.io_out_c_0(_mesh_29_27_io_out_c_0),
		.io_out_b_0(_mesh_29_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_27_io_out_id_0),
		.io_out_last_0(_mesh_29_27_io_out_last_0),
		.io_out_valid_0(_mesh_29_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10326 == GlobalFiModInstNr[0]) || (10326 == GlobalFiModInstNr[1]) || (10326 == GlobalFiModInstNr[2]) || (10326 == GlobalFiModInstNr[3]))));
	Tile mesh_29_28(
		.clock(clock),
		.io_in_a_0(r_956_0),
		.io_in_b_0(b_925_0),
		.io_in_d_0(b_1949_0),
		.io_in_control_0_dataflow(mesh_29_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2973_0),
		.io_in_last_0(r_3997_0),
		.io_in_valid_0(r_1949_0),
		.io_out_a_0(_mesh_29_28_io_out_a_0),
		.io_out_c_0(_mesh_29_28_io_out_c_0),
		.io_out_b_0(_mesh_29_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_28_io_out_id_0),
		.io_out_last_0(_mesh_29_28_io_out_last_0),
		.io_out_valid_0(_mesh_29_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10327 == GlobalFiModInstNr[0]) || (10327 == GlobalFiModInstNr[1]) || (10327 == GlobalFiModInstNr[2]) || (10327 == GlobalFiModInstNr[3]))));
	Tile mesh_29_29(
		.clock(clock),
		.io_in_a_0(r_957_0),
		.io_in_b_0(b_957_0),
		.io_in_d_0(b_1981_0),
		.io_in_control_0_dataflow(mesh_29_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3005_0),
		.io_in_last_0(r_4029_0),
		.io_in_valid_0(r_1981_0),
		.io_out_a_0(_mesh_29_29_io_out_a_0),
		.io_out_c_0(_mesh_29_29_io_out_c_0),
		.io_out_b_0(_mesh_29_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_29_io_out_id_0),
		.io_out_last_0(_mesh_29_29_io_out_last_0),
		.io_out_valid_0(_mesh_29_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10328 == GlobalFiModInstNr[0]) || (10328 == GlobalFiModInstNr[1]) || (10328 == GlobalFiModInstNr[2]) || (10328 == GlobalFiModInstNr[3]))));
	Tile mesh_29_30(
		.clock(clock),
		.io_in_a_0(r_958_0),
		.io_in_b_0(b_989_0),
		.io_in_d_0(b_2013_0),
		.io_in_control_0_dataflow(mesh_29_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3037_0),
		.io_in_last_0(r_4061_0),
		.io_in_valid_0(r_2013_0),
		.io_out_a_0(_mesh_29_30_io_out_a_0),
		.io_out_c_0(_mesh_29_30_io_out_c_0),
		.io_out_b_0(_mesh_29_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_30_io_out_id_0),
		.io_out_last_0(_mesh_29_30_io_out_last_0),
		.io_out_valid_0(_mesh_29_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10329 == GlobalFiModInstNr[0]) || (10329 == GlobalFiModInstNr[1]) || (10329 == GlobalFiModInstNr[2]) || (10329 == GlobalFiModInstNr[3]))));
	Tile mesh_29_31(
		.clock(clock),
		.io_in_a_0(r_959_0),
		.io_in_b_0(b_1021_0),
		.io_in_d_0(b_2045_0),
		.io_in_control_0_dataflow(mesh_29_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_29_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_29_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3069_0),
		.io_in_last_0(r_4093_0),
		.io_in_valid_0(r_2045_0),
		.io_out_a_0(_mesh_29_31_io_out_a_0),
		.io_out_c_0(_mesh_29_31_io_out_c_0),
		.io_out_b_0(_mesh_29_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_29_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_29_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_29_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_29_31_io_out_id_0),
		.io_out_last_0(_mesh_29_31_io_out_last_0),
		.io_out_valid_0(_mesh_29_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10330 == GlobalFiModInstNr[0]) || (10330 == GlobalFiModInstNr[1]) || (10330 == GlobalFiModInstNr[2]) || (10330 == GlobalFiModInstNr[3]))));
	Tile mesh_30_0(
		.clock(clock),
		.io_in_a_0(r_960_0),
		.io_in_b_0(b_30_0),
		.io_in_d_0(b_1054_0),
		.io_in_control_0_dataflow(mesh_30_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2078_0),
		.io_in_last_0(r_3102_0),
		.io_in_valid_0(r_1054_0),
		.io_out_a_0(_mesh_30_0_io_out_a_0),
		.io_out_c_0(_mesh_30_0_io_out_c_0),
		.io_out_b_0(_mesh_30_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_0_io_out_id_0),
		.io_out_last_0(_mesh_30_0_io_out_last_0),
		.io_out_valid_0(_mesh_30_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10331 == GlobalFiModInstNr[0]) || (10331 == GlobalFiModInstNr[1]) || (10331 == GlobalFiModInstNr[2]) || (10331 == GlobalFiModInstNr[3]))));
	Tile mesh_30_1(
		.clock(clock),
		.io_in_a_0(r_961_0),
		.io_in_b_0(b_62_0),
		.io_in_d_0(b_1086_0),
		.io_in_control_0_dataflow(mesh_30_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2110_0),
		.io_in_last_0(r_3134_0),
		.io_in_valid_0(r_1086_0),
		.io_out_a_0(_mesh_30_1_io_out_a_0),
		.io_out_c_0(_mesh_30_1_io_out_c_0),
		.io_out_b_0(_mesh_30_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_1_io_out_id_0),
		.io_out_last_0(_mesh_30_1_io_out_last_0),
		.io_out_valid_0(_mesh_30_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10332 == GlobalFiModInstNr[0]) || (10332 == GlobalFiModInstNr[1]) || (10332 == GlobalFiModInstNr[2]) || (10332 == GlobalFiModInstNr[3]))));
	Tile mesh_30_2(
		.clock(clock),
		.io_in_a_0(r_962_0),
		.io_in_b_0(b_94_0),
		.io_in_d_0(b_1118_0),
		.io_in_control_0_dataflow(mesh_30_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2142_0),
		.io_in_last_0(r_3166_0),
		.io_in_valid_0(r_1118_0),
		.io_out_a_0(_mesh_30_2_io_out_a_0),
		.io_out_c_0(_mesh_30_2_io_out_c_0),
		.io_out_b_0(_mesh_30_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_2_io_out_id_0),
		.io_out_last_0(_mesh_30_2_io_out_last_0),
		.io_out_valid_0(_mesh_30_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10333 == GlobalFiModInstNr[0]) || (10333 == GlobalFiModInstNr[1]) || (10333 == GlobalFiModInstNr[2]) || (10333 == GlobalFiModInstNr[3]))));
	Tile mesh_30_3(
		.clock(clock),
		.io_in_a_0(r_963_0),
		.io_in_b_0(b_126_0),
		.io_in_d_0(b_1150_0),
		.io_in_control_0_dataflow(mesh_30_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2174_0),
		.io_in_last_0(r_3198_0),
		.io_in_valid_0(r_1150_0),
		.io_out_a_0(_mesh_30_3_io_out_a_0),
		.io_out_c_0(_mesh_30_3_io_out_c_0),
		.io_out_b_0(_mesh_30_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_3_io_out_id_0),
		.io_out_last_0(_mesh_30_3_io_out_last_0),
		.io_out_valid_0(_mesh_30_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10334 == GlobalFiModInstNr[0]) || (10334 == GlobalFiModInstNr[1]) || (10334 == GlobalFiModInstNr[2]) || (10334 == GlobalFiModInstNr[3]))));
	Tile mesh_30_4(
		.clock(clock),
		.io_in_a_0(r_964_0),
		.io_in_b_0(b_158_0),
		.io_in_d_0(b_1182_0),
		.io_in_control_0_dataflow(mesh_30_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2206_0),
		.io_in_last_0(r_3230_0),
		.io_in_valid_0(r_1182_0),
		.io_out_a_0(_mesh_30_4_io_out_a_0),
		.io_out_c_0(_mesh_30_4_io_out_c_0),
		.io_out_b_0(_mesh_30_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_4_io_out_id_0),
		.io_out_last_0(_mesh_30_4_io_out_last_0),
		.io_out_valid_0(_mesh_30_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10335 == GlobalFiModInstNr[0]) || (10335 == GlobalFiModInstNr[1]) || (10335 == GlobalFiModInstNr[2]) || (10335 == GlobalFiModInstNr[3]))));
	Tile mesh_30_5(
		.clock(clock),
		.io_in_a_0(r_965_0),
		.io_in_b_0(b_190_0),
		.io_in_d_0(b_1214_0),
		.io_in_control_0_dataflow(mesh_30_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2238_0),
		.io_in_last_0(r_3262_0),
		.io_in_valid_0(r_1214_0),
		.io_out_a_0(_mesh_30_5_io_out_a_0),
		.io_out_c_0(_mesh_30_5_io_out_c_0),
		.io_out_b_0(_mesh_30_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_5_io_out_id_0),
		.io_out_last_0(_mesh_30_5_io_out_last_0),
		.io_out_valid_0(_mesh_30_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10336 == GlobalFiModInstNr[0]) || (10336 == GlobalFiModInstNr[1]) || (10336 == GlobalFiModInstNr[2]) || (10336 == GlobalFiModInstNr[3]))));
	Tile mesh_30_6(
		.clock(clock),
		.io_in_a_0(r_966_0),
		.io_in_b_0(b_222_0),
		.io_in_d_0(b_1246_0),
		.io_in_control_0_dataflow(mesh_30_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2270_0),
		.io_in_last_0(r_3294_0),
		.io_in_valid_0(r_1246_0),
		.io_out_a_0(_mesh_30_6_io_out_a_0),
		.io_out_c_0(_mesh_30_6_io_out_c_0),
		.io_out_b_0(_mesh_30_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_6_io_out_id_0),
		.io_out_last_0(_mesh_30_6_io_out_last_0),
		.io_out_valid_0(_mesh_30_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10337 == GlobalFiModInstNr[0]) || (10337 == GlobalFiModInstNr[1]) || (10337 == GlobalFiModInstNr[2]) || (10337 == GlobalFiModInstNr[3]))));
	Tile mesh_30_7(
		.clock(clock),
		.io_in_a_0(r_967_0),
		.io_in_b_0(b_254_0),
		.io_in_d_0(b_1278_0),
		.io_in_control_0_dataflow(mesh_30_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2302_0),
		.io_in_last_0(r_3326_0),
		.io_in_valid_0(r_1278_0),
		.io_out_a_0(_mesh_30_7_io_out_a_0),
		.io_out_c_0(_mesh_30_7_io_out_c_0),
		.io_out_b_0(_mesh_30_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_7_io_out_id_0),
		.io_out_last_0(_mesh_30_7_io_out_last_0),
		.io_out_valid_0(_mesh_30_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10338 == GlobalFiModInstNr[0]) || (10338 == GlobalFiModInstNr[1]) || (10338 == GlobalFiModInstNr[2]) || (10338 == GlobalFiModInstNr[3]))));
	Tile mesh_30_8(
		.clock(clock),
		.io_in_a_0(r_968_0),
		.io_in_b_0(b_286_0),
		.io_in_d_0(b_1310_0),
		.io_in_control_0_dataflow(mesh_30_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2334_0),
		.io_in_last_0(r_3358_0),
		.io_in_valid_0(r_1310_0),
		.io_out_a_0(_mesh_30_8_io_out_a_0),
		.io_out_c_0(_mesh_30_8_io_out_c_0),
		.io_out_b_0(_mesh_30_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_8_io_out_id_0),
		.io_out_last_0(_mesh_30_8_io_out_last_0),
		.io_out_valid_0(_mesh_30_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10339 == GlobalFiModInstNr[0]) || (10339 == GlobalFiModInstNr[1]) || (10339 == GlobalFiModInstNr[2]) || (10339 == GlobalFiModInstNr[3]))));
	Tile mesh_30_9(
		.clock(clock),
		.io_in_a_0(r_969_0),
		.io_in_b_0(b_318_0),
		.io_in_d_0(b_1342_0),
		.io_in_control_0_dataflow(mesh_30_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2366_0),
		.io_in_last_0(r_3390_0),
		.io_in_valid_0(r_1342_0),
		.io_out_a_0(_mesh_30_9_io_out_a_0),
		.io_out_c_0(_mesh_30_9_io_out_c_0),
		.io_out_b_0(_mesh_30_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_9_io_out_id_0),
		.io_out_last_0(_mesh_30_9_io_out_last_0),
		.io_out_valid_0(_mesh_30_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10340 == GlobalFiModInstNr[0]) || (10340 == GlobalFiModInstNr[1]) || (10340 == GlobalFiModInstNr[2]) || (10340 == GlobalFiModInstNr[3]))));
	Tile mesh_30_10(
		.clock(clock),
		.io_in_a_0(r_970_0),
		.io_in_b_0(b_350_0),
		.io_in_d_0(b_1374_0),
		.io_in_control_0_dataflow(mesh_30_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2398_0),
		.io_in_last_0(r_3422_0),
		.io_in_valid_0(r_1374_0),
		.io_out_a_0(_mesh_30_10_io_out_a_0),
		.io_out_c_0(_mesh_30_10_io_out_c_0),
		.io_out_b_0(_mesh_30_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_10_io_out_id_0),
		.io_out_last_0(_mesh_30_10_io_out_last_0),
		.io_out_valid_0(_mesh_30_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10341 == GlobalFiModInstNr[0]) || (10341 == GlobalFiModInstNr[1]) || (10341 == GlobalFiModInstNr[2]) || (10341 == GlobalFiModInstNr[3]))));
	Tile mesh_30_11(
		.clock(clock),
		.io_in_a_0(r_971_0),
		.io_in_b_0(b_382_0),
		.io_in_d_0(b_1406_0),
		.io_in_control_0_dataflow(mesh_30_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2430_0),
		.io_in_last_0(r_3454_0),
		.io_in_valid_0(r_1406_0),
		.io_out_a_0(_mesh_30_11_io_out_a_0),
		.io_out_c_0(_mesh_30_11_io_out_c_0),
		.io_out_b_0(_mesh_30_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_11_io_out_id_0),
		.io_out_last_0(_mesh_30_11_io_out_last_0),
		.io_out_valid_0(_mesh_30_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10342 == GlobalFiModInstNr[0]) || (10342 == GlobalFiModInstNr[1]) || (10342 == GlobalFiModInstNr[2]) || (10342 == GlobalFiModInstNr[3]))));
	Tile mesh_30_12(
		.clock(clock),
		.io_in_a_0(r_972_0),
		.io_in_b_0(b_414_0),
		.io_in_d_0(b_1438_0),
		.io_in_control_0_dataflow(mesh_30_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2462_0),
		.io_in_last_0(r_3486_0),
		.io_in_valid_0(r_1438_0),
		.io_out_a_0(_mesh_30_12_io_out_a_0),
		.io_out_c_0(_mesh_30_12_io_out_c_0),
		.io_out_b_0(_mesh_30_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_12_io_out_id_0),
		.io_out_last_0(_mesh_30_12_io_out_last_0),
		.io_out_valid_0(_mesh_30_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10343 == GlobalFiModInstNr[0]) || (10343 == GlobalFiModInstNr[1]) || (10343 == GlobalFiModInstNr[2]) || (10343 == GlobalFiModInstNr[3]))));
	Tile mesh_30_13(
		.clock(clock),
		.io_in_a_0(r_973_0),
		.io_in_b_0(b_446_0),
		.io_in_d_0(b_1470_0),
		.io_in_control_0_dataflow(mesh_30_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2494_0),
		.io_in_last_0(r_3518_0),
		.io_in_valid_0(r_1470_0),
		.io_out_a_0(_mesh_30_13_io_out_a_0),
		.io_out_c_0(_mesh_30_13_io_out_c_0),
		.io_out_b_0(_mesh_30_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_13_io_out_id_0),
		.io_out_last_0(_mesh_30_13_io_out_last_0),
		.io_out_valid_0(_mesh_30_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10344 == GlobalFiModInstNr[0]) || (10344 == GlobalFiModInstNr[1]) || (10344 == GlobalFiModInstNr[2]) || (10344 == GlobalFiModInstNr[3]))));
	Tile mesh_30_14(
		.clock(clock),
		.io_in_a_0(r_974_0),
		.io_in_b_0(b_478_0),
		.io_in_d_0(b_1502_0),
		.io_in_control_0_dataflow(mesh_30_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2526_0),
		.io_in_last_0(r_3550_0),
		.io_in_valid_0(r_1502_0),
		.io_out_a_0(_mesh_30_14_io_out_a_0),
		.io_out_c_0(_mesh_30_14_io_out_c_0),
		.io_out_b_0(_mesh_30_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_14_io_out_id_0),
		.io_out_last_0(_mesh_30_14_io_out_last_0),
		.io_out_valid_0(_mesh_30_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10345 == GlobalFiModInstNr[0]) || (10345 == GlobalFiModInstNr[1]) || (10345 == GlobalFiModInstNr[2]) || (10345 == GlobalFiModInstNr[3]))));
	Tile mesh_30_15(
		.clock(clock),
		.io_in_a_0(r_975_0),
		.io_in_b_0(b_510_0),
		.io_in_d_0(b_1534_0),
		.io_in_control_0_dataflow(mesh_30_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2558_0),
		.io_in_last_0(r_3582_0),
		.io_in_valid_0(r_1534_0),
		.io_out_a_0(_mesh_30_15_io_out_a_0),
		.io_out_c_0(_mesh_30_15_io_out_c_0),
		.io_out_b_0(_mesh_30_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_15_io_out_id_0),
		.io_out_last_0(_mesh_30_15_io_out_last_0),
		.io_out_valid_0(_mesh_30_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10346 == GlobalFiModInstNr[0]) || (10346 == GlobalFiModInstNr[1]) || (10346 == GlobalFiModInstNr[2]) || (10346 == GlobalFiModInstNr[3]))));
	Tile mesh_30_16(
		.clock(clock),
		.io_in_a_0(r_976_0),
		.io_in_b_0(b_542_0),
		.io_in_d_0(b_1566_0),
		.io_in_control_0_dataflow(mesh_30_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2590_0),
		.io_in_last_0(r_3614_0),
		.io_in_valid_0(r_1566_0),
		.io_out_a_0(_mesh_30_16_io_out_a_0),
		.io_out_c_0(_mesh_30_16_io_out_c_0),
		.io_out_b_0(_mesh_30_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_16_io_out_id_0),
		.io_out_last_0(_mesh_30_16_io_out_last_0),
		.io_out_valid_0(_mesh_30_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10347 == GlobalFiModInstNr[0]) || (10347 == GlobalFiModInstNr[1]) || (10347 == GlobalFiModInstNr[2]) || (10347 == GlobalFiModInstNr[3]))));
	Tile mesh_30_17(
		.clock(clock),
		.io_in_a_0(r_977_0),
		.io_in_b_0(b_574_0),
		.io_in_d_0(b_1598_0),
		.io_in_control_0_dataflow(mesh_30_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2622_0),
		.io_in_last_0(r_3646_0),
		.io_in_valid_0(r_1598_0),
		.io_out_a_0(_mesh_30_17_io_out_a_0),
		.io_out_c_0(_mesh_30_17_io_out_c_0),
		.io_out_b_0(_mesh_30_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_17_io_out_id_0),
		.io_out_last_0(_mesh_30_17_io_out_last_0),
		.io_out_valid_0(_mesh_30_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10348 == GlobalFiModInstNr[0]) || (10348 == GlobalFiModInstNr[1]) || (10348 == GlobalFiModInstNr[2]) || (10348 == GlobalFiModInstNr[3]))));
	Tile mesh_30_18(
		.clock(clock),
		.io_in_a_0(r_978_0),
		.io_in_b_0(b_606_0),
		.io_in_d_0(b_1630_0),
		.io_in_control_0_dataflow(mesh_30_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2654_0),
		.io_in_last_0(r_3678_0),
		.io_in_valid_0(r_1630_0),
		.io_out_a_0(_mesh_30_18_io_out_a_0),
		.io_out_c_0(_mesh_30_18_io_out_c_0),
		.io_out_b_0(_mesh_30_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_18_io_out_id_0),
		.io_out_last_0(_mesh_30_18_io_out_last_0),
		.io_out_valid_0(_mesh_30_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10349 == GlobalFiModInstNr[0]) || (10349 == GlobalFiModInstNr[1]) || (10349 == GlobalFiModInstNr[2]) || (10349 == GlobalFiModInstNr[3]))));
	Tile mesh_30_19(
		.clock(clock),
		.io_in_a_0(r_979_0),
		.io_in_b_0(b_638_0),
		.io_in_d_0(b_1662_0),
		.io_in_control_0_dataflow(mesh_30_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2686_0),
		.io_in_last_0(r_3710_0),
		.io_in_valid_0(r_1662_0),
		.io_out_a_0(_mesh_30_19_io_out_a_0),
		.io_out_c_0(_mesh_30_19_io_out_c_0),
		.io_out_b_0(_mesh_30_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_19_io_out_id_0),
		.io_out_last_0(_mesh_30_19_io_out_last_0),
		.io_out_valid_0(_mesh_30_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10350 == GlobalFiModInstNr[0]) || (10350 == GlobalFiModInstNr[1]) || (10350 == GlobalFiModInstNr[2]) || (10350 == GlobalFiModInstNr[3]))));
	Tile mesh_30_20(
		.clock(clock),
		.io_in_a_0(r_980_0),
		.io_in_b_0(b_670_0),
		.io_in_d_0(b_1694_0),
		.io_in_control_0_dataflow(mesh_30_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2718_0),
		.io_in_last_0(r_3742_0),
		.io_in_valid_0(r_1694_0),
		.io_out_a_0(_mesh_30_20_io_out_a_0),
		.io_out_c_0(_mesh_30_20_io_out_c_0),
		.io_out_b_0(_mesh_30_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_20_io_out_id_0),
		.io_out_last_0(_mesh_30_20_io_out_last_0),
		.io_out_valid_0(_mesh_30_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10351 == GlobalFiModInstNr[0]) || (10351 == GlobalFiModInstNr[1]) || (10351 == GlobalFiModInstNr[2]) || (10351 == GlobalFiModInstNr[3]))));
	Tile mesh_30_21(
		.clock(clock),
		.io_in_a_0(r_981_0),
		.io_in_b_0(b_702_0),
		.io_in_d_0(b_1726_0),
		.io_in_control_0_dataflow(mesh_30_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2750_0),
		.io_in_last_0(r_3774_0),
		.io_in_valid_0(r_1726_0),
		.io_out_a_0(_mesh_30_21_io_out_a_0),
		.io_out_c_0(_mesh_30_21_io_out_c_0),
		.io_out_b_0(_mesh_30_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_21_io_out_id_0),
		.io_out_last_0(_mesh_30_21_io_out_last_0),
		.io_out_valid_0(_mesh_30_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10352 == GlobalFiModInstNr[0]) || (10352 == GlobalFiModInstNr[1]) || (10352 == GlobalFiModInstNr[2]) || (10352 == GlobalFiModInstNr[3]))));
	Tile mesh_30_22(
		.clock(clock),
		.io_in_a_0(r_982_0),
		.io_in_b_0(b_734_0),
		.io_in_d_0(b_1758_0),
		.io_in_control_0_dataflow(mesh_30_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2782_0),
		.io_in_last_0(r_3806_0),
		.io_in_valid_0(r_1758_0),
		.io_out_a_0(_mesh_30_22_io_out_a_0),
		.io_out_c_0(_mesh_30_22_io_out_c_0),
		.io_out_b_0(_mesh_30_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_22_io_out_id_0),
		.io_out_last_0(_mesh_30_22_io_out_last_0),
		.io_out_valid_0(_mesh_30_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10353 == GlobalFiModInstNr[0]) || (10353 == GlobalFiModInstNr[1]) || (10353 == GlobalFiModInstNr[2]) || (10353 == GlobalFiModInstNr[3]))));
	Tile mesh_30_23(
		.clock(clock),
		.io_in_a_0(r_983_0),
		.io_in_b_0(b_766_0),
		.io_in_d_0(b_1790_0),
		.io_in_control_0_dataflow(mesh_30_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2814_0),
		.io_in_last_0(r_3838_0),
		.io_in_valid_0(r_1790_0),
		.io_out_a_0(_mesh_30_23_io_out_a_0),
		.io_out_c_0(_mesh_30_23_io_out_c_0),
		.io_out_b_0(_mesh_30_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_23_io_out_id_0),
		.io_out_last_0(_mesh_30_23_io_out_last_0),
		.io_out_valid_0(_mesh_30_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10354 == GlobalFiModInstNr[0]) || (10354 == GlobalFiModInstNr[1]) || (10354 == GlobalFiModInstNr[2]) || (10354 == GlobalFiModInstNr[3]))));
	Tile mesh_30_24(
		.clock(clock),
		.io_in_a_0(r_984_0),
		.io_in_b_0(b_798_0),
		.io_in_d_0(b_1822_0),
		.io_in_control_0_dataflow(mesh_30_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2846_0),
		.io_in_last_0(r_3870_0),
		.io_in_valid_0(r_1822_0),
		.io_out_a_0(_mesh_30_24_io_out_a_0),
		.io_out_c_0(_mesh_30_24_io_out_c_0),
		.io_out_b_0(_mesh_30_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_24_io_out_id_0),
		.io_out_last_0(_mesh_30_24_io_out_last_0),
		.io_out_valid_0(_mesh_30_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10355 == GlobalFiModInstNr[0]) || (10355 == GlobalFiModInstNr[1]) || (10355 == GlobalFiModInstNr[2]) || (10355 == GlobalFiModInstNr[3]))));
	Tile mesh_30_25(
		.clock(clock),
		.io_in_a_0(r_985_0),
		.io_in_b_0(b_830_0),
		.io_in_d_0(b_1854_0),
		.io_in_control_0_dataflow(mesh_30_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2878_0),
		.io_in_last_0(r_3902_0),
		.io_in_valid_0(r_1854_0),
		.io_out_a_0(_mesh_30_25_io_out_a_0),
		.io_out_c_0(_mesh_30_25_io_out_c_0),
		.io_out_b_0(_mesh_30_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_25_io_out_id_0),
		.io_out_last_0(_mesh_30_25_io_out_last_0),
		.io_out_valid_0(_mesh_30_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10356 == GlobalFiModInstNr[0]) || (10356 == GlobalFiModInstNr[1]) || (10356 == GlobalFiModInstNr[2]) || (10356 == GlobalFiModInstNr[3]))));
	Tile mesh_30_26(
		.clock(clock),
		.io_in_a_0(r_986_0),
		.io_in_b_0(b_862_0),
		.io_in_d_0(b_1886_0),
		.io_in_control_0_dataflow(mesh_30_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2910_0),
		.io_in_last_0(r_3934_0),
		.io_in_valid_0(r_1886_0),
		.io_out_a_0(_mesh_30_26_io_out_a_0),
		.io_out_c_0(_mesh_30_26_io_out_c_0),
		.io_out_b_0(_mesh_30_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_26_io_out_id_0),
		.io_out_last_0(_mesh_30_26_io_out_last_0),
		.io_out_valid_0(_mesh_30_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10357 == GlobalFiModInstNr[0]) || (10357 == GlobalFiModInstNr[1]) || (10357 == GlobalFiModInstNr[2]) || (10357 == GlobalFiModInstNr[3]))));
	Tile mesh_30_27(
		.clock(clock),
		.io_in_a_0(r_987_0),
		.io_in_b_0(b_894_0),
		.io_in_d_0(b_1918_0),
		.io_in_control_0_dataflow(mesh_30_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2942_0),
		.io_in_last_0(r_3966_0),
		.io_in_valid_0(r_1918_0),
		.io_out_a_0(_mesh_30_27_io_out_a_0),
		.io_out_c_0(_mesh_30_27_io_out_c_0),
		.io_out_b_0(_mesh_30_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_27_io_out_id_0),
		.io_out_last_0(_mesh_30_27_io_out_last_0),
		.io_out_valid_0(_mesh_30_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10358 == GlobalFiModInstNr[0]) || (10358 == GlobalFiModInstNr[1]) || (10358 == GlobalFiModInstNr[2]) || (10358 == GlobalFiModInstNr[3]))));
	Tile mesh_30_28(
		.clock(clock),
		.io_in_a_0(r_988_0),
		.io_in_b_0(b_926_0),
		.io_in_d_0(b_1950_0),
		.io_in_control_0_dataflow(mesh_30_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2974_0),
		.io_in_last_0(r_3998_0),
		.io_in_valid_0(r_1950_0),
		.io_out_a_0(_mesh_30_28_io_out_a_0),
		.io_out_c_0(_mesh_30_28_io_out_c_0),
		.io_out_b_0(_mesh_30_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_28_io_out_id_0),
		.io_out_last_0(_mesh_30_28_io_out_last_0),
		.io_out_valid_0(_mesh_30_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10359 == GlobalFiModInstNr[0]) || (10359 == GlobalFiModInstNr[1]) || (10359 == GlobalFiModInstNr[2]) || (10359 == GlobalFiModInstNr[3]))));
	Tile mesh_30_29(
		.clock(clock),
		.io_in_a_0(r_989_0),
		.io_in_b_0(b_958_0),
		.io_in_d_0(b_1982_0),
		.io_in_control_0_dataflow(mesh_30_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3006_0),
		.io_in_last_0(r_4030_0),
		.io_in_valid_0(r_1982_0),
		.io_out_a_0(_mesh_30_29_io_out_a_0),
		.io_out_c_0(_mesh_30_29_io_out_c_0),
		.io_out_b_0(_mesh_30_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_29_io_out_id_0),
		.io_out_last_0(_mesh_30_29_io_out_last_0),
		.io_out_valid_0(_mesh_30_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10360 == GlobalFiModInstNr[0]) || (10360 == GlobalFiModInstNr[1]) || (10360 == GlobalFiModInstNr[2]) || (10360 == GlobalFiModInstNr[3]))));
	Tile mesh_30_30(
		.clock(clock),
		.io_in_a_0(r_990_0),
		.io_in_b_0(b_990_0),
		.io_in_d_0(b_2014_0),
		.io_in_control_0_dataflow(mesh_30_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3038_0),
		.io_in_last_0(r_4062_0),
		.io_in_valid_0(r_2014_0),
		.io_out_a_0(_mesh_30_30_io_out_a_0),
		.io_out_c_0(_mesh_30_30_io_out_c_0),
		.io_out_b_0(_mesh_30_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_30_io_out_id_0),
		.io_out_last_0(_mesh_30_30_io_out_last_0),
		.io_out_valid_0(_mesh_30_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10361 == GlobalFiModInstNr[0]) || (10361 == GlobalFiModInstNr[1]) || (10361 == GlobalFiModInstNr[2]) || (10361 == GlobalFiModInstNr[3]))));
	Tile mesh_30_31(
		.clock(clock),
		.io_in_a_0(r_991_0),
		.io_in_b_0(b_1022_0),
		.io_in_d_0(b_2046_0),
		.io_in_control_0_dataflow(mesh_30_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_30_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_30_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3070_0),
		.io_in_last_0(r_4094_0),
		.io_in_valid_0(r_2046_0),
		.io_out_a_0(_mesh_30_31_io_out_a_0),
		.io_out_c_0(_mesh_30_31_io_out_c_0),
		.io_out_b_0(_mesh_30_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_30_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_30_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_30_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_30_31_io_out_id_0),
		.io_out_last_0(_mesh_30_31_io_out_last_0),
		.io_out_valid_0(_mesh_30_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10362 == GlobalFiModInstNr[0]) || (10362 == GlobalFiModInstNr[1]) || (10362 == GlobalFiModInstNr[2]) || (10362 == GlobalFiModInstNr[3]))));
	Tile mesh_31_0(
		.clock(clock),
		.io_in_a_0(r_992_0),
		.io_in_b_0(b_31_0),
		.io_in_d_0(b_1055_0),
		.io_in_control_0_dataflow(mesh_31_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_0_io_in_control_0_shift_b),
		.io_in_id_0(r_2079_0),
		.io_in_last_0(r_3103_0),
		.io_in_valid_0(r_1055_0),
		.io_out_a_0(_mesh_31_0_io_out_a_0),
		.io_out_c_0(_mesh_31_0_io_out_c_0),
		.io_out_b_0(_mesh_31_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_0_io_out_id_0),
		.io_out_last_0(_mesh_31_0_io_out_last_0),
		.io_out_valid_0(_mesh_31_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10363 == GlobalFiModInstNr[0]) || (10363 == GlobalFiModInstNr[1]) || (10363 == GlobalFiModInstNr[2]) || (10363 == GlobalFiModInstNr[3]))));
	Tile mesh_31_1(
		.clock(clock),
		.io_in_a_0(r_993_0),
		.io_in_b_0(b_63_0),
		.io_in_d_0(b_1087_0),
		.io_in_control_0_dataflow(mesh_31_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_1_io_in_control_0_shift_b),
		.io_in_id_0(r_2111_0),
		.io_in_last_0(r_3135_0),
		.io_in_valid_0(r_1087_0),
		.io_out_a_0(_mesh_31_1_io_out_a_0),
		.io_out_c_0(_mesh_31_1_io_out_c_0),
		.io_out_b_0(_mesh_31_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_1_io_out_id_0),
		.io_out_last_0(_mesh_31_1_io_out_last_0),
		.io_out_valid_0(_mesh_31_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10364 == GlobalFiModInstNr[0]) || (10364 == GlobalFiModInstNr[1]) || (10364 == GlobalFiModInstNr[2]) || (10364 == GlobalFiModInstNr[3]))));
	Tile mesh_31_2(
		.clock(clock),
		.io_in_a_0(r_994_0),
		.io_in_b_0(b_95_0),
		.io_in_d_0(b_1119_0),
		.io_in_control_0_dataflow(mesh_31_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_2_io_in_control_0_shift_b),
		.io_in_id_0(r_2143_0),
		.io_in_last_0(r_3167_0),
		.io_in_valid_0(r_1119_0),
		.io_out_a_0(_mesh_31_2_io_out_a_0),
		.io_out_c_0(_mesh_31_2_io_out_c_0),
		.io_out_b_0(_mesh_31_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_2_io_out_id_0),
		.io_out_last_0(_mesh_31_2_io_out_last_0),
		.io_out_valid_0(_mesh_31_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10365 == GlobalFiModInstNr[0]) || (10365 == GlobalFiModInstNr[1]) || (10365 == GlobalFiModInstNr[2]) || (10365 == GlobalFiModInstNr[3]))));
	Tile mesh_31_3(
		.clock(clock),
		.io_in_a_0(r_995_0),
		.io_in_b_0(b_127_0),
		.io_in_d_0(b_1151_0),
		.io_in_control_0_dataflow(mesh_31_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_3_io_in_control_0_shift_b),
		.io_in_id_0(r_2175_0),
		.io_in_last_0(r_3199_0),
		.io_in_valid_0(r_1151_0),
		.io_out_a_0(_mesh_31_3_io_out_a_0),
		.io_out_c_0(_mesh_31_3_io_out_c_0),
		.io_out_b_0(_mesh_31_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_3_io_out_id_0),
		.io_out_last_0(_mesh_31_3_io_out_last_0),
		.io_out_valid_0(_mesh_31_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10366 == GlobalFiModInstNr[0]) || (10366 == GlobalFiModInstNr[1]) || (10366 == GlobalFiModInstNr[2]) || (10366 == GlobalFiModInstNr[3]))));
	Tile mesh_31_4(
		.clock(clock),
		.io_in_a_0(r_996_0),
		.io_in_b_0(b_159_0),
		.io_in_d_0(b_1183_0),
		.io_in_control_0_dataflow(mesh_31_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_4_io_in_control_0_shift_b),
		.io_in_id_0(r_2207_0),
		.io_in_last_0(r_3231_0),
		.io_in_valid_0(r_1183_0),
		.io_out_a_0(_mesh_31_4_io_out_a_0),
		.io_out_c_0(_mesh_31_4_io_out_c_0),
		.io_out_b_0(_mesh_31_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_4_io_out_id_0),
		.io_out_last_0(_mesh_31_4_io_out_last_0),
		.io_out_valid_0(_mesh_31_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10367 == GlobalFiModInstNr[0]) || (10367 == GlobalFiModInstNr[1]) || (10367 == GlobalFiModInstNr[2]) || (10367 == GlobalFiModInstNr[3]))));
	Tile mesh_31_5(
		.clock(clock),
		.io_in_a_0(r_997_0),
		.io_in_b_0(b_191_0),
		.io_in_d_0(b_1215_0),
		.io_in_control_0_dataflow(mesh_31_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_5_io_in_control_0_shift_b),
		.io_in_id_0(r_2239_0),
		.io_in_last_0(r_3263_0),
		.io_in_valid_0(r_1215_0),
		.io_out_a_0(_mesh_31_5_io_out_a_0),
		.io_out_c_0(_mesh_31_5_io_out_c_0),
		.io_out_b_0(_mesh_31_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_5_io_out_id_0),
		.io_out_last_0(_mesh_31_5_io_out_last_0),
		.io_out_valid_0(_mesh_31_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10368 == GlobalFiModInstNr[0]) || (10368 == GlobalFiModInstNr[1]) || (10368 == GlobalFiModInstNr[2]) || (10368 == GlobalFiModInstNr[3]))));
	Tile mesh_31_6(
		.clock(clock),
		.io_in_a_0(r_998_0),
		.io_in_b_0(b_223_0),
		.io_in_d_0(b_1247_0),
		.io_in_control_0_dataflow(mesh_31_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_6_io_in_control_0_shift_b),
		.io_in_id_0(r_2271_0),
		.io_in_last_0(r_3295_0),
		.io_in_valid_0(r_1247_0),
		.io_out_a_0(_mesh_31_6_io_out_a_0),
		.io_out_c_0(_mesh_31_6_io_out_c_0),
		.io_out_b_0(_mesh_31_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_6_io_out_id_0),
		.io_out_last_0(_mesh_31_6_io_out_last_0),
		.io_out_valid_0(_mesh_31_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10369 == GlobalFiModInstNr[0]) || (10369 == GlobalFiModInstNr[1]) || (10369 == GlobalFiModInstNr[2]) || (10369 == GlobalFiModInstNr[3]))));
	Tile mesh_31_7(
		.clock(clock),
		.io_in_a_0(r_999_0),
		.io_in_b_0(b_255_0),
		.io_in_d_0(b_1279_0),
		.io_in_control_0_dataflow(mesh_31_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_7_io_in_control_0_shift_b),
		.io_in_id_0(r_2303_0),
		.io_in_last_0(r_3327_0),
		.io_in_valid_0(r_1279_0),
		.io_out_a_0(_mesh_31_7_io_out_a_0),
		.io_out_c_0(_mesh_31_7_io_out_c_0),
		.io_out_b_0(_mesh_31_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_7_io_out_id_0),
		.io_out_last_0(_mesh_31_7_io_out_last_0),
		.io_out_valid_0(_mesh_31_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10370 == GlobalFiModInstNr[0]) || (10370 == GlobalFiModInstNr[1]) || (10370 == GlobalFiModInstNr[2]) || (10370 == GlobalFiModInstNr[3]))));
	Tile mesh_31_8(
		.clock(clock),
		.io_in_a_0(r_1000_0),
		.io_in_b_0(b_287_0),
		.io_in_d_0(b_1311_0),
		.io_in_control_0_dataflow(mesh_31_8_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_8_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_8_io_in_control_0_shift_b),
		.io_in_id_0(r_2335_0),
		.io_in_last_0(r_3359_0),
		.io_in_valid_0(r_1311_0),
		.io_out_a_0(_mesh_31_8_io_out_a_0),
		.io_out_c_0(_mesh_31_8_io_out_c_0),
		.io_out_b_0(_mesh_31_8_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_8_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_8_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_8_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_8_io_out_id_0),
		.io_out_last_0(_mesh_31_8_io_out_last_0),
		.io_out_valid_0(_mesh_31_8_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10371 == GlobalFiModInstNr[0]) || (10371 == GlobalFiModInstNr[1]) || (10371 == GlobalFiModInstNr[2]) || (10371 == GlobalFiModInstNr[3]))));
	Tile mesh_31_9(
		.clock(clock),
		.io_in_a_0(r_1001_0),
		.io_in_b_0(b_319_0),
		.io_in_d_0(b_1343_0),
		.io_in_control_0_dataflow(mesh_31_9_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_9_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_9_io_in_control_0_shift_b),
		.io_in_id_0(r_2367_0),
		.io_in_last_0(r_3391_0),
		.io_in_valid_0(r_1343_0),
		.io_out_a_0(_mesh_31_9_io_out_a_0),
		.io_out_c_0(_mesh_31_9_io_out_c_0),
		.io_out_b_0(_mesh_31_9_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_9_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_9_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_9_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_9_io_out_id_0),
		.io_out_last_0(_mesh_31_9_io_out_last_0),
		.io_out_valid_0(_mesh_31_9_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10372 == GlobalFiModInstNr[0]) || (10372 == GlobalFiModInstNr[1]) || (10372 == GlobalFiModInstNr[2]) || (10372 == GlobalFiModInstNr[3]))));
	Tile mesh_31_10(
		.clock(clock),
		.io_in_a_0(r_1002_0),
		.io_in_b_0(b_351_0),
		.io_in_d_0(b_1375_0),
		.io_in_control_0_dataflow(mesh_31_10_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_10_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_10_io_in_control_0_shift_b),
		.io_in_id_0(r_2399_0),
		.io_in_last_0(r_3423_0),
		.io_in_valid_0(r_1375_0),
		.io_out_a_0(_mesh_31_10_io_out_a_0),
		.io_out_c_0(_mesh_31_10_io_out_c_0),
		.io_out_b_0(_mesh_31_10_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_10_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_10_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_10_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_10_io_out_id_0),
		.io_out_last_0(_mesh_31_10_io_out_last_0),
		.io_out_valid_0(_mesh_31_10_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10373 == GlobalFiModInstNr[0]) || (10373 == GlobalFiModInstNr[1]) || (10373 == GlobalFiModInstNr[2]) || (10373 == GlobalFiModInstNr[3]))));
	Tile mesh_31_11(
		.clock(clock),
		.io_in_a_0(r_1003_0),
		.io_in_b_0(b_383_0),
		.io_in_d_0(b_1407_0),
		.io_in_control_0_dataflow(mesh_31_11_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_11_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_11_io_in_control_0_shift_b),
		.io_in_id_0(r_2431_0),
		.io_in_last_0(r_3455_0),
		.io_in_valid_0(r_1407_0),
		.io_out_a_0(_mesh_31_11_io_out_a_0),
		.io_out_c_0(_mesh_31_11_io_out_c_0),
		.io_out_b_0(_mesh_31_11_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_11_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_11_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_11_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_11_io_out_id_0),
		.io_out_last_0(_mesh_31_11_io_out_last_0),
		.io_out_valid_0(_mesh_31_11_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10374 == GlobalFiModInstNr[0]) || (10374 == GlobalFiModInstNr[1]) || (10374 == GlobalFiModInstNr[2]) || (10374 == GlobalFiModInstNr[3]))));
	Tile mesh_31_12(
		.clock(clock),
		.io_in_a_0(r_1004_0),
		.io_in_b_0(b_415_0),
		.io_in_d_0(b_1439_0),
		.io_in_control_0_dataflow(mesh_31_12_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_12_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_12_io_in_control_0_shift_b),
		.io_in_id_0(r_2463_0),
		.io_in_last_0(r_3487_0),
		.io_in_valid_0(r_1439_0),
		.io_out_a_0(_mesh_31_12_io_out_a_0),
		.io_out_c_0(_mesh_31_12_io_out_c_0),
		.io_out_b_0(_mesh_31_12_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_12_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_12_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_12_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_12_io_out_id_0),
		.io_out_last_0(_mesh_31_12_io_out_last_0),
		.io_out_valid_0(_mesh_31_12_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10375 == GlobalFiModInstNr[0]) || (10375 == GlobalFiModInstNr[1]) || (10375 == GlobalFiModInstNr[2]) || (10375 == GlobalFiModInstNr[3]))));
	Tile mesh_31_13(
		.clock(clock),
		.io_in_a_0(r_1005_0),
		.io_in_b_0(b_447_0),
		.io_in_d_0(b_1471_0),
		.io_in_control_0_dataflow(mesh_31_13_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_13_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_13_io_in_control_0_shift_b),
		.io_in_id_0(r_2495_0),
		.io_in_last_0(r_3519_0),
		.io_in_valid_0(r_1471_0),
		.io_out_a_0(_mesh_31_13_io_out_a_0),
		.io_out_c_0(_mesh_31_13_io_out_c_0),
		.io_out_b_0(_mesh_31_13_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_13_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_13_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_13_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_13_io_out_id_0),
		.io_out_last_0(_mesh_31_13_io_out_last_0),
		.io_out_valid_0(_mesh_31_13_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10376 == GlobalFiModInstNr[0]) || (10376 == GlobalFiModInstNr[1]) || (10376 == GlobalFiModInstNr[2]) || (10376 == GlobalFiModInstNr[3]))));
	Tile mesh_31_14(
		.clock(clock),
		.io_in_a_0(r_1006_0),
		.io_in_b_0(b_479_0),
		.io_in_d_0(b_1503_0),
		.io_in_control_0_dataflow(mesh_31_14_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_14_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_14_io_in_control_0_shift_b),
		.io_in_id_0(r_2527_0),
		.io_in_last_0(r_3551_0),
		.io_in_valid_0(r_1503_0),
		.io_out_a_0(_mesh_31_14_io_out_a_0),
		.io_out_c_0(_mesh_31_14_io_out_c_0),
		.io_out_b_0(_mesh_31_14_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_14_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_14_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_14_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_14_io_out_id_0),
		.io_out_last_0(_mesh_31_14_io_out_last_0),
		.io_out_valid_0(_mesh_31_14_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10377 == GlobalFiModInstNr[0]) || (10377 == GlobalFiModInstNr[1]) || (10377 == GlobalFiModInstNr[2]) || (10377 == GlobalFiModInstNr[3]))));
	Tile mesh_31_15(
		.clock(clock),
		.io_in_a_0(r_1007_0),
		.io_in_b_0(b_511_0),
		.io_in_d_0(b_1535_0),
		.io_in_control_0_dataflow(mesh_31_15_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_15_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_15_io_in_control_0_shift_b),
		.io_in_id_0(r_2559_0),
		.io_in_last_0(r_3583_0),
		.io_in_valid_0(r_1535_0),
		.io_out_a_0(_mesh_31_15_io_out_a_0),
		.io_out_c_0(_mesh_31_15_io_out_c_0),
		.io_out_b_0(_mesh_31_15_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_15_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_15_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_15_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_15_io_out_id_0),
		.io_out_last_0(_mesh_31_15_io_out_last_0),
		.io_out_valid_0(_mesh_31_15_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10378 == GlobalFiModInstNr[0]) || (10378 == GlobalFiModInstNr[1]) || (10378 == GlobalFiModInstNr[2]) || (10378 == GlobalFiModInstNr[3]))));
	Tile mesh_31_16(
		.clock(clock),
		.io_in_a_0(r_1008_0),
		.io_in_b_0(b_543_0),
		.io_in_d_0(b_1567_0),
		.io_in_control_0_dataflow(mesh_31_16_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_16_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_16_io_in_control_0_shift_b),
		.io_in_id_0(r_2591_0),
		.io_in_last_0(r_3615_0),
		.io_in_valid_0(r_1567_0),
		.io_out_a_0(_mesh_31_16_io_out_a_0),
		.io_out_c_0(_mesh_31_16_io_out_c_0),
		.io_out_b_0(_mesh_31_16_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_16_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_16_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_16_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_16_io_out_id_0),
		.io_out_last_0(_mesh_31_16_io_out_last_0),
		.io_out_valid_0(_mesh_31_16_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10379 == GlobalFiModInstNr[0]) || (10379 == GlobalFiModInstNr[1]) || (10379 == GlobalFiModInstNr[2]) || (10379 == GlobalFiModInstNr[3]))));
	Tile mesh_31_17(
		.clock(clock),
		.io_in_a_0(r_1009_0),
		.io_in_b_0(b_575_0),
		.io_in_d_0(b_1599_0),
		.io_in_control_0_dataflow(mesh_31_17_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_17_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_17_io_in_control_0_shift_b),
		.io_in_id_0(r_2623_0),
		.io_in_last_0(r_3647_0),
		.io_in_valid_0(r_1599_0),
		.io_out_a_0(_mesh_31_17_io_out_a_0),
		.io_out_c_0(_mesh_31_17_io_out_c_0),
		.io_out_b_0(_mesh_31_17_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_17_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_17_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_17_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_17_io_out_id_0),
		.io_out_last_0(_mesh_31_17_io_out_last_0),
		.io_out_valid_0(_mesh_31_17_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10380 == GlobalFiModInstNr[0]) || (10380 == GlobalFiModInstNr[1]) || (10380 == GlobalFiModInstNr[2]) || (10380 == GlobalFiModInstNr[3]))));
	Tile mesh_31_18(
		.clock(clock),
		.io_in_a_0(r_1010_0),
		.io_in_b_0(b_607_0),
		.io_in_d_0(b_1631_0),
		.io_in_control_0_dataflow(mesh_31_18_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_18_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_18_io_in_control_0_shift_b),
		.io_in_id_0(r_2655_0),
		.io_in_last_0(r_3679_0),
		.io_in_valid_0(r_1631_0),
		.io_out_a_0(_mesh_31_18_io_out_a_0),
		.io_out_c_0(_mesh_31_18_io_out_c_0),
		.io_out_b_0(_mesh_31_18_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_18_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_18_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_18_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_18_io_out_id_0),
		.io_out_last_0(_mesh_31_18_io_out_last_0),
		.io_out_valid_0(_mesh_31_18_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10381 == GlobalFiModInstNr[0]) || (10381 == GlobalFiModInstNr[1]) || (10381 == GlobalFiModInstNr[2]) || (10381 == GlobalFiModInstNr[3]))));
	Tile mesh_31_19(
		.clock(clock),
		.io_in_a_0(r_1011_0),
		.io_in_b_0(b_639_0),
		.io_in_d_0(b_1663_0),
		.io_in_control_0_dataflow(mesh_31_19_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_19_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_19_io_in_control_0_shift_b),
		.io_in_id_0(r_2687_0),
		.io_in_last_0(r_3711_0),
		.io_in_valid_0(r_1663_0),
		.io_out_a_0(_mesh_31_19_io_out_a_0),
		.io_out_c_0(_mesh_31_19_io_out_c_0),
		.io_out_b_0(_mesh_31_19_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_19_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_19_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_19_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_19_io_out_id_0),
		.io_out_last_0(_mesh_31_19_io_out_last_0),
		.io_out_valid_0(_mesh_31_19_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10382 == GlobalFiModInstNr[0]) || (10382 == GlobalFiModInstNr[1]) || (10382 == GlobalFiModInstNr[2]) || (10382 == GlobalFiModInstNr[3]))));
	Tile mesh_31_20(
		.clock(clock),
		.io_in_a_0(r_1012_0),
		.io_in_b_0(b_671_0),
		.io_in_d_0(b_1695_0),
		.io_in_control_0_dataflow(mesh_31_20_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_20_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_20_io_in_control_0_shift_b),
		.io_in_id_0(r_2719_0),
		.io_in_last_0(r_3743_0),
		.io_in_valid_0(r_1695_0),
		.io_out_a_0(_mesh_31_20_io_out_a_0),
		.io_out_c_0(_mesh_31_20_io_out_c_0),
		.io_out_b_0(_mesh_31_20_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_20_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_20_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_20_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_20_io_out_id_0),
		.io_out_last_0(_mesh_31_20_io_out_last_0),
		.io_out_valid_0(_mesh_31_20_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10383 == GlobalFiModInstNr[0]) || (10383 == GlobalFiModInstNr[1]) || (10383 == GlobalFiModInstNr[2]) || (10383 == GlobalFiModInstNr[3]))));
	Tile mesh_31_21(
		.clock(clock),
		.io_in_a_0(r_1013_0),
		.io_in_b_0(b_703_0),
		.io_in_d_0(b_1727_0),
		.io_in_control_0_dataflow(mesh_31_21_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_21_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_21_io_in_control_0_shift_b),
		.io_in_id_0(r_2751_0),
		.io_in_last_0(r_3775_0),
		.io_in_valid_0(r_1727_0),
		.io_out_a_0(_mesh_31_21_io_out_a_0),
		.io_out_c_0(_mesh_31_21_io_out_c_0),
		.io_out_b_0(_mesh_31_21_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_21_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_21_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_21_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_21_io_out_id_0),
		.io_out_last_0(_mesh_31_21_io_out_last_0),
		.io_out_valid_0(_mesh_31_21_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10384 == GlobalFiModInstNr[0]) || (10384 == GlobalFiModInstNr[1]) || (10384 == GlobalFiModInstNr[2]) || (10384 == GlobalFiModInstNr[3]))));
	Tile mesh_31_22(
		.clock(clock),
		.io_in_a_0(r_1014_0),
		.io_in_b_0(b_735_0),
		.io_in_d_0(b_1759_0),
		.io_in_control_0_dataflow(mesh_31_22_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_22_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_22_io_in_control_0_shift_b),
		.io_in_id_0(r_2783_0),
		.io_in_last_0(r_3807_0),
		.io_in_valid_0(r_1759_0),
		.io_out_a_0(_mesh_31_22_io_out_a_0),
		.io_out_c_0(_mesh_31_22_io_out_c_0),
		.io_out_b_0(_mesh_31_22_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_22_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_22_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_22_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_22_io_out_id_0),
		.io_out_last_0(_mesh_31_22_io_out_last_0),
		.io_out_valid_0(_mesh_31_22_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10385 == GlobalFiModInstNr[0]) || (10385 == GlobalFiModInstNr[1]) || (10385 == GlobalFiModInstNr[2]) || (10385 == GlobalFiModInstNr[3]))));
	Tile mesh_31_23(
		.clock(clock),
		.io_in_a_0(r_1015_0),
		.io_in_b_0(b_767_0),
		.io_in_d_0(b_1791_0),
		.io_in_control_0_dataflow(mesh_31_23_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_23_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_23_io_in_control_0_shift_b),
		.io_in_id_0(r_2815_0),
		.io_in_last_0(r_3839_0),
		.io_in_valid_0(r_1791_0),
		.io_out_a_0(_mesh_31_23_io_out_a_0),
		.io_out_c_0(_mesh_31_23_io_out_c_0),
		.io_out_b_0(_mesh_31_23_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_23_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_23_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_23_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_23_io_out_id_0),
		.io_out_last_0(_mesh_31_23_io_out_last_0),
		.io_out_valid_0(_mesh_31_23_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10386 == GlobalFiModInstNr[0]) || (10386 == GlobalFiModInstNr[1]) || (10386 == GlobalFiModInstNr[2]) || (10386 == GlobalFiModInstNr[3]))));
	Tile mesh_31_24(
		.clock(clock),
		.io_in_a_0(r_1016_0),
		.io_in_b_0(b_799_0),
		.io_in_d_0(b_1823_0),
		.io_in_control_0_dataflow(mesh_31_24_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_24_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_24_io_in_control_0_shift_b),
		.io_in_id_0(r_2847_0),
		.io_in_last_0(r_3871_0),
		.io_in_valid_0(r_1823_0),
		.io_out_a_0(_mesh_31_24_io_out_a_0),
		.io_out_c_0(_mesh_31_24_io_out_c_0),
		.io_out_b_0(_mesh_31_24_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_24_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_24_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_24_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_24_io_out_id_0),
		.io_out_last_0(_mesh_31_24_io_out_last_0),
		.io_out_valid_0(_mesh_31_24_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10387 == GlobalFiModInstNr[0]) || (10387 == GlobalFiModInstNr[1]) || (10387 == GlobalFiModInstNr[2]) || (10387 == GlobalFiModInstNr[3]))));
	Tile mesh_31_25(
		.clock(clock),
		.io_in_a_0(r_1017_0),
		.io_in_b_0(b_831_0),
		.io_in_d_0(b_1855_0),
		.io_in_control_0_dataflow(mesh_31_25_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_25_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_25_io_in_control_0_shift_b),
		.io_in_id_0(r_2879_0),
		.io_in_last_0(r_3903_0),
		.io_in_valid_0(r_1855_0),
		.io_out_a_0(_mesh_31_25_io_out_a_0),
		.io_out_c_0(_mesh_31_25_io_out_c_0),
		.io_out_b_0(_mesh_31_25_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_25_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_25_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_25_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_25_io_out_id_0),
		.io_out_last_0(_mesh_31_25_io_out_last_0),
		.io_out_valid_0(_mesh_31_25_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10388 == GlobalFiModInstNr[0]) || (10388 == GlobalFiModInstNr[1]) || (10388 == GlobalFiModInstNr[2]) || (10388 == GlobalFiModInstNr[3]))));
	Tile mesh_31_26(
		.clock(clock),
		.io_in_a_0(r_1018_0),
		.io_in_b_0(b_863_0),
		.io_in_d_0(b_1887_0),
		.io_in_control_0_dataflow(mesh_31_26_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_26_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_26_io_in_control_0_shift_b),
		.io_in_id_0(r_2911_0),
		.io_in_last_0(r_3935_0),
		.io_in_valid_0(r_1887_0),
		.io_out_a_0(_mesh_31_26_io_out_a_0),
		.io_out_c_0(_mesh_31_26_io_out_c_0),
		.io_out_b_0(_mesh_31_26_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_26_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_26_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_26_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_26_io_out_id_0),
		.io_out_last_0(_mesh_31_26_io_out_last_0),
		.io_out_valid_0(_mesh_31_26_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10389 == GlobalFiModInstNr[0]) || (10389 == GlobalFiModInstNr[1]) || (10389 == GlobalFiModInstNr[2]) || (10389 == GlobalFiModInstNr[3]))));
	Tile mesh_31_27(
		.clock(clock),
		.io_in_a_0(r_1019_0),
		.io_in_b_0(b_895_0),
		.io_in_d_0(b_1919_0),
		.io_in_control_0_dataflow(mesh_31_27_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_27_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_27_io_in_control_0_shift_b),
		.io_in_id_0(r_2943_0),
		.io_in_last_0(r_3967_0),
		.io_in_valid_0(r_1919_0),
		.io_out_a_0(_mesh_31_27_io_out_a_0),
		.io_out_c_0(_mesh_31_27_io_out_c_0),
		.io_out_b_0(_mesh_31_27_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_27_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_27_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_27_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_27_io_out_id_0),
		.io_out_last_0(_mesh_31_27_io_out_last_0),
		.io_out_valid_0(_mesh_31_27_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10390 == GlobalFiModInstNr[0]) || (10390 == GlobalFiModInstNr[1]) || (10390 == GlobalFiModInstNr[2]) || (10390 == GlobalFiModInstNr[3]))));
	Tile mesh_31_28(
		.clock(clock),
		.io_in_a_0(r_1020_0),
		.io_in_b_0(b_927_0),
		.io_in_d_0(b_1951_0),
		.io_in_control_0_dataflow(mesh_31_28_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_28_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_28_io_in_control_0_shift_b),
		.io_in_id_0(r_2975_0),
		.io_in_last_0(r_3999_0),
		.io_in_valid_0(r_1951_0),
		.io_out_a_0(_mesh_31_28_io_out_a_0),
		.io_out_c_0(_mesh_31_28_io_out_c_0),
		.io_out_b_0(_mesh_31_28_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_28_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_28_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_28_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_28_io_out_id_0),
		.io_out_last_0(_mesh_31_28_io_out_last_0),
		.io_out_valid_0(_mesh_31_28_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10391 == GlobalFiModInstNr[0]) || (10391 == GlobalFiModInstNr[1]) || (10391 == GlobalFiModInstNr[2]) || (10391 == GlobalFiModInstNr[3]))));
	Tile mesh_31_29(
		.clock(clock),
		.io_in_a_0(r_1021_0),
		.io_in_b_0(b_959_0),
		.io_in_d_0(b_1983_0),
		.io_in_control_0_dataflow(mesh_31_29_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_29_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_29_io_in_control_0_shift_b),
		.io_in_id_0(r_3007_0),
		.io_in_last_0(r_4031_0),
		.io_in_valid_0(r_1983_0),
		.io_out_a_0(_mesh_31_29_io_out_a_0),
		.io_out_c_0(_mesh_31_29_io_out_c_0),
		.io_out_b_0(_mesh_31_29_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_29_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_29_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_29_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_29_io_out_id_0),
		.io_out_last_0(_mesh_31_29_io_out_last_0),
		.io_out_valid_0(_mesh_31_29_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10392 == GlobalFiModInstNr[0]) || (10392 == GlobalFiModInstNr[1]) || (10392 == GlobalFiModInstNr[2]) || (10392 == GlobalFiModInstNr[3]))));
	Tile mesh_31_30(
		.clock(clock),
		.io_in_a_0(r_1022_0),
		.io_in_b_0(b_991_0),
		.io_in_d_0(b_2015_0),
		.io_in_control_0_dataflow(mesh_31_30_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_30_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_30_io_in_control_0_shift_b),
		.io_in_id_0(r_3039_0),
		.io_in_last_0(r_4063_0),
		.io_in_valid_0(r_2015_0),
		.io_out_a_0(_mesh_31_30_io_out_a_0),
		.io_out_c_0(_mesh_31_30_io_out_c_0),
		.io_out_b_0(_mesh_31_30_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_30_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_30_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_30_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_30_io_out_id_0),
		.io_out_last_0(_mesh_31_30_io_out_last_0),
		.io_out_valid_0(_mesh_31_30_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10393 == GlobalFiModInstNr[0]) || (10393 == GlobalFiModInstNr[1]) || (10393 == GlobalFiModInstNr[2]) || (10393 == GlobalFiModInstNr[3]))));
	Tile mesh_31_31(
		.clock(clock),
		.io_in_a_0(r_1023_0),
		.io_in_b_0(b_1023_0),
		.io_in_d_0(b_2047_0),
		.io_in_control_0_dataflow(mesh_31_31_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_31_31_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_31_31_io_in_control_0_shift_b),
		.io_in_id_0(r_3071_0),
		.io_in_last_0(r_4095_0),
		.io_in_valid_0(r_2047_0),
		.io_out_a_0(_mesh_31_31_io_out_a_0),
		.io_out_c_0(_mesh_31_31_io_out_c_0),
		.io_out_b_0(_mesh_31_31_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_31_31_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_31_31_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_31_31_io_out_control_0_shift),
		.io_out_id_0(_mesh_31_31_io_out_id_0),
		.io_out_last_0(_mesh_31_31_io_out_last_0),
		.io_out_valid_0(_mesh_31_31_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((10394 == GlobalFiModInstNr[0]) || (10394 == GlobalFiModInstNr[1]) || (10394 == GlobalFiModInstNr[2]) || (10394 == GlobalFiModInstNr[3]))));
	assign io_out_b_0_0 =( r_4096_0) ^ ((fiEnable && (9301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_1_0 =( r_4102_0) ^ ((fiEnable && (9302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_2_0 =( r_4108_0) ^ ((fiEnable && (9303 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_3_0 =( r_4114_0) ^ ((fiEnable && (9304 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_4_0 =( r_4120_0) ^ ((fiEnable && (9305 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_5_0 =( r_4126_0) ^ ((fiEnable && (9306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_6_0 =( r_4132_0) ^ ((fiEnable && (9307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_7_0 =( r_4138_0) ^ ((fiEnable && (9308 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_8_0 =( r_4144_0) ^ ((fiEnable && (9309 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_9_0 =( r_4150_0) ^ ((fiEnable && (9310 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_10_0 =( r_4156_0) ^ ((fiEnable && (9311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_11_0 =( r_4162_0) ^ ((fiEnable && (9312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_12_0 =( r_4168_0) ^ ((fiEnable && (9313 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_13_0 =( r_4174_0) ^ ((fiEnable && (9314 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_14_0 =( r_4180_0) ^ ((fiEnable && (9315 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_15_0 =( r_4186_0) ^ ((fiEnable && (9316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_16_0 =( r_4192_0) ^ ((fiEnable && (9317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_17_0 =( r_4198_0) ^ ((fiEnable && (9318 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_18_0 =( r_4204_0) ^ ((fiEnable && (9319 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_19_0 =( r_4210_0) ^ ((fiEnable && (9320 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_20_0 =( r_4216_0) ^ ((fiEnable && (9321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_21_0 =( r_4222_0) ^ ((fiEnable && (9322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_22_0 =( r_4228_0) ^ ((fiEnable && (9323 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_23_0 =( r_4234_0) ^ ((fiEnable && (9324 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_24_0 =( r_4240_0) ^ ((fiEnable && (9325 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_25_0 =( r_4246_0) ^ ((fiEnable && (9326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_26_0 =( r_4252_0) ^ ((fiEnable && (9327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_27_0 =( r_4258_0) ^ ((fiEnable && (9328 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_28_0 =( r_4264_0) ^ ((fiEnable && (9329 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_29_0 =( r_4270_0) ^ ((fiEnable && (9330 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_30_0 =( r_4276_0) ^ ((fiEnable && (9331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_31_0 =( r_4282_0) ^ ((fiEnable && (9332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_0_0 =( r_4097_0) ^ ((fiEnable && (9333 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_1_0 =( r_4103_0) ^ ((fiEnable && (9334 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_2_0 =( r_4109_0) ^ ((fiEnable && (9335 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_3_0 =( r_4115_0) ^ ((fiEnable && (9336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_4_0 =( r_4121_0) ^ ((fiEnable && (9337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_5_0 =( r_4127_0) ^ ((fiEnable && (9338 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_6_0 =( r_4133_0) ^ ((fiEnable && (9339 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_7_0 =( r_4139_0) ^ ((fiEnable && (9340 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_8_0 =( r_4145_0) ^ ((fiEnable && (9341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_9_0 =( r_4151_0) ^ ((fiEnable && (9342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_10_0 =( r_4157_0) ^ ((fiEnable && (9343 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_11_0 =( r_4163_0) ^ ((fiEnable && (9344 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_12_0 =( r_4169_0) ^ ((fiEnable && (9345 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_13_0 =( r_4175_0) ^ ((fiEnable && (9346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_14_0 =( r_4181_0) ^ ((fiEnable && (9347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_15_0 =( r_4187_0) ^ ((fiEnable && (9348 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_16_0 =( r_4193_0) ^ ((fiEnable && (9349 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_17_0 =( r_4199_0) ^ ((fiEnable && (9350 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_18_0 =( r_4205_0) ^ ((fiEnable && (9351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_19_0 =( r_4211_0) ^ ((fiEnable && (9352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_20_0 =( r_4217_0) ^ ((fiEnable && (9353 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_21_0 =( r_4223_0) ^ ((fiEnable && (9354 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_22_0 =( r_4229_0) ^ ((fiEnable && (9355 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_23_0 =( r_4235_0) ^ ((fiEnable && (9356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_24_0 =( r_4241_0) ^ ((fiEnable && (9357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_25_0 =( r_4247_0) ^ ((fiEnable && (9358 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_26_0 =( r_4253_0) ^ ((fiEnable && (9359 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_27_0 =( r_4259_0) ^ ((fiEnable && (9360 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_28_0 =( r_4265_0) ^ ((fiEnable && (9361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_29_0 =( r_4271_0) ^ ((fiEnable && (9362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_30_0 =( r_4277_0) ^ ((fiEnable && (9363 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_31_0 =( r_4283_0) ^ ((fiEnable && (9364 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_valid_0_0 =( r_4098_0) ^ ((fiEnable && (9365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_0_0_dataflow =( r_4099_0_dataflow) ^ ((fiEnable && (9366 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_id_0_0 =( r_4100_0) ^ ((fiEnable && (9367 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last_0_0 =( r_4101_0) ^ ((fiEnable && (9368 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
endmodule