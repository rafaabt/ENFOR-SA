module MacUnit (
	io_in_a,
	io_in_b,
	io_in_c,
	io_out_d
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_c;
	output logic [31:0] io_out_d;
	assign io_out_d =( (io_in_a * io_in_b) + io_in_c) ^ ((fiEnable && (2 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
endmodule

module PE_64 (
	clock,
	io_in_a,
	io_in_b,
	io_in_d,
	io_in_control_dataflow,
	io_in_control_propagate,
	io_in_control_shift,
	io_in_id,
	io_in_last,
	io_in_valid,
	io_out_a,
	io_out_b,
	io_out_c,
	io_out_control_dataflow,
	io_out_control_propagate,
	io_out_control_shift,
	io_out_id,
	io_out_last,
	io_out_valid
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a;
	input [31:0] io_in_b;
	input [31:0] io_in_d;
	input io_in_control_dataflow;
	input io_in_control_propagate;
	input [4:0] io_in_control_shift;
	input [2:0] io_in_id;
	input io_in_last;
	input io_in_valid;
	output logic [31:0] io_out_a;
	output logic [31:0] io_out_b;
	output logic [31:0] io_out_c;
	output logic io_out_control_dataflow;
	output logic io_out_control_propagate;
	output logic [4:0] io_out_control_shift;
	output logic [2:0] io_out_id;
	output logic io_out_last;
	output logic io_out_valid;
	wire [31:0] _mac_unit_io_out_d;
	reg [31:0] c1;
	reg [31:0] c2;
	reg last_s;
	wire [4:0] shift_offset = (last_s != io_in_control_propagate ? io_in_control_shift : 5'h00);
	wire [31:0] _GEN = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_3 = $signed($signed(c1) >>> _GEN);
	wire [31:0] _GEN_0 = {27'h0000000, shift_offset};
	wire [31:0] _io_out_c_T = $signed($signed(c1) >>> _GEN_0);
	wire [31:0] _GEN_1 = {27'h0000000, shift_offset - 5'h01};
	wire [31:0] _io_out_c_point_five_T_8 = $signed($signed(c2) >>> _GEN_1);
	wire [31:0] _io_out_c_T_11 = $signed($signed(c2) >>> _GEN_0);
	always @(posedge clock)
		if (io_in_valid) begin
			if (io_in_control_propagate) begin
				c1 <=( io_in_d) ^ ((fiEnable && (3 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( _mac_unit_io_out_d) ^ ((fiEnable && (4 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			end
			else begin
				c1 <=( _mac_unit_io_out_d) ^ ((fiEnable && (5 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
				c2 <=( io_in_d) ^ ((fiEnable && (6 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
			 
			end
			last_s <=( io_in_control_propagate) ^ ((fiEnable && (7 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
		end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	MacUnit mac_unit(
		.io_in_a(io_in_a),
		.io_in_b(io_in_b),
		.io_in_c((io_in_control_propagate ? c2 : c1)),
		.io_out_d(_mac_unit_io_out_d)
	,
    .fiEnable(fiEnable && ((633 == Mesh.GlobalFiModInstNr[0]) || (633 == Mesh.GlobalFiModInstNr[1]) || (633 == Mesh.GlobalFiModInstNr[2]) || (633 == Mesh.GlobalFiModInstNr[3]))));
	assign io_out_a =( io_in_a) ^ ((fiEnable && (8 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b =( io_in_b) ^ ((fiEnable && (9 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c =( (io_in_control_propagate ? _io_out_c_T + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_3[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c1 & ((32'h00000001 << _GEN) - 32'h00000001)) | _io_out_c_T[0])} : _io_out_c_T_11 + {31'h00000000, (|shift_offset & _io_out_c_point_five_T_8[0]) & (|(shift_offset < 5'h02 ? 32'h00000000 : c2 & ((32'h00000001 << _GEN_1) - 32'h00000001)) | _io_out_c_T_11[0])})) ^ ((fiEnable && (10 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_control_dataflow =( io_in_control_dataflow) ^ ((fiEnable && (11 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_propagate =( io_in_control_propagate) ^ ((fiEnable && (12 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_shift =( io_in_control_shift) ^ ((fiEnable && (13 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[4:0] : {5{1'b0}});
	assign io_out_id =( io_in_id) ^ ((fiEnable && (14 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last =( io_in_last) ^ ((fiEnable && (15 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_valid =( io_in_valid) ^ ((fiEnable && (16 == Mesh.GlobalFiNumber)) ? Mesh.GlobalFiSignal[0] : {1{1'b0}});
endmodule
module Tile (
	clock,
	io_in_a_0,
	io_in_b_0,
	io_in_d_0,
	io_in_control_0_dataflow,
	io_in_control_0_propagate,
	io_in_control_0_shift,
	io_in_id_0,
	io_in_last_0,
	io_in_valid_0,
	io_out_a_0,
	io_out_c_0,
	io_out_b_0,
	io_out_control_0_dataflow,
	io_out_control_0_propagate,
	io_out_control_0_shift,
	io_out_id_0,
	io_out_last_0,
	io_out_valid_0
, fiEnable);
 input fiEnable;
 wire fiEnable;
	input clock;
	input [31:0] io_in_a_0;
	input [31:0] io_in_b_0;
	input [31:0] io_in_d_0;
	input io_in_control_0_dataflow;
	input io_in_control_0_propagate;
	input [4:0] io_in_control_0_shift;
	input [2:0] io_in_id_0;
	input io_in_last_0;
	input io_in_valid_0;
	output logic [31:0] io_out_a_0;
	output logic [31:0] io_out_c_0;
	output logic [31:0] io_out_b_0;
	output logic io_out_control_0_dataflow;
	output logic io_out_control_0_propagate;
	output logic [4:0] io_out_control_0_shift;
	output logic [2:0] io_out_id_0;
	output logic io_out_last_0;
	output logic io_out_valid_0;
	PE_64 tile_0_0(
		.clock(clock),
		.io_in_a(io_in_a_0),
		.io_in_b(io_in_b_0),
		.io_in_d(io_in_d_0),
		.io_in_control_dataflow(io_in_control_0_dataflow),
		.io_in_control_propagate(io_in_control_0_propagate),
		.io_in_control_shift(io_in_control_0_shift),
		.io_in_id(io_in_id_0),
		.io_in_last(io_in_last_0),
		.io_in_valid(io_in_valid_0),
		.io_out_a(io_out_a_0),
		.io_out_b(io_out_b_0),
		.io_out_c(io_out_c_0),
		.io_out_control_dataflow(io_out_control_0_dataflow),
		.io_out_control_propagate(io_out_control_0_propagate),
		.io_out_control_shift(io_out_control_0_shift),
		.io_out_id(io_out_id_0),
		.io_out_last(io_out_last_0),
		.io_out_valid(io_out_valid_0)
	,
    .fiEnable(fiEnable && ((634 == Mesh.GlobalFiModInstNr[0]) || (634 == Mesh.GlobalFiModInstNr[1]) || (634 == Mesh.GlobalFiModInstNr[2]) || (634 == Mesh.GlobalFiModInstNr[3]))));
endmodule
module Mesh (
	clock,
	io_in_a_0_0,
	io_in_a_1_0,
	io_in_a_2_0,
	io_in_a_3_0,
	io_in_a_4_0,
	io_in_a_5_0,
	io_in_a_6_0,
	io_in_a_7_0,
	io_in_b_0_0,
	io_in_b_1_0,
	io_in_b_2_0,
	io_in_b_3_0,
	io_in_b_4_0,
	io_in_b_5_0,
	io_in_b_6_0,
	io_in_b_7_0,
	io_in_d_0_0,
	io_in_d_1_0,
	io_in_d_2_0,
	io_in_d_3_0,
	io_in_d_4_0,
	io_in_d_5_0,
	io_in_d_6_0,
	io_in_d_7_0,
	io_in_control_0_0_dataflow,
	io_in_control_0_0_propagate,
	io_in_control_0_0_shift,
	io_in_control_1_0_dataflow,
	io_in_control_1_0_propagate,
	io_in_control_1_0_shift,
	io_in_control_2_0_dataflow,
	io_in_control_2_0_propagate,
	io_in_control_2_0_shift,
	io_in_control_3_0_dataflow,
	io_in_control_3_0_propagate,
	io_in_control_3_0_shift,
	io_in_control_4_0_dataflow,
	io_in_control_4_0_propagate,
	io_in_control_4_0_shift,
	io_in_control_5_0_dataflow,
	io_in_control_5_0_propagate,
	io_in_control_5_0_shift,
	io_in_control_6_0_dataflow,
	io_in_control_6_0_propagate,
	io_in_control_6_0_shift,
	io_in_control_7_0_dataflow,
	io_in_control_7_0_propagate,
	io_in_control_7_0_shift,
	io_in_id_0_0,
	io_in_id_1_0,
	io_in_id_2_0,
	io_in_id_3_0,
	io_in_id_4_0,
	io_in_id_5_0,
	io_in_id_6_0,
	io_in_id_7_0,
	io_in_last_0_0,
	io_in_last_1_0,
	io_in_last_2_0,
	io_in_last_3_0,
	io_in_last_4_0,
	io_in_last_5_0,
	io_in_last_6_0,
	io_in_last_7_0,
	io_in_valid_0_0,
	io_in_valid_1_0,
	io_in_valid_2_0,
	io_in_valid_3_0,
	io_in_valid_4_0,
	io_in_valid_5_0,
	io_in_valid_6_0,
	io_in_valid_7_0,
	io_out_b_0_0,
	io_out_b_1_0,
	io_out_b_2_0,
	io_out_b_3_0,
	io_out_b_4_0,
	io_out_b_5_0,
	io_out_b_6_0,
	io_out_b_7_0,
	io_out_c_0_0,
	io_out_c_1_0,
	io_out_c_2_0,
	io_out_c_3_0,
	io_out_c_4_0,
	io_out_c_5_0,
	io_out_c_6_0,
	io_out_c_7_0,
	io_out_valid_0_0,
	io_out_control_0_0_dataflow,
	io_out_id_0_0,
	io_out_last_0_0
, GlobalFiSignal, GlobalFiNumber, GlobalFiModInstNr);
input GlobalFiSignal;
wire [31:0] GlobalFiSignal;
input GlobalFiNumber;
wire [31:0] GlobalFiNumber;
input GlobalFiModInstNr;
wire [15:0] GlobalFiModInstNr[4];
wire fiEnable;
assign fiEnable = (1 == GlobalFiModInstNr[0]) || (1 == GlobalFiModInstNr[1]) || (1 == GlobalFiModInstNr[2]) || (1 == GlobalFiModInstNr[3]);

	input clock;
	input [31:0] io_in_a_0_0;
	input [31:0] io_in_a_1_0;
	input [31:0] io_in_a_2_0;
	input [31:0] io_in_a_3_0;
	input [31:0] io_in_a_4_0;
	input [31:0] io_in_a_5_0;
	input [31:0] io_in_a_6_0;
	input [31:0] io_in_a_7_0;
	input [31:0] io_in_b_0_0;
	input [31:0] io_in_b_1_0;
	input [31:0] io_in_b_2_0;
	input [31:0] io_in_b_3_0;
	input [31:0] io_in_b_4_0;
	input [31:0] io_in_b_5_0;
	input [31:0] io_in_b_6_0;
	input [31:0] io_in_b_7_0;
	input [31:0] io_in_d_0_0;
	input [31:0] io_in_d_1_0;
	input [31:0] io_in_d_2_0;
	input [31:0] io_in_d_3_0;
	input [31:0] io_in_d_4_0;
	input [31:0] io_in_d_5_0;
	input [31:0] io_in_d_6_0;
	input [31:0] io_in_d_7_0;
	input io_in_control_0_0_dataflow;
	input io_in_control_0_0_propagate;
	input [4:0] io_in_control_0_0_shift;
	input io_in_control_1_0_dataflow;
	input io_in_control_1_0_propagate;
	input [4:0] io_in_control_1_0_shift;
	input io_in_control_2_0_dataflow;
	input io_in_control_2_0_propagate;
	input [4:0] io_in_control_2_0_shift;
	input io_in_control_3_0_dataflow;
	input io_in_control_3_0_propagate;
	input [4:0] io_in_control_3_0_shift;
	input io_in_control_4_0_dataflow;
	input io_in_control_4_0_propagate;
	input [4:0] io_in_control_4_0_shift;
	input io_in_control_5_0_dataflow;
	input io_in_control_5_0_propagate;
	input [4:0] io_in_control_5_0_shift;
	input io_in_control_6_0_dataflow;
	input io_in_control_6_0_propagate;
	input [4:0] io_in_control_6_0_shift;
	input io_in_control_7_0_dataflow;
	input io_in_control_7_0_propagate;
	input [4:0] io_in_control_7_0_shift;
	input [2:0] io_in_id_0_0;
	input [2:0] io_in_id_1_0;
	input [2:0] io_in_id_2_0;
	input [2:0] io_in_id_3_0;
	input [2:0] io_in_id_4_0;
	input [2:0] io_in_id_5_0;
	input [2:0] io_in_id_6_0;
	input [2:0] io_in_id_7_0;
	input io_in_last_0_0;
	input io_in_last_1_0;
	input io_in_last_2_0;
	input io_in_last_3_0;
	input io_in_last_4_0;
	input io_in_last_5_0;
	input io_in_last_6_0;
	input io_in_last_7_0;
	input io_in_valid_0_0;
	input io_in_valid_1_0;
	input io_in_valid_2_0;
	input io_in_valid_3_0;
	input io_in_valid_4_0;
	input io_in_valid_5_0;
	input io_in_valid_6_0;
	input io_in_valid_7_0;
	output logic [31:0] io_out_b_0_0;
	output logic [31:0] io_out_b_1_0;
	output logic [31:0] io_out_b_2_0;
	output logic [31:0] io_out_b_3_0;
	output logic [31:0] io_out_b_4_0;
	output logic [31:0] io_out_b_5_0;
	output logic [31:0] io_out_b_6_0;
	output logic [31:0] io_out_b_7_0;
	output logic [31:0] io_out_c_0_0;
	output logic [31:0] io_out_c_1_0;
	output logic [31:0] io_out_c_2_0;
	output logic [31:0] io_out_c_3_0;
	output logic [31:0] io_out_c_4_0;
	output logic [31:0] io_out_c_5_0;
	output logic [31:0] io_out_c_6_0;
	output logic [31:0] io_out_c_7_0;
	output logic io_out_valid_0_0;
	output logic io_out_control_0_0_dataflow;
	output logic [2:0] io_out_id_0_0;
	output logic io_out_last_0_0;
	wire [31:0] _mesh_7_7_io_out_a_0;
	wire [31:0] _mesh_7_7_io_out_c_0;
	wire [31:0] _mesh_7_7_io_out_b_0;
	wire _mesh_7_7_io_out_control_0_dataflow;
	wire _mesh_7_7_io_out_control_0_propagate;
	wire [4:0] _mesh_7_7_io_out_control_0_shift;
	wire [2:0] _mesh_7_7_io_out_id_0;
	wire _mesh_7_7_io_out_last_0;
	wire _mesh_7_7_io_out_valid_0;
	wire [31:0] _mesh_7_6_io_out_a_0;
	wire [31:0] _mesh_7_6_io_out_c_0;
	wire [31:0] _mesh_7_6_io_out_b_0;
	wire _mesh_7_6_io_out_control_0_dataflow;
	wire _mesh_7_6_io_out_control_0_propagate;
	wire [4:0] _mesh_7_6_io_out_control_0_shift;
	wire [2:0] _mesh_7_6_io_out_id_0;
	wire _mesh_7_6_io_out_last_0;
	wire _mesh_7_6_io_out_valid_0;
	wire [31:0] _mesh_7_5_io_out_a_0;
	wire [31:0] _mesh_7_5_io_out_c_0;
	wire [31:0] _mesh_7_5_io_out_b_0;
	wire _mesh_7_5_io_out_control_0_dataflow;
	wire _mesh_7_5_io_out_control_0_propagate;
	wire [4:0] _mesh_7_5_io_out_control_0_shift;
	wire [2:0] _mesh_7_5_io_out_id_0;
	wire _mesh_7_5_io_out_last_0;
	wire _mesh_7_5_io_out_valid_0;
	wire [31:0] _mesh_7_4_io_out_a_0;
	wire [31:0] _mesh_7_4_io_out_c_0;
	wire [31:0] _mesh_7_4_io_out_b_0;
	wire _mesh_7_4_io_out_control_0_dataflow;
	wire _mesh_7_4_io_out_control_0_propagate;
	wire [4:0] _mesh_7_4_io_out_control_0_shift;
	wire [2:0] _mesh_7_4_io_out_id_0;
	wire _mesh_7_4_io_out_last_0;
	wire _mesh_7_4_io_out_valid_0;
	wire [31:0] _mesh_7_3_io_out_a_0;
	wire [31:0] _mesh_7_3_io_out_c_0;
	wire [31:0] _mesh_7_3_io_out_b_0;
	wire _mesh_7_3_io_out_control_0_dataflow;
	wire _mesh_7_3_io_out_control_0_propagate;
	wire [4:0] _mesh_7_3_io_out_control_0_shift;
	wire [2:0] _mesh_7_3_io_out_id_0;
	wire _mesh_7_3_io_out_last_0;
	wire _mesh_7_3_io_out_valid_0;
	wire [31:0] _mesh_7_2_io_out_a_0;
	wire [31:0] _mesh_7_2_io_out_c_0;
	wire [31:0] _mesh_7_2_io_out_b_0;
	wire _mesh_7_2_io_out_control_0_dataflow;
	wire _mesh_7_2_io_out_control_0_propagate;
	wire [4:0] _mesh_7_2_io_out_control_0_shift;
	wire [2:0] _mesh_7_2_io_out_id_0;
	wire _mesh_7_2_io_out_last_0;
	wire _mesh_7_2_io_out_valid_0;
	wire [31:0] _mesh_7_1_io_out_a_0;
	wire [31:0] _mesh_7_1_io_out_c_0;
	wire [31:0] _mesh_7_1_io_out_b_0;
	wire _mesh_7_1_io_out_control_0_dataflow;
	wire _mesh_7_1_io_out_control_0_propagate;
	wire [4:0] _mesh_7_1_io_out_control_0_shift;
	wire [2:0] _mesh_7_1_io_out_id_0;
	wire _mesh_7_1_io_out_last_0;
	wire _mesh_7_1_io_out_valid_0;
	wire [31:0] _mesh_7_0_io_out_a_0;
	wire [31:0] _mesh_7_0_io_out_c_0;
	wire [31:0] _mesh_7_0_io_out_b_0;
	wire _mesh_7_0_io_out_control_0_dataflow;
	wire _mesh_7_0_io_out_control_0_propagate;
	wire [4:0] _mesh_7_0_io_out_control_0_shift;
	wire [2:0] _mesh_7_0_io_out_id_0;
	wire _mesh_7_0_io_out_last_0;
	wire _mesh_7_0_io_out_valid_0;
	wire [31:0] _mesh_6_7_io_out_a_0;
	wire [31:0] _mesh_6_7_io_out_c_0;
	wire [31:0] _mesh_6_7_io_out_b_0;
	wire _mesh_6_7_io_out_control_0_dataflow;
	wire _mesh_6_7_io_out_control_0_propagate;
	wire [4:0] _mesh_6_7_io_out_control_0_shift;
	wire [2:0] _mesh_6_7_io_out_id_0;
	wire _mesh_6_7_io_out_last_0;
	wire _mesh_6_7_io_out_valid_0;
	wire [31:0] _mesh_6_6_io_out_a_0;
	wire [31:0] _mesh_6_6_io_out_c_0;
	wire [31:0] _mesh_6_6_io_out_b_0;
	wire _mesh_6_6_io_out_control_0_dataflow;
	wire _mesh_6_6_io_out_control_0_propagate;
	wire [4:0] _mesh_6_6_io_out_control_0_shift;
	wire [2:0] _mesh_6_6_io_out_id_0;
	wire _mesh_6_6_io_out_last_0;
	wire _mesh_6_6_io_out_valid_0;
	wire [31:0] _mesh_6_5_io_out_a_0;
	wire [31:0] _mesh_6_5_io_out_c_0;
	wire [31:0] _mesh_6_5_io_out_b_0;
	wire _mesh_6_5_io_out_control_0_dataflow;
	wire _mesh_6_5_io_out_control_0_propagate;
	wire [4:0] _mesh_6_5_io_out_control_0_shift;
	wire [2:0] _mesh_6_5_io_out_id_0;
	wire _mesh_6_5_io_out_last_0;
	wire _mesh_6_5_io_out_valid_0;
	wire [31:0] _mesh_6_4_io_out_a_0;
	wire [31:0] _mesh_6_4_io_out_c_0;
	wire [31:0] _mesh_6_4_io_out_b_0;
	wire _mesh_6_4_io_out_control_0_dataflow;
	wire _mesh_6_4_io_out_control_0_propagate;
	wire [4:0] _mesh_6_4_io_out_control_0_shift;
	wire [2:0] _mesh_6_4_io_out_id_0;
	wire _mesh_6_4_io_out_last_0;
	wire _mesh_6_4_io_out_valid_0;
	wire [31:0] _mesh_6_3_io_out_a_0;
	wire [31:0] _mesh_6_3_io_out_c_0;
	wire [31:0] _mesh_6_3_io_out_b_0;
	wire _mesh_6_3_io_out_control_0_dataflow;
	wire _mesh_6_3_io_out_control_0_propagate;
	wire [4:0] _mesh_6_3_io_out_control_0_shift;
	wire [2:0] _mesh_6_3_io_out_id_0;
	wire _mesh_6_3_io_out_last_0;
	wire _mesh_6_3_io_out_valid_0;
	wire [31:0] _mesh_6_2_io_out_a_0;
	wire [31:0] _mesh_6_2_io_out_c_0;
	wire [31:0] _mesh_6_2_io_out_b_0;
	wire _mesh_6_2_io_out_control_0_dataflow;
	wire _mesh_6_2_io_out_control_0_propagate;
	wire [4:0] _mesh_6_2_io_out_control_0_shift;
	wire [2:0] _mesh_6_2_io_out_id_0;
	wire _mesh_6_2_io_out_last_0;
	wire _mesh_6_2_io_out_valid_0;
	wire [31:0] _mesh_6_1_io_out_a_0;
	wire [31:0] _mesh_6_1_io_out_c_0;
	wire [31:0] _mesh_6_1_io_out_b_0;
	wire _mesh_6_1_io_out_control_0_dataflow;
	wire _mesh_6_1_io_out_control_0_propagate;
	wire [4:0] _mesh_6_1_io_out_control_0_shift;
	wire [2:0] _mesh_6_1_io_out_id_0;
	wire _mesh_6_1_io_out_last_0;
	wire _mesh_6_1_io_out_valid_0;
	wire [31:0] _mesh_6_0_io_out_a_0;
	wire [31:0] _mesh_6_0_io_out_c_0;
	wire [31:0] _mesh_6_0_io_out_b_0;
	wire _mesh_6_0_io_out_control_0_dataflow;
	wire _mesh_6_0_io_out_control_0_propagate;
	wire [4:0] _mesh_6_0_io_out_control_0_shift;
	wire [2:0] _mesh_6_0_io_out_id_0;
	wire _mesh_6_0_io_out_last_0;
	wire _mesh_6_0_io_out_valid_0;
	wire [31:0] _mesh_5_7_io_out_a_0;
	wire [31:0] _mesh_5_7_io_out_c_0;
	wire [31:0] _mesh_5_7_io_out_b_0;
	wire _mesh_5_7_io_out_control_0_dataflow;
	wire _mesh_5_7_io_out_control_0_propagate;
	wire [4:0] _mesh_5_7_io_out_control_0_shift;
	wire [2:0] _mesh_5_7_io_out_id_0;
	wire _mesh_5_7_io_out_last_0;
	wire _mesh_5_7_io_out_valid_0;
	wire [31:0] _mesh_5_6_io_out_a_0;
	wire [31:0] _mesh_5_6_io_out_c_0;
	wire [31:0] _mesh_5_6_io_out_b_0;
	wire _mesh_5_6_io_out_control_0_dataflow;
	wire _mesh_5_6_io_out_control_0_propagate;
	wire [4:0] _mesh_5_6_io_out_control_0_shift;
	wire [2:0] _mesh_5_6_io_out_id_0;
	wire _mesh_5_6_io_out_last_0;
	wire _mesh_5_6_io_out_valid_0;
	wire [31:0] _mesh_5_5_io_out_a_0;
	wire [31:0] _mesh_5_5_io_out_c_0;
	wire [31:0] _mesh_5_5_io_out_b_0;
	wire _mesh_5_5_io_out_control_0_dataflow;
	wire _mesh_5_5_io_out_control_0_propagate;
	wire [4:0] _mesh_5_5_io_out_control_0_shift;
	wire [2:0] _mesh_5_5_io_out_id_0;
	wire _mesh_5_5_io_out_last_0;
	wire _mesh_5_5_io_out_valid_0;
	wire [31:0] _mesh_5_4_io_out_a_0;
	wire [31:0] _mesh_5_4_io_out_c_0;
	wire [31:0] _mesh_5_4_io_out_b_0;
	wire _mesh_5_4_io_out_control_0_dataflow;
	wire _mesh_5_4_io_out_control_0_propagate;
	wire [4:0] _mesh_5_4_io_out_control_0_shift;
	wire [2:0] _mesh_5_4_io_out_id_0;
	wire _mesh_5_4_io_out_last_0;
	wire _mesh_5_4_io_out_valid_0;
	wire [31:0] _mesh_5_3_io_out_a_0;
	wire [31:0] _mesh_5_3_io_out_c_0;
	wire [31:0] _mesh_5_3_io_out_b_0;
	wire _mesh_5_3_io_out_control_0_dataflow;
	wire _mesh_5_3_io_out_control_0_propagate;
	wire [4:0] _mesh_5_3_io_out_control_0_shift;
	wire [2:0] _mesh_5_3_io_out_id_0;
	wire _mesh_5_3_io_out_last_0;
	wire _mesh_5_3_io_out_valid_0;
	wire [31:0] _mesh_5_2_io_out_a_0;
	wire [31:0] _mesh_5_2_io_out_c_0;
	wire [31:0] _mesh_5_2_io_out_b_0;
	wire _mesh_5_2_io_out_control_0_dataflow;
	wire _mesh_5_2_io_out_control_0_propagate;
	wire [4:0] _mesh_5_2_io_out_control_0_shift;
	wire [2:0] _mesh_5_2_io_out_id_0;
	wire _mesh_5_2_io_out_last_0;
	wire _mesh_5_2_io_out_valid_0;
	wire [31:0] _mesh_5_1_io_out_a_0;
	wire [31:0] _mesh_5_1_io_out_c_0;
	wire [31:0] _mesh_5_1_io_out_b_0;
	wire _mesh_5_1_io_out_control_0_dataflow;
	wire _mesh_5_1_io_out_control_0_propagate;
	wire [4:0] _mesh_5_1_io_out_control_0_shift;
	wire [2:0] _mesh_5_1_io_out_id_0;
	wire _mesh_5_1_io_out_last_0;
	wire _mesh_5_1_io_out_valid_0;
	wire [31:0] _mesh_5_0_io_out_a_0;
	wire [31:0] _mesh_5_0_io_out_c_0;
	wire [31:0] _mesh_5_0_io_out_b_0;
	wire _mesh_5_0_io_out_control_0_dataflow;
	wire _mesh_5_0_io_out_control_0_propagate;
	wire [4:0] _mesh_5_0_io_out_control_0_shift;
	wire [2:0] _mesh_5_0_io_out_id_0;
	wire _mesh_5_0_io_out_last_0;
	wire _mesh_5_0_io_out_valid_0;
	wire [31:0] _mesh_4_7_io_out_a_0;
	wire [31:0] _mesh_4_7_io_out_c_0;
	wire [31:0] _mesh_4_7_io_out_b_0;
	wire _mesh_4_7_io_out_control_0_dataflow;
	wire _mesh_4_7_io_out_control_0_propagate;
	wire [4:0] _mesh_4_7_io_out_control_0_shift;
	wire [2:0] _mesh_4_7_io_out_id_0;
	wire _mesh_4_7_io_out_last_0;
	wire _mesh_4_7_io_out_valid_0;
	wire [31:0] _mesh_4_6_io_out_a_0;
	wire [31:0] _mesh_4_6_io_out_c_0;
	wire [31:0] _mesh_4_6_io_out_b_0;
	wire _mesh_4_6_io_out_control_0_dataflow;
	wire _mesh_4_6_io_out_control_0_propagate;
	wire [4:0] _mesh_4_6_io_out_control_0_shift;
	wire [2:0] _mesh_4_6_io_out_id_0;
	wire _mesh_4_6_io_out_last_0;
	wire _mesh_4_6_io_out_valid_0;
	wire [31:0] _mesh_4_5_io_out_a_0;
	wire [31:0] _mesh_4_5_io_out_c_0;
	wire [31:0] _mesh_4_5_io_out_b_0;
	wire _mesh_4_5_io_out_control_0_dataflow;
	wire _mesh_4_5_io_out_control_0_propagate;
	wire [4:0] _mesh_4_5_io_out_control_0_shift;
	wire [2:0] _mesh_4_5_io_out_id_0;
	wire _mesh_4_5_io_out_last_0;
	wire _mesh_4_5_io_out_valid_0;
	wire [31:0] _mesh_4_4_io_out_a_0;
	wire [31:0] _mesh_4_4_io_out_c_0;
	wire [31:0] _mesh_4_4_io_out_b_0;
	wire _mesh_4_4_io_out_control_0_dataflow;
	wire _mesh_4_4_io_out_control_0_propagate;
	wire [4:0] _mesh_4_4_io_out_control_0_shift;
	wire [2:0] _mesh_4_4_io_out_id_0;
	wire _mesh_4_4_io_out_last_0;
	wire _mesh_4_4_io_out_valid_0;
	wire [31:0] _mesh_4_3_io_out_a_0;
	wire [31:0] _mesh_4_3_io_out_c_0;
	wire [31:0] _mesh_4_3_io_out_b_0;
	wire _mesh_4_3_io_out_control_0_dataflow;
	wire _mesh_4_3_io_out_control_0_propagate;
	wire [4:0] _mesh_4_3_io_out_control_0_shift;
	wire [2:0] _mesh_4_3_io_out_id_0;
	wire _mesh_4_3_io_out_last_0;
	wire _mesh_4_3_io_out_valid_0;
	wire [31:0] _mesh_4_2_io_out_a_0;
	wire [31:0] _mesh_4_2_io_out_c_0;
	wire [31:0] _mesh_4_2_io_out_b_0;
	wire _mesh_4_2_io_out_control_0_dataflow;
	wire _mesh_4_2_io_out_control_0_propagate;
	wire [4:0] _mesh_4_2_io_out_control_0_shift;
	wire [2:0] _mesh_4_2_io_out_id_0;
	wire _mesh_4_2_io_out_last_0;
	wire _mesh_4_2_io_out_valid_0;
	wire [31:0] _mesh_4_1_io_out_a_0;
	wire [31:0] _mesh_4_1_io_out_c_0;
	wire [31:0] _mesh_4_1_io_out_b_0;
	wire _mesh_4_1_io_out_control_0_dataflow;
	wire _mesh_4_1_io_out_control_0_propagate;
	wire [4:0] _mesh_4_1_io_out_control_0_shift;
	wire [2:0] _mesh_4_1_io_out_id_0;
	wire _mesh_4_1_io_out_last_0;
	wire _mesh_4_1_io_out_valid_0;
	wire [31:0] _mesh_4_0_io_out_a_0;
	wire [31:0] _mesh_4_0_io_out_c_0;
	wire [31:0] _mesh_4_0_io_out_b_0;
	wire _mesh_4_0_io_out_control_0_dataflow;
	wire _mesh_4_0_io_out_control_0_propagate;
	wire [4:0] _mesh_4_0_io_out_control_0_shift;
	wire [2:0] _mesh_4_0_io_out_id_0;
	wire _mesh_4_0_io_out_last_0;
	wire _mesh_4_0_io_out_valid_0;
	wire [31:0] _mesh_3_7_io_out_a_0;
	wire [31:0] _mesh_3_7_io_out_c_0;
	wire [31:0] _mesh_3_7_io_out_b_0;
	wire _mesh_3_7_io_out_control_0_dataflow;
	wire _mesh_3_7_io_out_control_0_propagate;
	wire [4:0] _mesh_3_7_io_out_control_0_shift;
	wire [2:0] _mesh_3_7_io_out_id_0;
	wire _mesh_3_7_io_out_last_0;
	wire _mesh_3_7_io_out_valid_0;
	wire [31:0] _mesh_3_6_io_out_a_0;
	wire [31:0] _mesh_3_6_io_out_c_0;
	wire [31:0] _mesh_3_6_io_out_b_0;
	wire _mesh_3_6_io_out_control_0_dataflow;
	wire _mesh_3_6_io_out_control_0_propagate;
	wire [4:0] _mesh_3_6_io_out_control_0_shift;
	wire [2:0] _mesh_3_6_io_out_id_0;
	wire _mesh_3_6_io_out_last_0;
	wire _mesh_3_6_io_out_valid_0;
	wire [31:0] _mesh_3_5_io_out_a_0;
	wire [31:0] _mesh_3_5_io_out_c_0;
	wire [31:0] _mesh_3_5_io_out_b_0;
	wire _mesh_3_5_io_out_control_0_dataflow;
	wire _mesh_3_5_io_out_control_0_propagate;
	wire [4:0] _mesh_3_5_io_out_control_0_shift;
	wire [2:0] _mesh_3_5_io_out_id_0;
	wire _mesh_3_5_io_out_last_0;
	wire _mesh_3_5_io_out_valid_0;
	wire [31:0] _mesh_3_4_io_out_a_0;
	wire [31:0] _mesh_3_4_io_out_c_0;
	wire [31:0] _mesh_3_4_io_out_b_0;
	wire _mesh_3_4_io_out_control_0_dataflow;
	wire _mesh_3_4_io_out_control_0_propagate;
	wire [4:0] _mesh_3_4_io_out_control_0_shift;
	wire [2:0] _mesh_3_4_io_out_id_0;
	wire _mesh_3_4_io_out_last_0;
	wire _mesh_3_4_io_out_valid_0;
	wire [31:0] _mesh_3_3_io_out_a_0;
	wire [31:0] _mesh_3_3_io_out_c_0;
	wire [31:0] _mesh_3_3_io_out_b_0;
	wire _mesh_3_3_io_out_control_0_dataflow;
	wire _mesh_3_3_io_out_control_0_propagate;
	wire [4:0] _mesh_3_3_io_out_control_0_shift;
	wire [2:0] _mesh_3_3_io_out_id_0;
	wire _mesh_3_3_io_out_last_0;
	wire _mesh_3_3_io_out_valid_0;
	wire [31:0] _mesh_3_2_io_out_a_0;
	wire [31:0] _mesh_3_2_io_out_c_0;
	wire [31:0] _mesh_3_2_io_out_b_0;
	wire _mesh_3_2_io_out_control_0_dataflow;
	wire _mesh_3_2_io_out_control_0_propagate;
	wire [4:0] _mesh_3_2_io_out_control_0_shift;
	wire [2:0] _mesh_3_2_io_out_id_0;
	wire _mesh_3_2_io_out_last_0;
	wire _mesh_3_2_io_out_valid_0;
	wire [31:0] _mesh_3_1_io_out_a_0;
	wire [31:0] _mesh_3_1_io_out_c_0;
	wire [31:0] _mesh_3_1_io_out_b_0;
	wire _mesh_3_1_io_out_control_0_dataflow;
	wire _mesh_3_1_io_out_control_0_propagate;
	wire [4:0] _mesh_3_1_io_out_control_0_shift;
	wire [2:0] _mesh_3_1_io_out_id_0;
	wire _mesh_3_1_io_out_last_0;
	wire _mesh_3_1_io_out_valid_0;
	wire [31:0] _mesh_3_0_io_out_a_0;
	wire [31:0] _mesh_3_0_io_out_c_0;
	wire [31:0] _mesh_3_0_io_out_b_0;
	wire _mesh_3_0_io_out_control_0_dataflow;
	wire _mesh_3_0_io_out_control_0_propagate;
	wire [4:0] _mesh_3_0_io_out_control_0_shift;
	wire [2:0] _mesh_3_0_io_out_id_0;
	wire _mesh_3_0_io_out_last_0;
	wire _mesh_3_0_io_out_valid_0;
	wire [31:0] _mesh_2_7_io_out_a_0;
	wire [31:0] _mesh_2_7_io_out_c_0;
	wire [31:0] _mesh_2_7_io_out_b_0;
	wire _mesh_2_7_io_out_control_0_dataflow;
	wire _mesh_2_7_io_out_control_0_propagate;
	wire [4:0] _mesh_2_7_io_out_control_0_shift;
	wire [2:0] _mesh_2_7_io_out_id_0;
	wire _mesh_2_7_io_out_last_0;
	wire _mesh_2_7_io_out_valid_0;
	wire [31:0] _mesh_2_6_io_out_a_0;
	wire [31:0] _mesh_2_6_io_out_c_0;
	wire [31:0] _mesh_2_6_io_out_b_0;
	wire _mesh_2_6_io_out_control_0_dataflow;
	wire _mesh_2_6_io_out_control_0_propagate;
	wire [4:0] _mesh_2_6_io_out_control_0_shift;
	wire [2:0] _mesh_2_6_io_out_id_0;
	wire _mesh_2_6_io_out_last_0;
	wire _mesh_2_6_io_out_valid_0;
	wire [31:0] _mesh_2_5_io_out_a_0;
	wire [31:0] _mesh_2_5_io_out_c_0;
	wire [31:0] _mesh_2_5_io_out_b_0;
	wire _mesh_2_5_io_out_control_0_dataflow;
	wire _mesh_2_5_io_out_control_0_propagate;
	wire [4:0] _mesh_2_5_io_out_control_0_shift;
	wire [2:0] _mesh_2_5_io_out_id_0;
	wire _mesh_2_5_io_out_last_0;
	wire _mesh_2_5_io_out_valid_0;
	wire [31:0] _mesh_2_4_io_out_a_0;
	wire [31:0] _mesh_2_4_io_out_c_0;
	wire [31:0] _mesh_2_4_io_out_b_0;
	wire _mesh_2_4_io_out_control_0_dataflow;
	wire _mesh_2_4_io_out_control_0_propagate;
	wire [4:0] _mesh_2_4_io_out_control_0_shift;
	wire [2:0] _mesh_2_4_io_out_id_0;
	wire _mesh_2_4_io_out_last_0;
	wire _mesh_2_4_io_out_valid_0;
	wire [31:0] _mesh_2_3_io_out_a_0;
	wire [31:0] _mesh_2_3_io_out_c_0;
	wire [31:0] _mesh_2_3_io_out_b_0;
	wire _mesh_2_3_io_out_control_0_dataflow;
	wire _mesh_2_3_io_out_control_0_propagate;
	wire [4:0] _mesh_2_3_io_out_control_0_shift;
	wire [2:0] _mesh_2_3_io_out_id_0;
	wire _mesh_2_3_io_out_last_0;
	wire _mesh_2_3_io_out_valid_0;
	wire [31:0] _mesh_2_2_io_out_a_0;
	wire [31:0] _mesh_2_2_io_out_c_0;
	wire [31:0] _mesh_2_2_io_out_b_0;
	wire _mesh_2_2_io_out_control_0_dataflow;
	wire _mesh_2_2_io_out_control_0_propagate;
	wire [4:0] _mesh_2_2_io_out_control_0_shift;
	wire [2:0] _mesh_2_2_io_out_id_0;
	wire _mesh_2_2_io_out_last_0;
	wire _mesh_2_2_io_out_valid_0;
	wire [31:0] _mesh_2_1_io_out_a_0;
	wire [31:0] _mesh_2_1_io_out_c_0;
	wire [31:0] _mesh_2_1_io_out_b_0;
	wire _mesh_2_1_io_out_control_0_dataflow;
	wire _mesh_2_1_io_out_control_0_propagate;
	wire [4:0] _mesh_2_1_io_out_control_0_shift;
	wire [2:0] _mesh_2_1_io_out_id_0;
	wire _mesh_2_1_io_out_last_0;
	wire _mesh_2_1_io_out_valid_0;
	wire [31:0] _mesh_2_0_io_out_a_0;
	wire [31:0] _mesh_2_0_io_out_c_0;
	wire [31:0] _mesh_2_0_io_out_b_0;
	wire _mesh_2_0_io_out_control_0_dataflow;
	wire _mesh_2_0_io_out_control_0_propagate;
	wire [4:0] _mesh_2_0_io_out_control_0_shift;
	wire [2:0] _mesh_2_0_io_out_id_0;
	wire _mesh_2_0_io_out_last_0;
	wire _mesh_2_0_io_out_valid_0;
	wire [31:0] _mesh_1_7_io_out_a_0;
	wire [31:0] _mesh_1_7_io_out_c_0;
	wire [31:0] _mesh_1_7_io_out_b_0;
	wire _mesh_1_7_io_out_control_0_dataflow;
	wire _mesh_1_7_io_out_control_0_propagate;
	wire [4:0] _mesh_1_7_io_out_control_0_shift;
	wire [2:0] _mesh_1_7_io_out_id_0;
	wire _mesh_1_7_io_out_last_0;
	wire _mesh_1_7_io_out_valid_0;
	wire [31:0] _mesh_1_6_io_out_a_0;
	wire [31:0] _mesh_1_6_io_out_c_0;
	wire [31:0] _mesh_1_6_io_out_b_0;
	wire _mesh_1_6_io_out_control_0_dataflow;
	wire _mesh_1_6_io_out_control_0_propagate;
	wire [4:0] _mesh_1_6_io_out_control_0_shift;
	wire [2:0] _mesh_1_6_io_out_id_0;
	wire _mesh_1_6_io_out_last_0;
	wire _mesh_1_6_io_out_valid_0;
	wire [31:0] _mesh_1_5_io_out_a_0;
	wire [31:0] _mesh_1_5_io_out_c_0;
	wire [31:0] _mesh_1_5_io_out_b_0;
	wire _mesh_1_5_io_out_control_0_dataflow;
	wire _mesh_1_5_io_out_control_0_propagate;
	wire [4:0] _mesh_1_5_io_out_control_0_shift;
	wire [2:0] _mesh_1_5_io_out_id_0;
	wire _mesh_1_5_io_out_last_0;
	wire _mesh_1_5_io_out_valid_0;
	wire [31:0] _mesh_1_4_io_out_a_0;
	wire [31:0] _mesh_1_4_io_out_c_0;
	wire [31:0] _mesh_1_4_io_out_b_0;
	wire _mesh_1_4_io_out_control_0_dataflow;
	wire _mesh_1_4_io_out_control_0_propagate;
	wire [4:0] _mesh_1_4_io_out_control_0_shift;
	wire [2:0] _mesh_1_4_io_out_id_0;
	wire _mesh_1_4_io_out_last_0;
	wire _mesh_1_4_io_out_valid_0;
	wire [31:0] _mesh_1_3_io_out_a_0;
	wire [31:0] _mesh_1_3_io_out_c_0;
	wire [31:0] _mesh_1_3_io_out_b_0;
	wire _mesh_1_3_io_out_control_0_dataflow;
	wire _mesh_1_3_io_out_control_0_propagate;
	wire [4:0] _mesh_1_3_io_out_control_0_shift;
	wire [2:0] _mesh_1_3_io_out_id_0;
	wire _mesh_1_3_io_out_last_0;
	wire _mesh_1_3_io_out_valid_0;
	wire [31:0] _mesh_1_2_io_out_a_0;
	wire [31:0] _mesh_1_2_io_out_c_0;
	wire [31:0] _mesh_1_2_io_out_b_0;
	wire _mesh_1_2_io_out_control_0_dataflow;
	wire _mesh_1_2_io_out_control_0_propagate;
	wire [4:0] _mesh_1_2_io_out_control_0_shift;
	wire [2:0] _mesh_1_2_io_out_id_0;
	wire _mesh_1_2_io_out_last_0;
	wire _mesh_1_2_io_out_valid_0;
	wire [31:0] _mesh_1_1_io_out_a_0;
	wire [31:0] _mesh_1_1_io_out_c_0;
	wire [31:0] _mesh_1_1_io_out_b_0;
	wire _mesh_1_1_io_out_control_0_dataflow;
	wire _mesh_1_1_io_out_control_0_propagate;
	wire [4:0] _mesh_1_1_io_out_control_0_shift;
	wire [2:0] _mesh_1_1_io_out_id_0;
	wire _mesh_1_1_io_out_last_0;
	wire _mesh_1_1_io_out_valid_0;
	wire [31:0] _mesh_1_0_io_out_a_0;
	wire [31:0] _mesh_1_0_io_out_c_0;
	wire [31:0] _mesh_1_0_io_out_b_0;
	wire _mesh_1_0_io_out_control_0_dataflow;
	wire _mesh_1_0_io_out_control_0_propagate;
	wire [4:0] _mesh_1_0_io_out_control_0_shift;
	wire [2:0] _mesh_1_0_io_out_id_0;
	wire _mesh_1_0_io_out_last_0;
	wire _mesh_1_0_io_out_valid_0;
	wire [31:0] _mesh_0_7_io_out_a_0;
	wire [31:0] _mesh_0_7_io_out_c_0;
	wire [31:0] _mesh_0_7_io_out_b_0;
	wire _mesh_0_7_io_out_control_0_dataflow;
	wire _mesh_0_7_io_out_control_0_propagate;
	wire [4:0] _mesh_0_7_io_out_control_0_shift;
	wire [2:0] _mesh_0_7_io_out_id_0;
	wire _mesh_0_7_io_out_last_0;
	wire _mesh_0_7_io_out_valid_0;
	wire [31:0] _mesh_0_6_io_out_a_0;
	wire [31:0] _mesh_0_6_io_out_c_0;
	wire [31:0] _mesh_0_6_io_out_b_0;
	wire _mesh_0_6_io_out_control_0_dataflow;
	wire _mesh_0_6_io_out_control_0_propagate;
	wire [4:0] _mesh_0_6_io_out_control_0_shift;
	wire [2:0] _mesh_0_6_io_out_id_0;
	wire _mesh_0_6_io_out_last_0;
	wire _mesh_0_6_io_out_valid_0;
	wire [31:0] _mesh_0_5_io_out_a_0;
	wire [31:0] _mesh_0_5_io_out_c_0;
	wire [31:0] _mesh_0_5_io_out_b_0;
	wire _mesh_0_5_io_out_control_0_dataflow;
	wire _mesh_0_5_io_out_control_0_propagate;
	wire [4:0] _mesh_0_5_io_out_control_0_shift;
	wire [2:0] _mesh_0_5_io_out_id_0;
	wire _mesh_0_5_io_out_last_0;
	wire _mesh_0_5_io_out_valid_0;
	wire [31:0] _mesh_0_4_io_out_a_0;
	wire [31:0] _mesh_0_4_io_out_c_0;
	wire [31:0] _mesh_0_4_io_out_b_0;
	wire _mesh_0_4_io_out_control_0_dataflow;
	wire _mesh_0_4_io_out_control_0_propagate;
	wire [4:0] _mesh_0_4_io_out_control_0_shift;
	wire [2:0] _mesh_0_4_io_out_id_0;
	wire _mesh_0_4_io_out_last_0;
	wire _mesh_0_4_io_out_valid_0;
	wire [31:0] _mesh_0_3_io_out_a_0;
	wire [31:0] _mesh_0_3_io_out_c_0;
	wire [31:0] _mesh_0_3_io_out_b_0;
	wire _mesh_0_3_io_out_control_0_dataflow;
	wire _mesh_0_3_io_out_control_0_propagate;
	wire [4:0] _mesh_0_3_io_out_control_0_shift;
	wire [2:0] _mesh_0_3_io_out_id_0;
	wire _mesh_0_3_io_out_last_0;
	wire _mesh_0_3_io_out_valid_0;
	wire [31:0] _mesh_0_2_io_out_a_0;
	wire [31:0] _mesh_0_2_io_out_c_0;
	wire [31:0] _mesh_0_2_io_out_b_0;
	wire _mesh_0_2_io_out_control_0_dataflow;
	wire _mesh_0_2_io_out_control_0_propagate;
	wire [4:0] _mesh_0_2_io_out_control_0_shift;
	wire [2:0] _mesh_0_2_io_out_id_0;
	wire _mesh_0_2_io_out_last_0;
	wire _mesh_0_2_io_out_valid_0;
	wire [31:0] _mesh_0_1_io_out_a_0;
	wire [31:0] _mesh_0_1_io_out_c_0;
	wire [31:0] _mesh_0_1_io_out_b_0;
	wire _mesh_0_1_io_out_control_0_dataflow;
	wire _mesh_0_1_io_out_control_0_propagate;
	wire [4:0] _mesh_0_1_io_out_control_0_shift;
	wire [2:0] _mesh_0_1_io_out_id_0;
	wire _mesh_0_1_io_out_last_0;
	wire _mesh_0_1_io_out_valid_0;
	wire [31:0] _mesh_0_0_io_out_a_0;
	wire [31:0] _mesh_0_0_io_out_c_0;
	wire [31:0] _mesh_0_0_io_out_b_0;
	wire _mesh_0_0_io_out_control_0_dataflow;
	wire _mesh_0_0_io_out_control_0_propagate;
	wire [4:0] _mesh_0_0_io_out_control_0_shift;
	wire [2:0] _mesh_0_0_io_out_id_0;
	wire _mesh_0_0_io_out_last_0;
	wire _mesh_0_0_io_out_valid_0;
	reg [31:0] r_0;
	reg [31:0] r_1_0;
	reg [31:0] r_2_0;
	reg [31:0] r_3_0;
	reg [31:0] r_4_0;
	reg [31:0] r_5_0;
	reg [31:0] r_6_0;
	reg [31:0] r_7_0;
	reg [31:0] r_8_0;
	reg [31:0] r_9_0;
	reg [31:0] r_10_0;
	reg [31:0] r_11_0;
	reg [31:0] r_12_0;
	reg [31:0] r_13_0;
	reg [31:0] r_14_0;
	reg [31:0] r_15_0;
	reg [31:0] r_16_0;
	reg [31:0] r_17_0;
	reg [31:0] r_18_0;
	reg [31:0] r_19_0;
	reg [31:0] r_20_0;
	reg [31:0] r_21_0;
	reg [31:0] r_22_0;
	reg [31:0] r_23_0;
	reg [31:0] r_24_0;
	reg [31:0] r_25_0;
	reg [31:0] r_26_0;
	reg [31:0] r_27_0;
	reg [31:0] r_28_0;
	reg [31:0] r_29_0;
	reg [31:0] r_30_0;
	reg [31:0] r_31_0;
	reg [31:0] r_32_0;
	reg [31:0] r_33_0;
	reg [31:0] r_34_0;
	reg [31:0] r_35_0;
	reg [31:0] r_36_0;
	reg [31:0] r_37_0;
	reg [31:0] r_38_0;
	reg [31:0] r_39_0;
	reg [31:0] r_40_0;
	reg [31:0] r_41_0;
	reg [31:0] r_42_0;
	reg [31:0] r_43_0;
	reg [31:0] r_44_0;
	reg [31:0] r_45_0;
	reg [31:0] r_46_0;
	reg [31:0] r_47_0;
	reg [31:0] r_48_0;
	reg [31:0] r_49_0;
	reg [31:0] r_50_0;
	reg [31:0] r_51_0;
	reg [31:0] r_52_0;
	reg [31:0] r_53_0;
	reg [31:0] r_54_0;
	reg [31:0] r_55_0;
	reg [31:0] r_56_0;
	reg [31:0] r_57_0;
	reg [31:0] r_58_0;
	reg [31:0] r_59_0;
	reg [31:0] r_60_0;
	reg [31:0] r_61_0;
	reg [31:0] r_62_0;
	reg [31:0] r_63_0;
	reg [31:0] b_0;
	reg [31:0] b_1_0;
	reg [31:0] b_2_0;
	reg [31:0] b_3_0;
	reg [31:0] b_4_0;
	reg [31:0] b_5_0;
	reg [31:0] b_6_0;
	reg [31:0] b_7_0;
	reg [31:0] b_8_0;
	reg [31:0] b_9_0;
	reg [31:0] b_10_0;
	reg [31:0] b_11_0;
	reg [31:0] b_12_0;
	reg [31:0] b_13_0;
	reg [31:0] b_14_0;
	reg [31:0] b_15_0;
	reg [31:0] b_16_0;
	reg [31:0] b_17_0;
	reg [31:0] b_18_0;
	reg [31:0] b_19_0;
	reg [31:0] b_20_0;
	reg [31:0] b_21_0;
	reg [31:0] b_22_0;
	reg [31:0] b_23_0;
	reg [31:0] b_24_0;
	reg [31:0] b_25_0;
	reg [31:0] b_26_0;
	reg [31:0] b_27_0;
	reg [31:0] b_28_0;
	reg [31:0] b_29_0;
	reg [31:0] b_30_0;
	reg [31:0] b_31_0;
	reg [31:0] b_32_0;
	reg [31:0] b_33_0;
	reg [31:0] b_34_0;
	reg [31:0] b_35_0;
	reg [31:0] b_36_0;
	reg [31:0] b_37_0;
	reg [31:0] b_38_0;
	reg [31:0] b_39_0;
	reg [31:0] b_40_0;
	reg [31:0] b_41_0;
	reg [31:0] b_42_0;
	reg [31:0] b_43_0;
	reg [31:0] b_44_0;
	reg [31:0] b_45_0;
	reg [31:0] b_46_0;
	reg [31:0] b_47_0;
	reg [31:0] b_48_0;
	reg [31:0] b_49_0;
	reg [31:0] b_50_0;
	reg [31:0] b_51_0;
	reg [31:0] b_52_0;
	reg [31:0] b_53_0;
	reg [31:0] b_54_0;
	reg [31:0] b_55_0;
	reg [31:0] b_56_0;
	reg [31:0] b_57_0;
	reg [31:0] b_58_0;
	reg [31:0] b_59_0;
	reg [31:0] b_60_0;
	reg [31:0] b_61_0;
	reg [31:0] b_62_0;
	reg [31:0] b_63_0;
	reg [31:0] b_64_0;
	reg [31:0] b_65_0;
	reg [31:0] b_66_0;
	reg [31:0] b_67_0;
	reg [31:0] b_68_0;
	reg [31:0] b_69_0;
	reg [31:0] b_70_0;
	reg [31:0] b_71_0;
	reg [31:0] b_72_0;
	reg [31:0] b_73_0;
	reg [31:0] b_74_0;
	reg [31:0] b_75_0;
	reg [31:0] b_76_0;
	reg [31:0] b_77_0;
	reg [31:0] b_78_0;
	reg [31:0] b_79_0;
	reg [31:0] b_80_0;
	reg [31:0] b_81_0;
	reg [31:0] b_82_0;
	reg [31:0] b_83_0;
	reg [31:0] b_84_0;
	reg [31:0] b_85_0;
	reg [31:0] b_86_0;
	reg [31:0] b_87_0;
	reg [31:0] b_88_0;
	reg [31:0] b_89_0;
	reg [31:0] b_90_0;
	reg [31:0] b_91_0;
	reg [31:0] b_92_0;
	reg [31:0] b_93_0;
	reg [31:0] b_94_0;
	reg [31:0] b_95_0;
	reg [31:0] b_96_0;
	reg [31:0] b_97_0;
	reg [31:0] b_98_0;
	reg [31:0] b_99_0;
	reg [31:0] b_100_0;
	reg [31:0] b_101_0;
	reg [31:0] b_102_0;
	reg [31:0] b_103_0;
	reg [31:0] b_104_0;
	reg [31:0] b_105_0;
	reg [31:0] b_106_0;
	reg [31:0] b_107_0;
	reg [31:0] b_108_0;
	reg [31:0] b_109_0;
	reg [31:0] b_110_0;
	reg [31:0] b_111_0;
	reg [31:0] b_112_0;
	reg [31:0] b_113_0;
	reg [31:0] b_114_0;
	reg [31:0] b_115_0;
	reg [31:0] b_116_0;
	reg [31:0] b_117_0;
	reg [31:0] b_118_0;
	reg [31:0] b_119_0;
	reg [31:0] b_120_0;
	reg [31:0] b_121_0;
	reg [31:0] b_122_0;
	reg [31:0] b_123_0;
	reg [31:0] b_124_0;
	reg [31:0] b_125_0;
	reg [31:0] b_126_0;
	reg [31:0] b_127_0;
	reg [4:0] mesh_0_0_io_in_control_0_shift_b;
	reg mesh_0_0_io_in_control_0_dataflow_b;
	reg mesh_0_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_0_io_in_control_0_shift_b;
	reg mesh_1_0_io_in_control_0_dataflow_b;
	reg mesh_1_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_0_io_in_control_0_shift_b;
	reg mesh_2_0_io_in_control_0_dataflow_b;
	reg mesh_2_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_0_io_in_control_0_shift_b;
	reg mesh_3_0_io_in_control_0_dataflow_b;
	reg mesh_3_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_0_io_in_control_0_shift_b;
	reg mesh_4_0_io_in_control_0_dataflow_b;
	reg mesh_4_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_0_io_in_control_0_shift_b;
	reg mesh_5_0_io_in_control_0_dataflow_b;
	reg mesh_5_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_0_io_in_control_0_shift_b;
	reg mesh_6_0_io_in_control_0_dataflow_b;
	reg mesh_6_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_0_io_in_control_0_shift_b;
	reg mesh_7_0_io_in_control_0_dataflow_b;
	reg mesh_7_0_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_1_io_in_control_0_shift_b;
	reg mesh_0_1_io_in_control_0_dataflow_b;
	reg mesh_0_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_1_io_in_control_0_shift_b;
	reg mesh_1_1_io_in_control_0_dataflow_b;
	reg mesh_1_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_1_io_in_control_0_shift_b;
	reg mesh_2_1_io_in_control_0_dataflow_b;
	reg mesh_2_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_1_io_in_control_0_shift_b;
	reg mesh_3_1_io_in_control_0_dataflow_b;
	reg mesh_3_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_1_io_in_control_0_shift_b;
	reg mesh_4_1_io_in_control_0_dataflow_b;
	reg mesh_4_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_1_io_in_control_0_shift_b;
	reg mesh_5_1_io_in_control_0_dataflow_b;
	reg mesh_5_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_1_io_in_control_0_shift_b;
	reg mesh_6_1_io_in_control_0_dataflow_b;
	reg mesh_6_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_1_io_in_control_0_shift_b;
	reg mesh_7_1_io_in_control_0_dataflow_b;
	reg mesh_7_1_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_2_io_in_control_0_shift_b;
	reg mesh_0_2_io_in_control_0_dataflow_b;
	reg mesh_0_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_2_io_in_control_0_shift_b;
	reg mesh_1_2_io_in_control_0_dataflow_b;
	reg mesh_1_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_2_io_in_control_0_shift_b;
	reg mesh_2_2_io_in_control_0_dataflow_b;
	reg mesh_2_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_2_io_in_control_0_shift_b;
	reg mesh_3_2_io_in_control_0_dataflow_b;
	reg mesh_3_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_2_io_in_control_0_shift_b;
	reg mesh_4_2_io_in_control_0_dataflow_b;
	reg mesh_4_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_2_io_in_control_0_shift_b;
	reg mesh_5_2_io_in_control_0_dataflow_b;
	reg mesh_5_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_2_io_in_control_0_shift_b;
	reg mesh_6_2_io_in_control_0_dataflow_b;
	reg mesh_6_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_2_io_in_control_0_shift_b;
	reg mesh_7_2_io_in_control_0_dataflow_b;
	reg mesh_7_2_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_3_io_in_control_0_shift_b;
	reg mesh_0_3_io_in_control_0_dataflow_b;
	reg mesh_0_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_3_io_in_control_0_shift_b;
	reg mesh_1_3_io_in_control_0_dataflow_b;
	reg mesh_1_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_3_io_in_control_0_shift_b;
	reg mesh_2_3_io_in_control_0_dataflow_b;
	reg mesh_2_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_3_io_in_control_0_shift_b;
	reg mesh_3_3_io_in_control_0_dataflow_b;
	reg mesh_3_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_3_io_in_control_0_shift_b;
	reg mesh_4_3_io_in_control_0_dataflow_b;
	reg mesh_4_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_3_io_in_control_0_shift_b;
	reg mesh_5_3_io_in_control_0_dataflow_b;
	reg mesh_5_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_3_io_in_control_0_shift_b;
	reg mesh_6_3_io_in_control_0_dataflow_b;
	reg mesh_6_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_3_io_in_control_0_shift_b;
	reg mesh_7_3_io_in_control_0_dataflow_b;
	reg mesh_7_3_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_4_io_in_control_0_shift_b;
	reg mesh_0_4_io_in_control_0_dataflow_b;
	reg mesh_0_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_4_io_in_control_0_shift_b;
	reg mesh_1_4_io_in_control_0_dataflow_b;
	reg mesh_1_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_4_io_in_control_0_shift_b;
	reg mesh_2_4_io_in_control_0_dataflow_b;
	reg mesh_2_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_4_io_in_control_0_shift_b;
	reg mesh_3_4_io_in_control_0_dataflow_b;
	reg mesh_3_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_4_io_in_control_0_shift_b;
	reg mesh_4_4_io_in_control_0_dataflow_b;
	reg mesh_4_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_4_io_in_control_0_shift_b;
	reg mesh_5_4_io_in_control_0_dataflow_b;
	reg mesh_5_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_4_io_in_control_0_shift_b;
	reg mesh_6_4_io_in_control_0_dataflow_b;
	reg mesh_6_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_4_io_in_control_0_shift_b;
	reg mesh_7_4_io_in_control_0_dataflow_b;
	reg mesh_7_4_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_5_io_in_control_0_shift_b;
	reg mesh_0_5_io_in_control_0_dataflow_b;
	reg mesh_0_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_5_io_in_control_0_shift_b;
	reg mesh_1_5_io_in_control_0_dataflow_b;
	reg mesh_1_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_5_io_in_control_0_shift_b;
	reg mesh_2_5_io_in_control_0_dataflow_b;
	reg mesh_2_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_5_io_in_control_0_shift_b;
	reg mesh_3_5_io_in_control_0_dataflow_b;
	reg mesh_3_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_5_io_in_control_0_shift_b;
	reg mesh_4_5_io_in_control_0_dataflow_b;
	reg mesh_4_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_5_io_in_control_0_shift_b;
	reg mesh_5_5_io_in_control_0_dataflow_b;
	reg mesh_5_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_5_io_in_control_0_shift_b;
	reg mesh_6_5_io_in_control_0_dataflow_b;
	reg mesh_6_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_5_io_in_control_0_shift_b;
	reg mesh_7_5_io_in_control_0_dataflow_b;
	reg mesh_7_5_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_6_io_in_control_0_shift_b;
	reg mesh_0_6_io_in_control_0_dataflow_b;
	reg mesh_0_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_6_io_in_control_0_shift_b;
	reg mesh_1_6_io_in_control_0_dataflow_b;
	reg mesh_1_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_6_io_in_control_0_shift_b;
	reg mesh_2_6_io_in_control_0_dataflow_b;
	reg mesh_2_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_6_io_in_control_0_shift_b;
	reg mesh_3_6_io_in_control_0_dataflow_b;
	reg mesh_3_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_6_io_in_control_0_shift_b;
	reg mesh_4_6_io_in_control_0_dataflow_b;
	reg mesh_4_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_6_io_in_control_0_shift_b;
	reg mesh_5_6_io_in_control_0_dataflow_b;
	reg mesh_5_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_6_io_in_control_0_shift_b;
	reg mesh_6_6_io_in_control_0_dataflow_b;
	reg mesh_6_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_6_io_in_control_0_shift_b;
	reg mesh_7_6_io_in_control_0_dataflow_b;
	reg mesh_7_6_io_in_control_0_propagate_b;
	reg [4:0] mesh_0_7_io_in_control_0_shift_b;
	reg mesh_0_7_io_in_control_0_dataflow_b;
	reg mesh_0_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_1_7_io_in_control_0_shift_b;
	reg mesh_1_7_io_in_control_0_dataflow_b;
	reg mesh_1_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_2_7_io_in_control_0_shift_b;
	reg mesh_2_7_io_in_control_0_dataflow_b;
	reg mesh_2_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_3_7_io_in_control_0_shift_b;
	reg mesh_3_7_io_in_control_0_dataflow_b;
	reg mesh_3_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_4_7_io_in_control_0_shift_b;
	reg mesh_4_7_io_in_control_0_dataflow_b;
	reg mesh_4_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_5_7_io_in_control_0_shift_b;
	reg mesh_5_7_io_in_control_0_dataflow_b;
	reg mesh_5_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_6_7_io_in_control_0_shift_b;
	reg mesh_6_7_io_in_control_0_dataflow_b;
	reg mesh_6_7_io_in_control_0_propagate_b;
	reg [4:0] mesh_7_7_io_in_control_0_shift_b;
	reg mesh_7_7_io_in_control_0_dataflow_b;
	reg mesh_7_7_io_in_control_0_propagate_b;
	reg r_64_0;
	reg r_65_0;
	reg r_66_0;
	reg r_67_0;
	reg r_68_0;
	reg r_69_0;
	reg r_70_0;
	reg r_71_0;
	reg r_72_0;
	reg r_73_0;
	reg r_74_0;
	reg r_75_0;
	reg r_76_0;
	reg r_77_0;
	reg r_78_0;
	reg r_79_0;
	reg r_80_0;
	reg r_81_0;
	reg r_82_0;
	reg r_83_0;
	reg r_84_0;
	reg r_85_0;
	reg r_86_0;
	reg r_87_0;
	reg r_88_0;
	reg r_89_0;
	reg r_90_0;
	reg r_91_0;
	reg r_92_0;
	reg r_93_0;
	reg r_94_0;
	reg r_95_0;
	reg r_96_0;
	reg r_97_0;
	reg r_98_0;
	reg r_99_0;
	reg r_100_0;
	reg r_101_0;
	reg r_102_0;
	reg r_103_0;
	reg r_104_0;
	reg r_105_0;
	reg r_106_0;
	reg r_107_0;
	reg r_108_0;
	reg r_109_0;
	reg r_110_0;
	reg r_111_0;
	reg r_112_0;
	reg r_113_0;
	reg r_114_0;
	reg r_115_0;
	reg r_116_0;
	reg r_117_0;
	reg r_118_0;
	reg r_119_0;
	reg r_120_0;
	reg r_121_0;
	reg r_122_0;
	reg r_123_0;
	reg r_124_0;
	reg r_125_0;
	reg r_126_0;
	reg r_127_0;
	reg [2:0] r_128_0;
	reg [2:0] r_129_0;
	reg [2:0] r_130_0;
	reg [2:0] r_131_0;
	reg [2:0] r_132_0;
	reg [2:0] r_133_0;
	reg [2:0] r_134_0;
	reg [2:0] r_135_0;
	reg [2:0] r_136_0;
	reg [2:0] r_137_0;
	reg [2:0] r_138_0;
	reg [2:0] r_139_0;
	reg [2:0] r_140_0;
	reg [2:0] r_141_0;
	reg [2:0] r_142_0;
	reg [2:0] r_143_0;
	reg [2:0] r_144_0;
	reg [2:0] r_145_0;
	reg [2:0] r_146_0;
	reg [2:0] r_147_0;
	reg [2:0] r_148_0;
	reg [2:0] r_149_0;
	reg [2:0] r_150_0;
	reg [2:0] r_151_0;
	reg [2:0] r_152_0;
	reg [2:0] r_153_0;
	reg [2:0] r_154_0;
	reg [2:0] r_155_0;
	reg [2:0] r_156_0;
	reg [2:0] r_157_0;
	reg [2:0] r_158_0;
	reg [2:0] r_159_0;
	reg [2:0] r_160_0;
	reg [2:0] r_161_0;
	reg [2:0] r_162_0;
	reg [2:0] r_163_0;
	reg [2:0] r_164_0;
	reg [2:0] r_165_0;
	reg [2:0] r_166_0;
	reg [2:0] r_167_0;
	reg [2:0] r_168_0;
	reg [2:0] r_169_0;
	reg [2:0] r_170_0;
	reg [2:0] r_171_0;
	reg [2:0] r_172_0;
	reg [2:0] r_173_0;
	reg [2:0] r_174_0;
	reg [2:0] r_175_0;
	reg [2:0] r_176_0;
	reg [2:0] r_177_0;
	reg [2:0] r_178_0;
	reg [2:0] r_179_0;
	reg [2:0] r_180_0;
	reg [2:0] r_181_0;
	reg [2:0] r_182_0;
	reg [2:0] r_183_0;
	reg [2:0] r_184_0;
	reg [2:0] r_185_0;
	reg [2:0] r_186_0;
	reg [2:0] r_187_0;
	reg [2:0] r_188_0;
	reg [2:0] r_189_0;
	reg [2:0] r_190_0;
	reg [2:0] r_191_0;
	reg r_192_0;
	reg r_193_0;
	reg r_194_0;
	reg r_195_0;
	reg r_196_0;
	reg r_197_0;
	reg r_198_0;
	reg r_199_0;
	reg r_200_0;
	reg r_201_0;
	reg r_202_0;
	reg r_203_0;
	reg r_204_0;
	reg r_205_0;
	reg r_206_0;
	reg r_207_0;
	reg r_208_0;
	reg r_209_0;
	reg r_210_0;
	reg r_211_0;
	reg r_212_0;
	reg r_213_0;
	reg r_214_0;
	reg r_215_0;
	reg r_216_0;
	reg r_217_0;
	reg r_218_0;
	reg r_219_0;
	reg r_220_0;
	reg r_221_0;
	reg r_222_0;
	reg r_223_0;
	reg r_224_0;
	reg r_225_0;
	reg r_226_0;
	reg r_227_0;
	reg r_228_0;
	reg r_229_0;
	reg r_230_0;
	reg r_231_0;
	reg r_232_0;
	reg r_233_0;
	reg r_234_0;
	reg r_235_0;
	reg r_236_0;
	reg r_237_0;
	reg r_238_0;
	reg r_239_0;
	reg r_240_0;
	reg r_241_0;
	reg r_242_0;
	reg r_243_0;
	reg r_244_0;
	reg r_245_0;
	reg r_246_0;
	reg r_247_0;
	reg r_248_0;
	reg r_249_0;
	reg r_250_0;
	reg r_251_0;
	reg r_252_0;
	reg r_253_0;
	reg r_254_0;
	reg r_255_0;
	reg [31:0] r_256_0;
	reg [31:0] r_257_0;
	reg r_258_0;
	reg r_259_0_dataflow;
	reg [2:0] r_260_0;
	reg r_261_0;
	reg [31:0] r_262_0;
	reg [31:0] r_263_0;
	reg [31:0] r_268_0;
	reg [31:0] r_269_0;
	reg [31:0] r_274_0;
	reg [31:0] r_275_0;
	reg [31:0] r_280_0;
	reg [31:0] r_281_0;
	reg [31:0] r_286_0;
	reg [31:0] r_287_0;
	reg [31:0] r_292_0;
	reg [31:0] r_293_0;
	reg [31:0] r_298_0;
	reg [31:0] r_299_0;
	always @(posedge clock) begin
		r_0 <=( io_in_a_0_0) ^ ((fiEnable && (17 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_1_0 <=( _mesh_0_0_io_out_a_0) ^ ((fiEnable && (18 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_2_0 <=( _mesh_0_1_io_out_a_0) ^ ((fiEnable && (19 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_3_0 <=( _mesh_0_2_io_out_a_0) ^ ((fiEnable && (20 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_4_0 <=( _mesh_0_3_io_out_a_0) ^ ((fiEnable && (21 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_5_0 <=( _mesh_0_4_io_out_a_0) ^ ((fiEnable && (22 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_6_0 <=( _mesh_0_5_io_out_a_0) ^ ((fiEnable && (23 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_7_0 <=( _mesh_0_6_io_out_a_0) ^ ((fiEnable && (24 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_8_0 <=( io_in_a_1_0) ^ ((fiEnable && (25 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_9_0 <=( _mesh_1_0_io_out_a_0) ^ ((fiEnable && (26 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_10_0 <=( _mesh_1_1_io_out_a_0) ^ ((fiEnable && (27 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_11_0 <=( _mesh_1_2_io_out_a_0) ^ ((fiEnable && (28 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_12_0 <=( _mesh_1_3_io_out_a_0) ^ ((fiEnable && (29 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_13_0 <=( _mesh_1_4_io_out_a_0) ^ ((fiEnable && (30 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_14_0 <=( _mesh_1_5_io_out_a_0) ^ ((fiEnable && (31 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_15_0 <=( _mesh_1_6_io_out_a_0) ^ ((fiEnable && (32 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_16_0 <=( io_in_a_2_0) ^ ((fiEnable && (33 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_17_0 <=( _mesh_2_0_io_out_a_0) ^ ((fiEnable && (34 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_18_0 <=( _mesh_2_1_io_out_a_0) ^ ((fiEnable && (35 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_19_0 <=( _mesh_2_2_io_out_a_0) ^ ((fiEnable && (36 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_20_0 <=( _mesh_2_3_io_out_a_0) ^ ((fiEnable && (37 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_21_0 <=( _mesh_2_4_io_out_a_0) ^ ((fiEnable && (38 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_22_0 <=( _mesh_2_5_io_out_a_0) ^ ((fiEnable && (39 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_23_0 <=( _mesh_2_6_io_out_a_0) ^ ((fiEnable && (40 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_24_0 <=( io_in_a_3_0) ^ ((fiEnable && (41 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_25_0 <=( _mesh_3_0_io_out_a_0) ^ ((fiEnable && (42 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_26_0 <=( _mesh_3_1_io_out_a_0) ^ ((fiEnable && (43 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_27_0 <=( _mesh_3_2_io_out_a_0) ^ ((fiEnable && (44 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_28_0 <=( _mesh_3_3_io_out_a_0) ^ ((fiEnable && (45 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_29_0 <=( _mesh_3_4_io_out_a_0) ^ ((fiEnable && (46 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_30_0 <=( _mesh_3_5_io_out_a_0) ^ ((fiEnable && (47 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_31_0 <=( _mesh_3_6_io_out_a_0) ^ ((fiEnable && (48 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_32_0 <=( io_in_a_4_0) ^ ((fiEnable && (49 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_33_0 <=( _mesh_4_0_io_out_a_0) ^ ((fiEnable && (50 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_34_0 <=( _mesh_4_1_io_out_a_0) ^ ((fiEnable && (51 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_35_0 <=( _mesh_4_2_io_out_a_0) ^ ((fiEnable && (52 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_36_0 <=( _mesh_4_3_io_out_a_0) ^ ((fiEnable && (53 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_37_0 <=( _mesh_4_4_io_out_a_0) ^ ((fiEnable && (54 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_38_0 <=( _mesh_4_5_io_out_a_0) ^ ((fiEnable && (55 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_39_0 <=( _mesh_4_6_io_out_a_0) ^ ((fiEnable && (56 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_40_0 <=( io_in_a_5_0) ^ ((fiEnable && (57 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_41_0 <=( _mesh_5_0_io_out_a_0) ^ ((fiEnable && (58 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_42_0 <=( _mesh_5_1_io_out_a_0) ^ ((fiEnable && (59 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_43_0 <=( _mesh_5_2_io_out_a_0) ^ ((fiEnable && (60 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_44_0 <=( _mesh_5_3_io_out_a_0) ^ ((fiEnable && (61 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_45_0 <=( _mesh_5_4_io_out_a_0) ^ ((fiEnable && (62 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_46_0 <=( _mesh_5_5_io_out_a_0) ^ ((fiEnable && (63 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_47_0 <=( _mesh_5_6_io_out_a_0) ^ ((fiEnable && (64 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_48_0 <=( io_in_a_6_0) ^ ((fiEnable && (65 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_49_0 <=( _mesh_6_0_io_out_a_0) ^ ((fiEnable && (66 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_50_0 <=( _mesh_6_1_io_out_a_0) ^ ((fiEnable && (67 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_51_0 <=( _mesh_6_2_io_out_a_0) ^ ((fiEnable && (68 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_52_0 <=( _mesh_6_3_io_out_a_0) ^ ((fiEnable && (69 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_53_0 <=( _mesh_6_4_io_out_a_0) ^ ((fiEnable && (70 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_54_0 <=( _mesh_6_5_io_out_a_0) ^ ((fiEnable && (71 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_55_0 <=( _mesh_6_6_io_out_a_0) ^ ((fiEnable && (72 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_56_0 <=( io_in_a_7_0) ^ ((fiEnable && (73 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_57_0 <=( _mesh_7_0_io_out_a_0) ^ ((fiEnable && (74 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_58_0 <=( _mesh_7_1_io_out_a_0) ^ ((fiEnable && (75 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_59_0 <=( _mesh_7_2_io_out_a_0) ^ ((fiEnable && (76 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_60_0 <=( _mesh_7_3_io_out_a_0) ^ ((fiEnable && (77 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_61_0 <=( _mesh_7_4_io_out_a_0) ^ ((fiEnable && (78 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_62_0 <=( _mesh_7_5_io_out_a_0) ^ ((fiEnable && (79 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_63_0 <=( _mesh_7_6_io_out_a_0) ^ ((fiEnable && (80 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		if (io_in_valid_0_0) begin
			b_0 <=( io_in_b_0_0) ^ ((fiEnable && (81 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_64_0 <=( io_in_d_0_0) ^ ((fiEnable && (82 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_0_io_in_control_0_shift_b <=( io_in_control_0_0_shift) ^ ((fiEnable && (83 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_0_io_in_control_0_dataflow_b <=( io_in_control_0_0_dataflow) ^ ((fiEnable && (84 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_0_io_in_control_0_propagate_b <=( io_in_control_0_0_propagate) ^ ((fiEnable && (85 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_0_io_out_valid_0) begin 
			b_1_0 <=( _mesh_0_0_io_out_b_0) ^ ((fiEnable && (86 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_65_0 <=( _mesh_0_0_io_out_c_0) ^ ((fiEnable && (87 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_0_io_in_control_0_shift_b <=( _mesh_0_0_io_out_control_0_shift) ^ ((fiEnable && (88 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_0_io_in_control_0_dataflow_b <=( _mesh_0_0_io_out_control_0_dataflow) ^ ((fiEnable && (89 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_0_io_in_control_0_propagate_b <=( _mesh_0_0_io_out_control_0_propagate) ^ ((fiEnable && (90 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_0_io_out_valid_0) begin
			b_2_0 <=( _mesh_1_0_io_out_b_0) ^ ((fiEnable && (91 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_66_0 <=( _mesh_1_0_io_out_c_0) ^ ((fiEnable && (92 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_0_io_in_control_0_shift_b <=( _mesh_1_0_io_out_control_0_shift) ^ ((fiEnable && (93 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_0_io_in_control_0_dataflow_b <=( _mesh_1_0_io_out_control_0_dataflow) ^ ((fiEnable && (94 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_0_io_in_control_0_propagate_b <=( _mesh_1_0_io_out_control_0_propagate) ^ ((fiEnable && (95 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_0_io_out_valid_0) begin
			b_3_0 <=( _mesh_2_0_io_out_b_0) ^ ((fiEnable && (96 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_67_0 <=( _mesh_2_0_io_out_c_0) ^ ((fiEnable && (97 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_0_io_in_control_0_shift_b <=( _mesh_2_0_io_out_control_0_shift) ^ ((fiEnable && (98 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_0_io_in_control_0_dataflow_b <=( _mesh_2_0_io_out_control_0_dataflow) ^ ((fiEnable && (99 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_0_io_in_control_0_propagate_b <=( _mesh_2_0_io_out_control_0_propagate) ^ ((fiEnable && (100 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_0_io_out_valid_0) begin
			b_4_0 <=( _mesh_3_0_io_out_b_0) ^ ((fiEnable && (101 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_68_0 <=( _mesh_3_0_io_out_c_0) ^ ((fiEnable && (102 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_0_io_in_control_0_shift_b <=( _mesh_3_0_io_out_control_0_shift) ^ ((fiEnable && (103 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_0_io_in_control_0_dataflow_b <=( _mesh_3_0_io_out_control_0_dataflow) ^ ((fiEnable && (104 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_0_io_in_control_0_propagate_b <=( _mesh_3_0_io_out_control_0_propagate) ^ ((fiEnable && (105 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_0_io_out_valid_0) begin
			b_5_0 <=( _mesh_4_0_io_out_b_0) ^ ((fiEnable && (106 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_69_0 <=( _mesh_4_0_io_out_c_0) ^ ((fiEnable && (107 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_0_io_in_control_0_shift_b <=( _mesh_4_0_io_out_control_0_shift) ^ ((fiEnable && (108 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_0_io_in_control_0_dataflow_b <=( _mesh_4_0_io_out_control_0_dataflow) ^ ((fiEnable && (109 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_0_io_in_control_0_propagate_b <=( _mesh_4_0_io_out_control_0_propagate) ^ ((fiEnable && (110 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_0_io_out_valid_0) begin
			b_6_0 <=( _mesh_5_0_io_out_b_0) ^ ((fiEnable && (111 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_70_0 <=( _mesh_5_0_io_out_c_0) ^ ((fiEnable && (112 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_0_io_in_control_0_shift_b <=( _mesh_5_0_io_out_control_0_shift) ^ ((fiEnable && (113 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_0_io_in_control_0_dataflow_b <=( _mesh_5_0_io_out_control_0_dataflow) ^ ((fiEnable && (114 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_0_io_in_control_0_propagate_b <=( _mesh_5_0_io_out_control_0_propagate) ^ ((fiEnable && (115 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_0_io_out_valid_0) begin
			b_7_0 <=( _mesh_6_0_io_out_b_0) ^ ((fiEnable && (116 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_71_0 <=( _mesh_6_0_io_out_c_0) ^ ((fiEnable && (117 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_0_io_in_control_0_shift_b <=( _mesh_6_0_io_out_control_0_shift) ^ ((fiEnable && (118 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_0_io_in_control_0_dataflow_b <=( _mesh_6_0_io_out_control_0_dataflow) ^ ((fiEnable && (119 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_0_io_in_control_0_propagate_b <=( _mesh_6_0_io_out_control_0_propagate) ^ ((fiEnable && (120 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_1_0) begin
			b_8_0 <=( io_in_b_1_0) ^ ((fiEnable && (121 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_72_0 <=( io_in_d_1_0) ^ ((fiEnable && (122 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_1_io_in_control_0_shift_b <=( io_in_control_1_0_shift) ^ ((fiEnable && (123 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_1_io_in_control_0_dataflow_b <=( io_in_control_1_0_dataflow) ^ ((fiEnable && (124 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_1_io_in_control_0_propagate_b <=( io_in_control_1_0_propagate) ^ ((fiEnable && (125 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_1_io_out_valid_0) begin
			b_9_0 <=( _mesh_0_1_io_out_b_0) ^ ((fiEnable && (126 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_73_0 <=( _mesh_0_1_io_out_c_0) ^ ((fiEnable && (127 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_1_io_in_control_0_shift_b <=( _mesh_0_1_io_out_control_0_shift) ^ ((fiEnable && (128 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_1_io_in_control_0_dataflow_b <=( _mesh_0_1_io_out_control_0_dataflow) ^ ((fiEnable && (129 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_1_io_in_control_0_propagate_b <=( _mesh_0_1_io_out_control_0_propagate) ^ ((fiEnable && (130 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_1_io_out_valid_0) begin
			b_10_0 <=( _mesh_1_1_io_out_b_0) ^ ((fiEnable && (131 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_74_0 <=( _mesh_1_1_io_out_c_0) ^ ((fiEnable && (132 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_1_io_in_control_0_shift_b <=( _mesh_1_1_io_out_control_0_shift) ^ ((fiEnable && (133 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_1_io_in_control_0_dataflow_b <=( _mesh_1_1_io_out_control_0_dataflow) ^ ((fiEnable && (134 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_1_io_in_control_0_propagate_b <=( _mesh_1_1_io_out_control_0_propagate) ^ ((fiEnable && (135 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_1_io_out_valid_0) begin
			b_11_0 <=( _mesh_2_1_io_out_b_0) ^ ((fiEnable && (136 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_75_0 <=( _mesh_2_1_io_out_c_0) ^ ((fiEnable && (137 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_1_io_in_control_0_shift_b <=( _mesh_2_1_io_out_control_0_shift) ^ ((fiEnable && (138 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_1_io_in_control_0_dataflow_b <=( _mesh_2_1_io_out_control_0_dataflow) ^ ((fiEnable && (139 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_1_io_in_control_0_propagate_b <=( _mesh_2_1_io_out_control_0_propagate) ^ ((fiEnable && (140 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_1_io_out_valid_0) begin
			b_12_0 <=( _mesh_3_1_io_out_b_0) ^ ((fiEnable && (141 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_76_0 <=( _mesh_3_1_io_out_c_0) ^ ((fiEnable && (142 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_1_io_in_control_0_shift_b <=( _mesh_3_1_io_out_control_0_shift) ^ ((fiEnable && (143 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_1_io_in_control_0_dataflow_b <=( _mesh_3_1_io_out_control_0_dataflow) ^ ((fiEnable && (144 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_1_io_in_control_0_propagate_b <=( _mesh_3_1_io_out_control_0_propagate) ^ ((fiEnable && (145 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_1_io_out_valid_0) begin
			b_13_0 <=( _mesh_4_1_io_out_b_0) ^ ((fiEnable && (146 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_77_0 <=( _mesh_4_1_io_out_c_0) ^ ((fiEnable && (147 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_1_io_in_control_0_shift_b <=( _mesh_4_1_io_out_control_0_shift) ^ ((fiEnable && (148 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_1_io_in_control_0_dataflow_b <=( _mesh_4_1_io_out_control_0_dataflow) ^ ((fiEnable && (149 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_1_io_in_control_0_propagate_b <=( _mesh_4_1_io_out_control_0_propagate) ^ ((fiEnable && (150 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_1_io_out_valid_0) begin
			b_14_0 <=( _mesh_5_1_io_out_b_0) ^ ((fiEnable && (151 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_78_0 <=( _mesh_5_1_io_out_c_0) ^ ((fiEnable && (152 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_1_io_in_control_0_shift_b <=( _mesh_5_1_io_out_control_0_shift) ^ ((fiEnable && (153 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_1_io_in_control_0_dataflow_b <=( _mesh_5_1_io_out_control_0_dataflow) ^ ((fiEnable && (154 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_1_io_in_control_0_propagate_b <=( _mesh_5_1_io_out_control_0_propagate) ^ ((fiEnable && (155 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_1_io_out_valid_0) begin
			b_15_0 <=( _mesh_6_1_io_out_b_0) ^ ((fiEnable && (156 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_79_0 <=( _mesh_6_1_io_out_c_0) ^ ((fiEnable && (157 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_1_io_in_control_0_shift_b <=( _mesh_6_1_io_out_control_0_shift) ^ ((fiEnable && (158 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_1_io_in_control_0_dataflow_b <=( _mesh_6_1_io_out_control_0_dataflow) ^ ((fiEnable && (159 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_1_io_in_control_0_propagate_b <=( _mesh_6_1_io_out_control_0_propagate) ^ ((fiEnable && (160 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_2_0) begin
			b_16_0 <=( io_in_b_2_0) ^ ((fiEnable && (161 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_80_0 <=( io_in_d_2_0) ^ ((fiEnable && (162 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_2_io_in_control_0_shift_b <=( io_in_control_2_0_shift) ^ ((fiEnable && (163 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_2_io_in_control_0_dataflow_b <=( io_in_control_2_0_dataflow) ^ ((fiEnable && (164 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_2_io_in_control_0_propagate_b <=( io_in_control_2_0_propagate) ^ ((fiEnable && (165 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_2_io_out_valid_0) begin
			b_17_0 <=( _mesh_0_2_io_out_b_0) ^ ((fiEnable && (166 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_81_0 <=( _mesh_0_2_io_out_c_0) ^ ((fiEnable && (167 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_2_io_in_control_0_shift_b <=( _mesh_0_2_io_out_control_0_shift) ^ ((fiEnable && (168 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_2_io_in_control_0_dataflow_b <=( _mesh_0_2_io_out_control_0_dataflow) ^ ((fiEnable && (169 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_2_io_in_control_0_propagate_b <=( _mesh_0_2_io_out_control_0_propagate) ^ ((fiEnable && (170 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_2_io_out_valid_0) begin
			b_18_0 <=( _mesh_1_2_io_out_b_0) ^ ((fiEnable && (171 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_82_0 <=( _mesh_1_2_io_out_c_0) ^ ((fiEnable && (172 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_2_io_in_control_0_shift_b <=( _mesh_1_2_io_out_control_0_shift) ^ ((fiEnable && (173 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_2_io_in_control_0_dataflow_b <=( _mesh_1_2_io_out_control_0_dataflow) ^ ((fiEnable && (174 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_2_io_in_control_0_propagate_b <=( _mesh_1_2_io_out_control_0_propagate) ^ ((fiEnable && (175 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_2_io_out_valid_0) begin
			b_19_0 <=( _mesh_2_2_io_out_b_0) ^ ((fiEnable && (176 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_83_0 <=( _mesh_2_2_io_out_c_0) ^ ((fiEnable && (177 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_2_io_in_control_0_shift_b <=( _mesh_2_2_io_out_control_0_shift) ^ ((fiEnable && (178 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_2_io_in_control_0_dataflow_b <=( _mesh_2_2_io_out_control_0_dataflow) ^ ((fiEnable && (179 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_2_io_in_control_0_propagate_b <=( _mesh_2_2_io_out_control_0_propagate) ^ ((fiEnable && (180 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_2_io_out_valid_0) begin
			b_20_0 <=( _mesh_3_2_io_out_b_0) ^ ((fiEnable && (181 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_84_0 <=( _mesh_3_2_io_out_c_0) ^ ((fiEnable && (182 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_2_io_in_control_0_shift_b <=( _mesh_3_2_io_out_control_0_shift) ^ ((fiEnable && (183 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_2_io_in_control_0_dataflow_b <=( _mesh_3_2_io_out_control_0_dataflow) ^ ((fiEnable && (184 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_2_io_in_control_0_propagate_b <=( _mesh_3_2_io_out_control_0_propagate) ^ ((fiEnable && (185 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_2_io_out_valid_0) begin
			b_21_0 <=( _mesh_4_2_io_out_b_0) ^ ((fiEnable && (186 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_85_0 <=( _mesh_4_2_io_out_c_0) ^ ((fiEnable && (187 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_2_io_in_control_0_shift_b <=( _mesh_4_2_io_out_control_0_shift) ^ ((fiEnable && (188 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_2_io_in_control_0_dataflow_b <=( _mesh_4_2_io_out_control_0_dataflow) ^ ((fiEnable && (189 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_2_io_in_control_0_propagate_b <=( _mesh_4_2_io_out_control_0_propagate) ^ ((fiEnable && (190 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_2_io_out_valid_0) begin
			b_22_0 <=( _mesh_5_2_io_out_b_0) ^ ((fiEnable && (191 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_86_0 <=( _mesh_5_2_io_out_c_0) ^ ((fiEnable && (192 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_2_io_in_control_0_shift_b <=( _mesh_5_2_io_out_control_0_shift) ^ ((fiEnable && (193 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_2_io_in_control_0_dataflow_b <=( _mesh_5_2_io_out_control_0_dataflow) ^ ((fiEnable && (194 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_2_io_in_control_0_propagate_b <=( _mesh_5_2_io_out_control_0_propagate) ^ ((fiEnable && (195 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_2_io_out_valid_0) begin
			b_23_0 <=( _mesh_6_2_io_out_b_0) ^ ((fiEnable && (196 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_87_0 <=( _mesh_6_2_io_out_c_0) ^ ((fiEnable && (197 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_2_io_in_control_0_shift_b <=( _mesh_6_2_io_out_control_0_shift) ^ ((fiEnable && (198 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_2_io_in_control_0_dataflow_b <=( _mesh_6_2_io_out_control_0_dataflow) ^ ((fiEnable && (199 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_2_io_in_control_0_propagate_b <=( _mesh_6_2_io_out_control_0_propagate) ^ ((fiEnable && (200 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_3_0) begin
			b_24_0 <=( io_in_b_3_0) ^ ((fiEnable && (201 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_88_0 <=( io_in_d_3_0) ^ ((fiEnable && (202 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_3_io_in_control_0_shift_b <=( io_in_control_3_0_shift) ^ ((fiEnable && (203 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_3_io_in_control_0_dataflow_b <=( io_in_control_3_0_dataflow) ^ ((fiEnable && (204 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_3_io_in_control_0_propagate_b <=( io_in_control_3_0_propagate) ^ ((fiEnable && (205 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_3_io_out_valid_0) begin
			b_25_0 <=( _mesh_0_3_io_out_b_0) ^ ((fiEnable && (206 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_89_0 <=( _mesh_0_3_io_out_c_0) ^ ((fiEnable && (207 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_3_io_in_control_0_shift_b <=( _mesh_0_3_io_out_control_0_shift) ^ ((fiEnable && (208 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_3_io_in_control_0_dataflow_b <=( _mesh_0_3_io_out_control_0_dataflow) ^ ((fiEnable && (209 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_3_io_in_control_0_propagate_b <=( _mesh_0_3_io_out_control_0_propagate) ^ ((fiEnable && (210 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_3_io_out_valid_0) begin
			b_26_0 <=( _mesh_1_3_io_out_b_0) ^ ((fiEnable && (211 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_90_0 <=( _mesh_1_3_io_out_c_0) ^ ((fiEnable && (212 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_3_io_in_control_0_shift_b <=( _mesh_1_3_io_out_control_0_shift) ^ ((fiEnable && (213 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_3_io_in_control_0_dataflow_b <=( _mesh_1_3_io_out_control_0_dataflow) ^ ((fiEnable && (214 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_3_io_in_control_0_propagate_b <=( _mesh_1_3_io_out_control_0_propagate) ^ ((fiEnable && (215 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_3_io_out_valid_0) begin
			b_27_0 <=( _mesh_2_3_io_out_b_0) ^ ((fiEnable && (216 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_91_0 <=( _mesh_2_3_io_out_c_0) ^ ((fiEnable && (217 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_3_io_in_control_0_shift_b <=( _mesh_2_3_io_out_control_0_shift) ^ ((fiEnable && (218 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_3_io_in_control_0_dataflow_b <=( _mesh_2_3_io_out_control_0_dataflow) ^ ((fiEnable && (219 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_3_io_in_control_0_propagate_b <=( _mesh_2_3_io_out_control_0_propagate) ^ ((fiEnable && (220 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_3_io_out_valid_0) begin
			b_28_0 <=( _mesh_3_3_io_out_b_0) ^ ((fiEnable && (221 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_92_0 <=( _mesh_3_3_io_out_c_0) ^ ((fiEnable && (222 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_3_io_in_control_0_shift_b <=( _mesh_3_3_io_out_control_0_shift) ^ ((fiEnable && (223 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_3_io_in_control_0_dataflow_b <=( _mesh_3_3_io_out_control_0_dataflow) ^ ((fiEnable && (224 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_3_io_in_control_0_propagate_b <=( _mesh_3_3_io_out_control_0_propagate) ^ ((fiEnable && (225 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_3_io_out_valid_0) begin
			b_29_0 <=( _mesh_4_3_io_out_b_0) ^ ((fiEnable && (226 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_93_0 <=( _mesh_4_3_io_out_c_0) ^ ((fiEnable && (227 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_3_io_in_control_0_shift_b <=( _mesh_4_3_io_out_control_0_shift) ^ ((fiEnable && (228 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_3_io_in_control_0_dataflow_b <=( _mesh_4_3_io_out_control_0_dataflow) ^ ((fiEnable && (229 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_3_io_in_control_0_propagate_b <=( _mesh_4_3_io_out_control_0_propagate) ^ ((fiEnable && (230 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_3_io_out_valid_0) begin
			b_30_0 <=( _mesh_5_3_io_out_b_0) ^ ((fiEnable && (231 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_94_0 <=( _mesh_5_3_io_out_c_0) ^ ((fiEnable && (232 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_3_io_in_control_0_shift_b <=( _mesh_5_3_io_out_control_0_shift) ^ ((fiEnable && (233 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_3_io_in_control_0_dataflow_b <=( _mesh_5_3_io_out_control_0_dataflow) ^ ((fiEnable && (234 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_3_io_in_control_0_propagate_b <=( _mesh_5_3_io_out_control_0_propagate) ^ ((fiEnable && (235 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_3_io_out_valid_0) begin
			b_31_0 <=( _mesh_6_3_io_out_b_0) ^ ((fiEnable && (236 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_95_0 <=( _mesh_6_3_io_out_c_0) ^ ((fiEnable && (237 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_3_io_in_control_0_shift_b <=( _mesh_6_3_io_out_control_0_shift) ^ ((fiEnable && (238 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_3_io_in_control_0_dataflow_b <=( _mesh_6_3_io_out_control_0_dataflow) ^ ((fiEnable && (239 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_3_io_in_control_0_propagate_b <=( _mesh_6_3_io_out_control_0_propagate) ^ ((fiEnable && (240 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_4_0) begin
			b_32_0 <=( io_in_b_4_0) ^ ((fiEnable && (241 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_96_0 <=( io_in_d_4_0) ^ ((fiEnable && (242 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_4_io_in_control_0_shift_b <=( io_in_control_4_0_shift) ^ ((fiEnable && (243 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_4_io_in_control_0_dataflow_b <=( io_in_control_4_0_dataflow) ^ ((fiEnable && (244 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_4_io_in_control_0_propagate_b <=( io_in_control_4_0_propagate) ^ ((fiEnable && (245 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_4_io_out_valid_0) begin
			b_33_0 <=( _mesh_0_4_io_out_b_0) ^ ((fiEnable && (246 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_97_0 <=( _mesh_0_4_io_out_c_0) ^ ((fiEnable && (247 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_4_io_in_control_0_shift_b <=( _mesh_0_4_io_out_control_0_shift) ^ ((fiEnable && (248 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_4_io_in_control_0_dataflow_b <=( _mesh_0_4_io_out_control_0_dataflow) ^ ((fiEnable && (249 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_4_io_in_control_0_propagate_b <=( _mesh_0_4_io_out_control_0_propagate) ^ ((fiEnable && (250 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_4_io_out_valid_0) begin
			b_34_0 <=( _mesh_1_4_io_out_b_0) ^ ((fiEnable && (251 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_98_0 <=( _mesh_1_4_io_out_c_0) ^ ((fiEnable && (252 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_4_io_in_control_0_shift_b <=( _mesh_1_4_io_out_control_0_shift) ^ ((fiEnable && (253 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_4_io_in_control_0_dataflow_b <=( _mesh_1_4_io_out_control_0_dataflow) ^ ((fiEnable && (254 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_4_io_in_control_0_propagate_b <=( _mesh_1_4_io_out_control_0_propagate) ^ ((fiEnable && (255 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_4_io_out_valid_0) begin
			b_35_0 <=( _mesh_2_4_io_out_b_0) ^ ((fiEnable && (256 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_99_0 <=( _mesh_2_4_io_out_c_0) ^ ((fiEnable && (257 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_4_io_in_control_0_shift_b <=( _mesh_2_4_io_out_control_0_shift) ^ ((fiEnable && (258 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_4_io_in_control_0_dataflow_b <=( _mesh_2_4_io_out_control_0_dataflow) ^ ((fiEnable && (259 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_4_io_in_control_0_propagate_b <=( _mesh_2_4_io_out_control_0_propagate) ^ ((fiEnable && (260 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_4_io_out_valid_0) begin
			b_36_0 <=( _mesh_3_4_io_out_b_0) ^ ((fiEnable && (261 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_100_0 <=( _mesh_3_4_io_out_c_0) ^ ((fiEnable && (262 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_4_io_in_control_0_shift_b <=( _mesh_3_4_io_out_control_0_shift) ^ ((fiEnable && (263 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_4_io_in_control_0_dataflow_b <=( _mesh_3_4_io_out_control_0_dataflow) ^ ((fiEnable && (264 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_4_io_in_control_0_propagate_b <=( _mesh_3_4_io_out_control_0_propagate) ^ ((fiEnable && (265 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_4_io_out_valid_0) begin
			b_37_0 <=( _mesh_4_4_io_out_b_0) ^ ((fiEnable && (266 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_101_0 <=( _mesh_4_4_io_out_c_0) ^ ((fiEnable && (267 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_4_io_in_control_0_shift_b <=( _mesh_4_4_io_out_control_0_shift) ^ ((fiEnable && (268 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_4_io_in_control_0_dataflow_b <=( _mesh_4_4_io_out_control_0_dataflow) ^ ((fiEnable && (269 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_4_io_in_control_0_propagate_b <=( _mesh_4_4_io_out_control_0_propagate) ^ ((fiEnable && (270 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_4_io_out_valid_0) begin
			b_38_0 <=( _mesh_5_4_io_out_b_0) ^ ((fiEnable && (271 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_102_0 <=( _mesh_5_4_io_out_c_0) ^ ((fiEnable && (272 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_4_io_in_control_0_shift_b <=( _mesh_5_4_io_out_control_0_shift) ^ ((fiEnable && (273 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_4_io_in_control_0_dataflow_b <=( _mesh_5_4_io_out_control_0_dataflow) ^ ((fiEnable && (274 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_4_io_in_control_0_propagate_b <=( _mesh_5_4_io_out_control_0_propagate) ^ ((fiEnable && (275 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_4_io_out_valid_0) begin
			b_39_0 <=( _mesh_6_4_io_out_b_0) ^ ((fiEnable && (276 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_103_0 <=( _mesh_6_4_io_out_c_0) ^ ((fiEnable && (277 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_4_io_in_control_0_shift_b <=( _mesh_6_4_io_out_control_0_shift) ^ ((fiEnable && (278 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_4_io_in_control_0_dataflow_b <=( _mesh_6_4_io_out_control_0_dataflow) ^ ((fiEnable && (279 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_4_io_in_control_0_propagate_b <=( _mesh_6_4_io_out_control_0_propagate) ^ ((fiEnable && (280 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_5_0) begin
			b_40_0 <=( io_in_b_5_0) ^ ((fiEnable && (281 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_104_0 <=( io_in_d_5_0) ^ ((fiEnable && (282 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_5_io_in_control_0_shift_b <=( io_in_control_5_0_shift) ^ ((fiEnable && (283 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_5_io_in_control_0_dataflow_b <=( io_in_control_5_0_dataflow) ^ ((fiEnable && (284 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_5_io_in_control_0_propagate_b <=( io_in_control_5_0_propagate) ^ ((fiEnable && (285 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_5_io_out_valid_0) begin
			b_41_0 <=( _mesh_0_5_io_out_b_0) ^ ((fiEnable && (286 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_105_0 <=( _mesh_0_5_io_out_c_0) ^ ((fiEnable && (287 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_5_io_in_control_0_shift_b <=( _mesh_0_5_io_out_control_0_shift) ^ ((fiEnable && (288 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_5_io_in_control_0_dataflow_b <=( _mesh_0_5_io_out_control_0_dataflow) ^ ((fiEnable && (289 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_5_io_in_control_0_propagate_b <=( _mesh_0_5_io_out_control_0_propagate) ^ ((fiEnable && (290 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_5_io_out_valid_0) begin
			b_42_0 <=( _mesh_1_5_io_out_b_0) ^ ((fiEnable && (291 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_106_0 <=( _mesh_1_5_io_out_c_0) ^ ((fiEnable && (292 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_5_io_in_control_0_shift_b <=( _mesh_1_5_io_out_control_0_shift) ^ ((fiEnable && (293 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_5_io_in_control_0_dataflow_b <=( _mesh_1_5_io_out_control_0_dataflow) ^ ((fiEnable && (294 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_5_io_in_control_0_propagate_b <=( _mesh_1_5_io_out_control_0_propagate) ^ ((fiEnable && (295 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_5_io_out_valid_0) begin
			b_43_0 <=( _mesh_2_5_io_out_b_0) ^ ((fiEnable && (296 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_107_0 <=( _mesh_2_5_io_out_c_0) ^ ((fiEnable && (297 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_5_io_in_control_0_shift_b <=( _mesh_2_5_io_out_control_0_shift) ^ ((fiEnable && (298 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_5_io_in_control_0_dataflow_b <=( _mesh_2_5_io_out_control_0_dataflow) ^ ((fiEnable && (299 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_5_io_in_control_0_propagate_b <=( _mesh_2_5_io_out_control_0_propagate) ^ ((fiEnable && (300 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_5_io_out_valid_0) begin
			b_44_0 <=( _mesh_3_5_io_out_b_0) ^ ((fiEnable && (301 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_108_0 <=( _mesh_3_5_io_out_c_0) ^ ((fiEnable && (302 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_5_io_in_control_0_shift_b <=( _mesh_3_5_io_out_control_0_shift) ^ ((fiEnable && (303 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_5_io_in_control_0_dataflow_b <=( _mesh_3_5_io_out_control_0_dataflow) ^ ((fiEnable && (304 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_5_io_in_control_0_propagate_b <=( _mesh_3_5_io_out_control_0_propagate) ^ ((fiEnable && (305 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_5_io_out_valid_0) begin
			b_45_0 <=( _mesh_4_5_io_out_b_0) ^ ((fiEnable && (306 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_109_0 <=( _mesh_4_5_io_out_c_0) ^ ((fiEnable && (307 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_5_io_in_control_0_shift_b <=( _mesh_4_5_io_out_control_0_shift) ^ ((fiEnable && (308 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_5_io_in_control_0_dataflow_b <=( _mesh_4_5_io_out_control_0_dataflow) ^ ((fiEnable && (309 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_5_io_in_control_0_propagate_b <=( _mesh_4_5_io_out_control_0_propagate) ^ ((fiEnable && (310 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_5_io_out_valid_0) begin
			b_46_0 <=( _mesh_5_5_io_out_b_0) ^ ((fiEnable && (311 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_110_0 <=( _mesh_5_5_io_out_c_0) ^ ((fiEnable && (312 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_5_io_in_control_0_shift_b <=( _mesh_5_5_io_out_control_0_shift) ^ ((fiEnable && (313 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_5_io_in_control_0_dataflow_b <=( _mesh_5_5_io_out_control_0_dataflow) ^ ((fiEnable && (314 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_5_io_in_control_0_propagate_b <=( _mesh_5_5_io_out_control_0_propagate) ^ ((fiEnable && (315 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_5_io_out_valid_0) begin
			b_47_0 <=( _mesh_6_5_io_out_b_0) ^ ((fiEnable && (316 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_111_0 <=( _mesh_6_5_io_out_c_0) ^ ((fiEnable && (317 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_5_io_in_control_0_shift_b <=( _mesh_6_5_io_out_control_0_shift) ^ ((fiEnable && (318 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_5_io_in_control_0_dataflow_b <=( _mesh_6_5_io_out_control_0_dataflow) ^ ((fiEnable && (319 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_5_io_in_control_0_propagate_b <=( _mesh_6_5_io_out_control_0_propagate) ^ ((fiEnable && (320 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_6_0) begin
			b_48_0 <=( io_in_b_6_0) ^ ((fiEnable && (321 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_112_0 <=( io_in_d_6_0) ^ ((fiEnable && (322 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_6_io_in_control_0_shift_b <=( io_in_control_6_0_shift) ^ ((fiEnable && (323 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_6_io_in_control_0_dataflow_b <=( io_in_control_6_0_dataflow) ^ ((fiEnable && (324 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_6_io_in_control_0_propagate_b <=( io_in_control_6_0_propagate) ^ ((fiEnable && (325 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_6_io_out_valid_0) begin
			b_49_0 <=( _mesh_0_6_io_out_b_0) ^ ((fiEnable && (326 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_113_0 <=( _mesh_0_6_io_out_c_0) ^ ((fiEnable && (327 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_6_io_in_control_0_shift_b <=( _mesh_0_6_io_out_control_0_shift) ^ ((fiEnable && (328 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_6_io_in_control_0_dataflow_b <=( _mesh_0_6_io_out_control_0_dataflow) ^ ((fiEnable && (329 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_6_io_in_control_0_propagate_b <=( _mesh_0_6_io_out_control_0_propagate) ^ ((fiEnable && (330 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_6_io_out_valid_0) begin
			b_50_0 <=( _mesh_1_6_io_out_b_0) ^ ((fiEnable && (331 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_114_0 <=( _mesh_1_6_io_out_c_0) ^ ((fiEnable && (332 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_6_io_in_control_0_shift_b <=( _mesh_1_6_io_out_control_0_shift) ^ ((fiEnable && (333 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_6_io_in_control_0_dataflow_b <=( _mesh_1_6_io_out_control_0_dataflow) ^ ((fiEnable && (334 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_6_io_in_control_0_propagate_b <=( _mesh_1_6_io_out_control_0_propagate) ^ ((fiEnable && (335 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_6_io_out_valid_0) begin
			b_51_0 <=( _mesh_2_6_io_out_b_0) ^ ((fiEnable && (336 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_115_0 <=( _mesh_2_6_io_out_c_0) ^ ((fiEnable && (337 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_6_io_in_control_0_shift_b <=( _mesh_2_6_io_out_control_0_shift) ^ ((fiEnable && (338 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_6_io_in_control_0_dataflow_b <=( _mesh_2_6_io_out_control_0_dataflow) ^ ((fiEnable && (339 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_6_io_in_control_0_propagate_b <=( _mesh_2_6_io_out_control_0_propagate) ^ ((fiEnable && (340 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_6_io_out_valid_0) begin
			b_52_0 <=( _mesh_3_6_io_out_b_0) ^ ((fiEnable && (341 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_116_0 <=( _mesh_3_6_io_out_c_0) ^ ((fiEnable && (342 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_6_io_in_control_0_shift_b <=( _mesh_3_6_io_out_control_0_shift) ^ ((fiEnable && (343 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_6_io_in_control_0_dataflow_b <=( _mesh_3_6_io_out_control_0_dataflow) ^ ((fiEnable && (344 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_6_io_in_control_0_propagate_b <=( _mesh_3_6_io_out_control_0_propagate) ^ ((fiEnable && (345 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_6_io_out_valid_0) begin
			b_53_0 <=( _mesh_4_6_io_out_b_0) ^ ((fiEnable && (346 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_117_0 <=( _mesh_4_6_io_out_c_0) ^ ((fiEnable && (347 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_6_io_in_control_0_shift_b <=( _mesh_4_6_io_out_control_0_shift) ^ ((fiEnable && (348 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_6_io_in_control_0_dataflow_b <=( _mesh_4_6_io_out_control_0_dataflow) ^ ((fiEnable && (349 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_6_io_in_control_0_propagate_b <=( _mesh_4_6_io_out_control_0_propagate) ^ ((fiEnable && (350 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_6_io_out_valid_0) begin
			b_54_0 <=( _mesh_5_6_io_out_b_0) ^ ((fiEnable && (351 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_118_0 <=( _mesh_5_6_io_out_c_0) ^ ((fiEnable && (352 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_6_io_in_control_0_shift_b <=( _mesh_5_6_io_out_control_0_shift) ^ ((fiEnable && (353 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_6_io_in_control_0_dataflow_b <=( _mesh_5_6_io_out_control_0_dataflow) ^ ((fiEnable && (354 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_6_io_in_control_0_propagate_b <=( _mesh_5_6_io_out_control_0_propagate) ^ ((fiEnable && (355 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_6_io_out_valid_0) begin
			b_55_0 <=( _mesh_6_6_io_out_b_0) ^ ((fiEnable && (356 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_119_0 <=( _mesh_6_6_io_out_c_0) ^ ((fiEnable && (357 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_6_io_in_control_0_shift_b <=( _mesh_6_6_io_out_control_0_shift) ^ ((fiEnable && (358 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_6_io_in_control_0_dataflow_b <=( _mesh_6_6_io_out_control_0_dataflow) ^ ((fiEnable && (359 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_6_io_in_control_0_propagate_b <=( _mesh_6_6_io_out_control_0_propagate) ^ ((fiEnable && (360 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (io_in_valid_7_0) begin
			b_56_0 <=( io_in_b_7_0) ^ ((fiEnable && (361 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_120_0 <=( io_in_d_7_0) ^ ((fiEnable && (362 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_0_7_io_in_control_0_shift_b <=( io_in_control_7_0_shift) ^ ((fiEnable && (363 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_0_7_io_in_control_0_dataflow_b <=( io_in_control_7_0_dataflow) ^ ((fiEnable && (364 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_0_7_io_in_control_0_propagate_b <=( io_in_control_7_0_propagate) ^ ((fiEnable && (365 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_0_7_io_out_valid_0) begin
			b_57_0 <=( _mesh_0_7_io_out_b_0) ^ ((fiEnable && (366 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_121_0 <=( _mesh_0_7_io_out_c_0) ^ ((fiEnable && (367 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_1_7_io_in_control_0_shift_b <=( _mesh_0_7_io_out_control_0_shift) ^ ((fiEnable && (368 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_1_7_io_in_control_0_dataflow_b <=( _mesh_0_7_io_out_control_0_dataflow) ^ ((fiEnable && (369 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_1_7_io_in_control_0_propagate_b <=( _mesh_0_7_io_out_control_0_propagate) ^ ((fiEnable && (370 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_1_7_io_out_valid_0) begin
			b_58_0 <=( _mesh_1_7_io_out_b_0) ^ ((fiEnable && (371 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_122_0 <=( _mesh_1_7_io_out_c_0) ^ ((fiEnable && (372 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_2_7_io_in_control_0_shift_b <=( _mesh_1_7_io_out_control_0_shift) ^ ((fiEnable && (373 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_2_7_io_in_control_0_dataflow_b <=( _mesh_1_7_io_out_control_0_dataflow) ^ ((fiEnable && (374 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_2_7_io_in_control_0_propagate_b <=( _mesh_1_7_io_out_control_0_propagate) ^ ((fiEnable && (375 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_2_7_io_out_valid_0) begin
			b_59_0 <=( _mesh_2_7_io_out_b_0) ^ ((fiEnable && (376 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_123_0 <=( _mesh_2_7_io_out_c_0) ^ ((fiEnable && (377 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_3_7_io_in_control_0_shift_b <=( _mesh_2_7_io_out_control_0_shift) ^ ((fiEnable && (378 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_3_7_io_in_control_0_dataflow_b <=( _mesh_2_7_io_out_control_0_dataflow) ^ ((fiEnable && (379 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_3_7_io_in_control_0_propagate_b <=( _mesh_2_7_io_out_control_0_propagate) ^ ((fiEnable && (380 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_3_7_io_out_valid_0) begin
			b_60_0 <=( _mesh_3_7_io_out_b_0) ^ ((fiEnable && (381 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_124_0 <=( _mesh_3_7_io_out_c_0) ^ ((fiEnable && (382 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_4_7_io_in_control_0_shift_b <=( _mesh_3_7_io_out_control_0_shift) ^ ((fiEnable && (383 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_4_7_io_in_control_0_dataflow_b <=( _mesh_3_7_io_out_control_0_dataflow) ^ ((fiEnable && (384 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_4_7_io_in_control_0_propagate_b <=( _mesh_3_7_io_out_control_0_propagate) ^ ((fiEnable && (385 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_4_7_io_out_valid_0) begin
			b_61_0 <=( _mesh_4_7_io_out_b_0) ^ ((fiEnable && (386 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_125_0 <=( _mesh_4_7_io_out_c_0) ^ ((fiEnable && (387 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_5_7_io_in_control_0_shift_b <=( _mesh_4_7_io_out_control_0_shift) ^ ((fiEnable && (388 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_5_7_io_in_control_0_dataflow_b <=( _mesh_4_7_io_out_control_0_dataflow) ^ ((fiEnable && (389 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_5_7_io_in_control_0_propagate_b <=( _mesh_4_7_io_out_control_0_propagate) ^ ((fiEnable && (390 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_5_7_io_out_valid_0) begin
			b_62_0 <=( _mesh_5_7_io_out_b_0) ^ ((fiEnable && (391 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_126_0 <=( _mesh_5_7_io_out_c_0) ^ ((fiEnable && (392 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_6_7_io_in_control_0_shift_b <=( _mesh_5_7_io_out_control_0_shift) ^ ((fiEnable && (393 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_6_7_io_in_control_0_dataflow_b <=( _mesh_5_7_io_out_control_0_dataflow) ^ ((fiEnable && (394 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_6_7_io_in_control_0_propagate_b <=( _mesh_5_7_io_out_control_0_propagate) ^ ((fiEnable && (395 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		if (_mesh_6_7_io_out_valid_0) begin
			b_63_0 <=( _mesh_6_7_io_out_b_0) ^ ((fiEnable && (396 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			b_127_0 <=( _mesh_6_7_io_out_c_0) ^ ((fiEnable && (397 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
			mesh_7_7_io_in_control_0_shift_b <=( _mesh_6_7_io_out_control_0_shift) ^ ((fiEnable && (398 == GlobalFiNumber)) ? GlobalFiSignal[4:0] : {5{1'b0}});
			mesh_7_7_io_in_control_0_dataflow_b <=( _mesh_6_7_io_out_control_0_dataflow) ^ ((fiEnable && (399 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
			mesh_7_7_io_in_control_0_propagate_b <=( _mesh_6_7_io_out_control_0_propagate) ^ ((fiEnable && (400 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		end
		r_64_0 <=( io_in_valid_0_0) ^ ((fiEnable && (401 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_65_0 <=( _mesh_0_0_io_out_valid_0) ^ ((fiEnable && (402 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_66_0 <=( _mesh_1_0_io_out_valid_0) ^ ((fiEnable && (403 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_67_0 <=( _mesh_2_0_io_out_valid_0) ^ ((fiEnable && (404 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_68_0 <=( _mesh_3_0_io_out_valid_0) ^ ((fiEnable && (405 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_69_0 <=( _mesh_4_0_io_out_valid_0) ^ ((fiEnable && (406 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_70_0 <=( _mesh_5_0_io_out_valid_0) ^ ((fiEnable && (407 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_71_0 <=( _mesh_6_0_io_out_valid_0) ^ ((fiEnable && (408 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_72_0 <=( io_in_valid_1_0) ^ ((fiEnable && (409 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_73_0 <=( _mesh_0_1_io_out_valid_0) ^ ((fiEnable && (410 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_74_0 <=( _mesh_1_1_io_out_valid_0) ^ ((fiEnable && (411 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_75_0 <=( _mesh_2_1_io_out_valid_0) ^ ((fiEnable && (412 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_76_0 <=( _mesh_3_1_io_out_valid_0) ^ ((fiEnable && (413 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_77_0 <=( _mesh_4_1_io_out_valid_0) ^ ((fiEnable && (414 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_78_0 <=( _mesh_5_1_io_out_valid_0) ^ ((fiEnable && (415 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_79_0 <=( _mesh_6_1_io_out_valid_0) ^ ((fiEnable && (416 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_80_0 <=( io_in_valid_2_0) ^ ((fiEnable && (417 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_81_0 <=( _mesh_0_2_io_out_valid_0) ^ ((fiEnable && (418 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_82_0 <=( _mesh_1_2_io_out_valid_0) ^ ((fiEnable && (419 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_83_0 <=( _mesh_2_2_io_out_valid_0) ^ ((fiEnable && (420 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_84_0 <=( _mesh_3_2_io_out_valid_0) ^ ((fiEnable && (421 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_85_0 <=( _mesh_4_2_io_out_valid_0) ^ ((fiEnable && (422 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_86_0 <=( _mesh_5_2_io_out_valid_0) ^ ((fiEnable && (423 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_87_0 <=( _mesh_6_2_io_out_valid_0) ^ ((fiEnable && (424 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_88_0 <=( io_in_valid_3_0) ^ ((fiEnable && (425 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_89_0 <=( _mesh_0_3_io_out_valid_0) ^ ((fiEnable && (426 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_90_0 <=( _mesh_1_3_io_out_valid_0) ^ ((fiEnable && (427 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_91_0 <=( _mesh_2_3_io_out_valid_0) ^ ((fiEnable && (428 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_92_0 <=( _mesh_3_3_io_out_valid_0) ^ ((fiEnable && (429 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_93_0 <=( _mesh_4_3_io_out_valid_0) ^ ((fiEnable && (430 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_94_0 <=( _mesh_5_3_io_out_valid_0) ^ ((fiEnable && (431 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_95_0 <=( _mesh_6_3_io_out_valid_0) ^ ((fiEnable && (432 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_96_0 <=( io_in_valid_4_0) ^ ((fiEnable && (433 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_97_0 <=( _mesh_0_4_io_out_valid_0) ^ ((fiEnable && (434 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_98_0 <=( _mesh_1_4_io_out_valid_0) ^ ((fiEnable && (435 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_99_0 <=( _mesh_2_4_io_out_valid_0) ^ ((fiEnable && (436 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_100_0 <=( _mesh_3_4_io_out_valid_0) ^ ((fiEnable && (437 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_101_0 <=( _mesh_4_4_io_out_valid_0) ^ ((fiEnable && (438 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_102_0 <=( _mesh_5_4_io_out_valid_0) ^ ((fiEnable && (439 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_103_0 <=( _mesh_6_4_io_out_valid_0) ^ ((fiEnable && (440 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_104_0 <=( io_in_valid_5_0) ^ ((fiEnable && (441 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_105_0 <=( _mesh_0_5_io_out_valid_0) ^ ((fiEnable && (442 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_106_0 <=( _mesh_1_5_io_out_valid_0) ^ ((fiEnable && (443 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_107_0 <=( _mesh_2_5_io_out_valid_0) ^ ((fiEnable && (444 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_108_0 <=( _mesh_3_5_io_out_valid_0) ^ ((fiEnable && (445 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_109_0 <=( _mesh_4_5_io_out_valid_0) ^ ((fiEnable && (446 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_110_0 <=( _mesh_5_5_io_out_valid_0) ^ ((fiEnable && (447 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_111_0 <=( _mesh_6_5_io_out_valid_0) ^ ((fiEnable && (448 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_112_0 <=( io_in_valid_6_0) ^ ((fiEnable && (449 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_113_0 <=( _mesh_0_6_io_out_valid_0) ^ ((fiEnable && (450 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_114_0 <=( _mesh_1_6_io_out_valid_0) ^ ((fiEnable && (451 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_115_0 <=( _mesh_2_6_io_out_valid_0) ^ ((fiEnable && (452 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_116_0 <=( _mesh_3_6_io_out_valid_0) ^ ((fiEnable && (453 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_117_0 <=( _mesh_4_6_io_out_valid_0) ^ ((fiEnable && (454 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_118_0 <=( _mesh_5_6_io_out_valid_0) ^ ((fiEnable && (455 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_119_0 <=( _mesh_6_6_io_out_valid_0) ^ ((fiEnable && (456 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_120_0 <=( io_in_valid_7_0) ^ ((fiEnable && (457 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_121_0 <=( _mesh_0_7_io_out_valid_0) ^ ((fiEnable && (458 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_122_0 <=( _mesh_1_7_io_out_valid_0) ^ ((fiEnable && (459 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_123_0 <=( _mesh_2_7_io_out_valid_0) ^ ((fiEnable && (460 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_124_0 <=( _mesh_3_7_io_out_valid_0) ^ ((fiEnable && (461 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_125_0 <=( _mesh_4_7_io_out_valid_0) ^ ((fiEnable && (462 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_126_0 <=( _mesh_5_7_io_out_valid_0) ^ ((fiEnable && (463 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_127_0 <=( _mesh_6_7_io_out_valid_0) ^ ((fiEnable && (464 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_128_0 <=( io_in_id_0_0) ^ ((fiEnable && (465 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_129_0 <=( _mesh_0_0_io_out_id_0) ^ ((fiEnable && (466 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_130_0 <=( _mesh_1_0_io_out_id_0) ^ ((fiEnable && (467 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_131_0 <=( _mesh_2_0_io_out_id_0) ^ ((fiEnable && (468 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_132_0 <=( _mesh_3_0_io_out_id_0) ^ ((fiEnable && (469 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_133_0 <=( _mesh_4_0_io_out_id_0) ^ ((fiEnable && (470 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_134_0 <=( _mesh_5_0_io_out_id_0) ^ ((fiEnable && (471 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_135_0 <=( _mesh_6_0_io_out_id_0) ^ ((fiEnable && (472 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_136_0 <=( io_in_id_1_0) ^ ((fiEnable && (473 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_137_0 <=( _mesh_0_1_io_out_id_0) ^ ((fiEnable && (474 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_138_0 <=( _mesh_1_1_io_out_id_0) ^ ((fiEnable && (475 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_139_0 <=( _mesh_2_1_io_out_id_0) ^ ((fiEnable && (476 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_140_0 <=( _mesh_3_1_io_out_id_0) ^ ((fiEnable && (477 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_141_0 <=( _mesh_4_1_io_out_id_0) ^ ((fiEnable && (478 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_142_0 <=( _mesh_5_1_io_out_id_0) ^ ((fiEnable && (479 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_143_0 <=( _mesh_6_1_io_out_id_0) ^ ((fiEnable && (480 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_144_0 <=( io_in_id_2_0) ^ ((fiEnable && (481 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_145_0 <=( _mesh_0_2_io_out_id_0) ^ ((fiEnable && (482 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_146_0 <=( _mesh_1_2_io_out_id_0) ^ ((fiEnable && (483 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_147_0 <=( _mesh_2_2_io_out_id_0) ^ ((fiEnable && (484 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_148_0 <=( _mesh_3_2_io_out_id_0) ^ ((fiEnable && (485 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_149_0 <=( _mesh_4_2_io_out_id_0) ^ ((fiEnable && (486 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_150_0 <=( _mesh_5_2_io_out_id_0) ^ ((fiEnable && (487 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_151_0 <=( _mesh_6_2_io_out_id_0) ^ ((fiEnable && (488 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_152_0 <=( io_in_id_3_0) ^ ((fiEnable && (489 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_153_0 <=( _mesh_0_3_io_out_id_0) ^ ((fiEnable && (490 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_154_0 <=( _mesh_1_3_io_out_id_0) ^ ((fiEnable && (491 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_155_0 <=( _mesh_2_3_io_out_id_0) ^ ((fiEnable && (492 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_156_0 <=( _mesh_3_3_io_out_id_0) ^ ((fiEnable && (493 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_157_0 <=( _mesh_4_3_io_out_id_0) ^ ((fiEnable && (494 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_158_0 <=( _mesh_5_3_io_out_id_0) ^ ((fiEnable && (495 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_159_0 <=( _mesh_6_3_io_out_id_0) ^ ((fiEnable && (496 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_160_0 <=( io_in_id_4_0) ^ ((fiEnable && (497 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_161_0 <=( _mesh_0_4_io_out_id_0) ^ ((fiEnable && (498 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_162_0 <=( _mesh_1_4_io_out_id_0) ^ ((fiEnable && (499 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_163_0 <=( _mesh_2_4_io_out_id_0) ^ ((fiEnable && (500 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_164_0 <=( _mesh_3_4_io_out_id_0) ^ ((fiEnable && (501 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_165_0 <=( _mesh_4_4_io_out_id_0) ^ ((fiEnable && (502 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_166_0 <=( _mesh_5_4_io_out_id_0) ^ ((fiEnable && (503 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_167_0 <=( _mesh_6_4_io_out_id_0) ^ ((fiEnable && (504 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_168_0 <=( io_in_id_5_0) ^ ((fiEnable && (505 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_169_0 <=( _mesh_0_5_io_out_id_0) ^ ((fiEnable && (506 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_170_0 <=( _mesh_1_5_io_out_id_0) ^ ((fiEnable && (507 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_171_0 <=( _mesh_2_5_io_out_id_0) ^ ((fiEnable && (508 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_172_0 <=( _mesh_3_5_io_out_id_0) ^ ((fiEnable && (509 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_173_0 <=( _mesh_4_5_io_out_id_0) ^ ((fiEnable && (510 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_174_0 <=( _mesh_5_5_io_out_id_0) ^ ((fiEnable && (511 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_175_0 <=( _mesh_6_5_io_out_id_0) ^ ((fiEnable && (512 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_176_0 <=( io_in_id_6_0) ^ ((fiEnable && (513 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_177_0 <=( _mesh_0_6_io_out_id_0) ^ ((fiEnable && (514 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_178_0 <=( _mesh_1_6_io_out_id_0) ^ ((fiEnable && (515 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_179_0 <=( _mesh_2_6_io_out_id_0) ^ ((fiEnable && (516 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_180_0 <=( _mesh_3_6_io_out_id_0) ^ ((fiEnable && (517 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_181_0 <=( _mesh_4_6_io_out_id_0) ^ ((fiEnable && (518 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_182_0 <=( _mesh_5_6_io_out_id_0) ^ ((fiEnable && (519 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_183_0 <=( _mesh_6_6_io_out_id_0) ^ ((fiEnable && (520 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_184_0 <=( io_in_id_7_0) ^ ((fiEnable && (521 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_185_0 <=( _mesh_0_7_io_out_id_0) ^ ((fiEnable && (522 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_186_0 <=( _mesh_1_7_io_out_id_0) ^ ((fiEnable && (523 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_187_0 <=( _mesh_2_7_io_out_id_0) ^ ((fiEnable && (524 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_188_0 <=( _mesh_3_7_io_out_id_0) ^ ((fiEnable && (525 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_189_0 <=( _mesh_4_7_io_out_id_0) ^ ((fiEnable && (526 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_190_0 <=( _mesh_5_7_io_out_id_0) ^ ((fiEnable && (527 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_191_0 <=( _mesh_6_7_io_out_id_0) ^ ((fiEnable && (528 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_192_0 <=( io_in_last_0_0) ^ ((fiEnable && (529 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_193_0 <=( _mesh_0_0_io_out_last_0) ^ ((fiEnable && (530 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_194_0 <=( _mesh_1_0_io_out_last_0) ^ ((fiEnable && (531 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_195_0 <=( _mesh_2_0_io_out_last_0) ^ ((fiEnable && (532 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_196_0 <=( _mesh_3_0_io_out_last_0) ^ ((fiEnable && (533 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_197_0 <=( _mesh_4_0_io_out_last_0) ^ ((fiEnable && (534 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_198_0 <=( _mesh_5_0_io_out_last_0) ^ ((fiEnable && (535 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_199_0 <=( _mesh_6_0_io_out_last_0) ^ ((fiEnable && (536 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_200_0 <=( io_in_last_1_0) ^ ((fiEnable && (537 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_201_0 <=( _mesh_0_1_io_out_last_0) ^ ((fiEnable && (538 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_202_0 <=( _mesh_1_1_io_out_last_0) ^ ((fiEnable && (539 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_203_0 <=( _mesh_2_1_io_out_last_0) ^ ((fiEnable && (540 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_204_0 <=( _mesh_3_1_io_out_last_0) ^ ((fiEnable && (541 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_205_0 <=( _mesh_4_1_io_out_last_0) ^ ((fiEnable && (542 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_206_0 <=( _mesh_5_1_io_out_last_0) ^ ((fiEnable && (543 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_207_0 <=( _mesh_6_1_io_out_last_0) ^ ((fiEnable && (544 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_208_0 <=( io_in_last_2_0) ^ ((fiEnable && (545 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_209_0 <=( _mesh_0_2_io_out_last_0) ^ ((fiEnable && (546 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_210_0 <=( _mesh_1_2_io_out_last_0) ^ ((fiEnable && (547 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_211_0 <=( _mesh_2_2_io_out_last_0) ^ ((fiEnable && (548 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_212_0 <=( _mesh_3_2_io_out_last_0) ^ ((fiEnable && (549 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_213_0 <=( _mesh_4_2_io_out_last_0) ^ ((fiEnable && (550 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_214_0 <=( _mesh_5_2_io_out_last_0) ^ ((fiEnable && (551 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_215_0 <=( _mesh_6_2_io_out_last_0) ^ ((fiEnable && (552 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_216_0 <=( io_in_last_3_0) ^ ((fiEnable && (553 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_217_0 <=( _mesh_0_3_io_out_last_0) ^ ((fiEnable && (554 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_218_0 <=( _mesh_1_3_io_out_last_0) ^ ((fiEnable && (555 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_219_0 <=( _mesh_2_3_io_out_last_0) ^ ((fiEnable && (556 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_220_0 <=( _mesh_3_3_io_out_last_0) ^ ((fiEnable && (557 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_221_0 <=( _mesh_4_3_io_out_last_0) ^ ((fiEnable && (558 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_222_0 <=( _mesh_5_3_io_out_last_0) ^ ((fiEnable && (559 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_223_0 <=( _mesh_6_3_io_out_last_0) ^ ((fiEnable && (560 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_224_0 <=( io_in_last_4_0) ^ ((fiEnable && (561 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_225_0 <=( _mesh_0_4_io_out_last_0) ^ ((fiEnable && (562 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_226_0 <=( _mesh_1_4_io_out_last_0) ^ ((fiEnable && (563 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_227_0 <=( _mesh_2_4_io_out_last_0) ^ ((fiEnable && (564 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_228_0 <=( _mesh_3_4_io_out_last_0) ^ ((fiEnable && (565 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_229_0 <=( _mesh_4_4_io_out_last_0) ^ ((fiEnable && (566 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_230_0 <=( _mesh_5_4_io_out_last_0) ^ ((fiEnable && (567 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_231_0 <=( _mesh_6_4_io_out_last_0) ^ ((fiEnable && (568 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_232_0 <=( io_in_last_5_0) ^ ((fiEnable && (569 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_233_0 <=( _mesh_0_5_io_out_last_0) ^ ((fiEnable && (570 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_234_0 <=( _mesh_1_5_io_out_last_0) ^ ((fiEnable && (571 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_235_0 <=( _mesh_2_5_io_out_last_0) ^ ((fiEnable && (572 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_236_0 <=( _mesh_3_5_io_out_last_0) ^ ((fiEnable && (573 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_237_0 <=( _mesh_4_5_io_out_last_0) ^ ((fiEnable && (574 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_238_0 <=( _mesh_5_5_io_out_last_0) ^ ((fiEnable && (575 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_239_0 <=( _mesh_6_5_io_out_last_0) ^ ((fiEnable && (576 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_240_0 <=( io_in_last_6_0) ^ ((fiEnable && (577 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_241_0 <=( _mesh_0_6_io_out_last_0) ^ ((fiEnable && (578 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_242_0 <=( _mesh_1_6_io_out_last_0) ^ ((fiEnable && (579 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_243_0 <=( _mesh_2_6_io_out_last_0) ^ ((fiEnable && (580 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_244_0 <=( _mesh_3_6_io_out_last_0) ^ ((fiEnable && (581 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_245_0 <=( _mesh_4_6_io_out_last_0) ^ ((fiEnable && (582 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_246_0 <=( _mesh_5_6_io_out_last_0) ^ ((fiEnable && (583 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_247_0 <=( _mesh_6_6_io_out_last_0) ^ ((fiEnable && (584 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_248_0 <=( io_in_last_7_0) ^ ((fiEnable && (585 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_249_0 <=( _mesh_0_7_io_out_last_0) ^ ((fiEnable && (586 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_250_0 <=( _mesh_1_7_io_out_last_0) ^ ((fiEnable && (587 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_251_0 <=( _mesh_2_7_io_out_last_0) ^ ((fiEnable && (588 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_252_0 <=( _mesh_3_7_io_out_last_0) ^ ((fiEnable && (589 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_253_0 <=( _mesh_4_7_io_out_last_0) ^ ((fiEnable && (590 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_254_0 <=( _mesh_5_7_io_out_last_0) ^ ((fiEnable && (591 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_255_0 <=( _mesh_6_7_io_out_last_0) ^ ((fiEnable && (592 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_256_0 <=( _mesh_7_0_io_out_b_0) ^ ((fiEnable && (593 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_257_0 <=( _mesh_7_0_io_out_c_0) ^ ((fiEnable && (594 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_258_0 <=( _mesh_7_0_io_out_valid_0) ^ ((fiEnable && (595 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_259_0_dataflow <=( _mesh_7_0_io_out_control_0_dataflow) ^ ((fiEnable && (596 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_260_0 <=( _mesh_7_0_io_out_id_0) ^ ((fiEnable && (597 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
		r_261_0 <=( _mesh_7_0_io_out_last_0) ^ ((fiEnable && (598 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
		r_262_0 <=( _mesh_7_1_io_out_b_0) ^ ((fiEnable && (599 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_263_0 <=( _mesh_7_1_io_out_c_0) ^ ((fiEnable && (600 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_268_0 <=( _mesh_7_2_io_out_b_0) ^ ((fiEnable && (601 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_269_0 <=( _mesh_7_2_io_out_c_0) ^ ((fiEnable && (602 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_274_0 <=( _mesh_7_3_io_out_b_0) ^ ((fiEnable && (603 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_275_0 <=( _mesh_7_3_io_out_c_0) ^ ((fiEnable && (604 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_280_0 <=( _mesh_7_4_io_out_b_0) ^ ((fiEnable && (605 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_281_0 <=( _mesh_7_4_io_out_c_0) ^ ((fiEnable && (606 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_286_0 <=( _mesh_7_5_io_out_b_0) ^ ((fiEnable && (607 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_287_0 <=( _mesh_7_5_io_out_c_0) ^ ((fiEnable && (608 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_292_0 <=( _mesh_7_6_io_out_b_0) ^ ((fiEnable && (609 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_293_0 <=( _mesh_7_6_io_out_c_0) ^ ((fiEnable && (610 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_298_0 <=( _mesh_7_7_io_out_b_0) ^ ((fiEnable && (611 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
		r_299_0 <=( _mesh_7_7_io_out_c_0) ^ ((fiEnable && (612 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	end
	logic [31:0] _RANDOM_0;
	logic [31:0] _RANDOM_1;
	logic [31:0] _RANDOM_2;
	logic [31:0] _RANDOM_3;
	logic [31:0] _RANDOM_4;
	logic [31:0] _RANDOM_5;
	logic [31:0] _RANDOM_6;
	logic [31:0] _RANDOM_7;
	logic [31:0] _RANDOM_8;
	logic [31:0] _RANDOM_9;
	logic [31:0] _RANDOM_10;
	logic [31:0] _RANDOM_11;
	logic [31:0] _RANDOM_12;
	logic [31:0] _RANDOM_13;
	logic [31:0] _RANDOM_14;
	logic [31:0] _RANDOM_15;
	logic [31:0] _RANDOM_16;
	logic [31:0] _RANDOM_17;
	logic [31:0] _RANDOM_18;
	logic [31:0] _RANDOM_19;
	logic [31:0] _RANDOM_20;
	logic [31:0] _RANDOM_21;
	logic [31:0] _RANDOM_22;
	logic [31:0] _RANDOM_23;
	logic [31:0] _RANDOM_24;
	logic [31:0] _RANDOM_25;
	logic [31:0] _RANDOM_26;
	logic [31:0] _RANDOM_27;
	logic [31:0] _RANDOM_28;
	logic [31:0] _RANDOM_29;
	logic [31:0] _RANDOM_30;
	logic [31:0] _RANDOM_31;
	logic [31:0] _RANDOM_32;
	logic [31:0] _RANDOM_33;
	logic [31:0] _RANDOM_34;
	logic [31:0] _RANDOM_35;
	logic [31:0] _RANDOM_36;
	logic [31:0] _RANDOM_37;
	logic [31:0] _RANDOM_38;
	logic [31:0] _RANDOM_39;
	logic [31:0] _RANDOM_40;
	logic [31:0] _RANDOM_41;
	logic [31:0] _RANDOM_42;
	logic [31:0] _RANDOM_43;
	logic [31:0] _RANDOM_44;
	logic [31:0] _RANDOM_45;
	logic [31:0] _RANDOM_46;
	logic [31:0] _RANDOM_47;
	logic [31:0] _RANDOM_48;
	logic [31:0] _RANDOM_49;
	logic [31:0] _RANDOM_50;
	logic [31:0] _RANDOM_51;
	logic [31:0] _RANDOM_52;
	logic [31:0] _RANDOM_53;
	logic [31:0] _RANDOM_54;
	logic [31:0] _RANDOM_55;
	logic [31:0] _RANDOM_56;
	logic [31:0] _RANDOM_57;
	logic [31:0] _RANDOM_58;
	logic [31:0] _RANDOM_59;
	logic [31:0] _RANDOM_60;
	logic [31:0] _RANDOM_61;
	logic [31:0] _RANDOM_62;
	logic [31:0] _RANDOM_63;
	logic [31:0] _RANDOM_64;
	logic [31:0] _RANDOM_65;
	logic [31:0] _RANDOM_66;
	logic [31:0] _RANDOM_67;
	logic [31:0] _RANDOM_68;
	logic [31:0] _RANDOM_69;
	logic [31:0] _RANDOM_70;
	logic [31:0] _RANDOM_71;
	logic [31:0] _RANDOM_72;
	logic [31:0] _RANDOM_73;
	logic [31:0] _RANDOM_74;
	logic [31:0] _RANDOM_75;
	logic [31:0] _RANDOM_76;
	logic [31:0] _RANDOM_77;
	logic [31:0] _RANDOM_78;
	logic [31:0] _RANDOM_79;
	logic [31:0] _RANDOM_80;
	logic [31:0] _RANDOM_81;
	logic [31:0] _RANDOM_82;
	logic [31:0] _RANDOM_83;
	logic [31:0] _RANDOM_84;
	logic [31:0] _RANDOM_85;
	logic [31:0] _RANDOM_86;
	logic [31:0] _RANDOM_87;
	logic [31:0] _RANDOM_88;
	logic [31:0] _RANDOM_89;
	logic [31:0] _RANDOM_90;
	logic [31:0] _RANDOM_91;
	logic [31:0] _RANDOM_92;
	logic [31:0] _RANDOM_93;
	logic [31:0] _RANDOM_94;
	logic [31:0] _RANDOM_95;
	logic [31:0] _RANDOM_96;
	logic [31:0] _RANDOM_97;
	logic [31:0] _RANDOM_98;
	logic [31:0] _RANDOM_99;
	logic [31:0] _RANDOM_100;
	logic [31:0] _RANDOM_101;
	logic [31:0] _RANDOM_102;
	logic [31:0] _RANDOM_103;
	logic [31:0] _RANDOM_104;
	logic [31:0] _RANDOM_105;
	logic [31:0] _RANDOM_106;
	logic [31:0] _RANDOM_107;
	logic [31:0] _RANDOM_108;
	logic [31:0] _RANDOM_109;
	logic [31:0] _RANDOM_110;
	logic [31:0] _RANDOM_111;
	logic [31:0] _RANDOM_112;
	logic [31:0] _RANDOM_113;
	logic [31:0] _RANDOM_114;
	logic [31:0] _RANDOM_115;
	logic [31:0] _RANDOM_116;
	logic [31:0] _RANDOM_117;
	logic [31:0] _RANDOM_118;
	logic [31:0] _RANDOM_119;
	logic [31:0] _RANDOM_120;
	logic [31:0] _RANDOM_121;
	logic [31:0] _RANDOM_122;
	logic [31:0] _RANDOM_123;
	logic [31:0] _RANDOM_124;
	logic [31:0] _RANDOM_125;
	logic [31:0] _RANDOM_126;
	logic [31:0] _RANDOM_127;
	logic [31:0] _RANDOM_128;
	logic [31:0] _RANDOM_129;
	logic [31:0] _RANDOM_130;
	logic [31:0] _RANDOM_131;
	logic [31:0] _RANDOM_132;
	logic [31:0] _RANDOM_133;
	logic [31:0] _RANDOM_134;
	logic [31:0] _RANDOM_135;
	logic [31:0] _RANDOM_136;
	logic [31:0] _RANDOM_137;
	logic [31:0] _RANDOM_138;
	logic [31:0] _RANDOM_139;
	logic [31:0] _RANDOM_140;
	logic [31:0] _RANDOM_141;
	logic [31:0] _RANDOM_142;
	logic [31:0] _RANDOM_143;
	logic [31:0] _RANDOM_144;
	logic [31:0] _RANDOM_145;
	logic [31:0] _RANDOM_146;
	logic [31:0] _RANDOM_147;
	logic [31:0] _RANDOM_148;
	logic [31:0] _RANDOM_149;
	logic [31:0] _RANDOM_150;
	logic [31:0] _RANDOM_151;
	logic [31:0] _RANDOM_152;
	logic [31:0] _RANDOM_153;
	logic [31:0] _RANDOM_154;
	logic [31:0] _RANDOM_155;
	logic [31:0] _RANDOM_156;
	logic [31:0] _RANDOM_157;
	logic [31:0] _RANDOM_158;
	logic [31:0] _RANDOM_159;
	logic [31:0] _RANDOM_160;
	logic [31:0] _RANDOM_161;
	logic [31:0] _RANDOM_162;
	logic [31:0] _RANDOM_163;
	logic [31:0] _RANDOM_164;
	logic [31:0] _RANDOM_165;
	logic [31:0] _RANDOM_166;
	logic [31:0] _RANDOM_167;
	logic [31:0] _RANDOM_168;
	logic [31:0] _RANDOM_169;
	logic [31:0] _RANDOM_170;
	logic [31:0] _RANDOM_171;
	logic [31:0] _RANDOM_172;
	logic [31:0] _RANDOM_173;
	logic [31:0] _RANDOM_174;
	logic [31:0] _RANDOM_175;
	logic [31:0] _RANDOM_176;
	logic [31:0] _RANDOM_177;
	logic [31:0] _RANDOM_178;
	logic [31:0] _RANDOM_179;
	logic [31:0] _RANDOM_180;
	logic [31:0] _RANDOM_181;
	logic [31:0] _RANDOM_182;
	logic [31:0] _RANDOM_183;
	logic [31:0] _RANDOM_184;
	logic [31:0] _RANDOM_185;
	logic [31:0] _RANDOM_186;
	logic [31:0] _RANDOM_187;
	logic [31:0] _RANDOM_188;
	logic [31:0] _RANDOM_189;
	logic [31:0] _RANDOM_190;
	logic [31:0] _RANDOM_191;
	logic [31:0] _RANDOM_192;
	logic [31:0] _RANDOM_193;
	logic [31:0] _RANDOM_194;
	logic [31:0] _RANDOM_195;
	logic [31:0] _RANDOM_196;
	logic [31:0] _RANDOM_197;
	logic [31:0] _RANDOM_198;
	logic [31:0] _RANDOM_199;
	logic [31:0] _RANDOM_200;
	logic [31:0] _RANDOM_201;
	logic [31:0] _RANDOM_202;
	logic [31:0] _RANDOM_203;
	logic [31:0] _RANDOM_204;
	logic [31:0] _RANDOM_205;
	logic [31:0] _RANDOM_206;
	logic [31:0] _RANDOM_207;
	logic [31:0] _RANDOM_208;
	logic [31:0] _RANDOM_209;
	logic [31:0] _RANDOM_210;
	logic [31:0] _RANDOM_211;
	logic [31:0] _RANDOM_212;
	logic [31:0] _RANDOM_213;
	logic [31:0] _RANDOM_214;
	logic [31:0] _RANDOM_215;
	logic [31:0] _RANDOM_216;
	logic [31:0] _RANDOM_217;
	logic [31:0] _RANDOM_218;
	logic [31:0] _RANDOM_219;
	logic [31:0] _RANDOM_220;
	logic [31:0] _RANDOM_221;
	logic [31:0] _RANDOM_222;
	logic [31:0] _RANDOM_223;
	logic [31:0] _RANDOM_224;
	logic [31:0] _RANDOM_225;
	logic [31:0] _RANDOM_226;
	logic [31:0] _RANDOM_227;
	logic [31:0] _RANDOM_228;
	logic [31:0] _RANDOM_229;
	logic [31:0] _RANDOM_230;
	logic [31:0] _RANDOM_231;
	logic [31:0] _RANDOM_232;
	logic [31:0] _RANDOM_233;
	logic [31:0] _RANDOM_234;
	logic [31:0] _RANDOM_235;
	logic [31:0] _RANDOM_236;
	logic [31:0] _RANDOM_237;
	logic [31:0] _RANDOM_238;
	logic [31:0] _RANDOM_239;
	logic [31:0] _RANDOM_240;
	logic [31:0] _RANDOM_241;
	logic [31:0] _RANDOM_242;
	logic [31:0] _RANDOM_243;
	logic [31:0] _RANDOM_244;
	Tile mesh_0_0(
		.clock(clock),
		.io_in_a_0(r_0),
		.io_in_b_0(b_0),
		.io_in_d_0(b_64_0),
		.io_in_control_0_dataflow(mesh_0_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_0_io_in_control_0_shift_b),
		.io_in_id_0(r_128_0),
		.io_in_last_0(r_192_0),
		.io_in_valid_0(r_64_0),
		.io_out_a_0(_mesh_0_0_io_out_a_0),
		.io_out_c_0(_mesh_0_0_io_out_c_0),
		.io_out_b_0(_mesh_0_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_0_io_out_id_0),
		.io_out_last_0(_mesh_0_0_io_out_last_0),
		.io_out_valid_0(_mesh_0_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((635 == GlobalFiModInstNr[0]) || (635 == GlobalFiModInstNr[1]) || (635 == GlobalFiModInstNr[2]) || (635 == GlobalFiModInstNr[3]))));
	Tile mesh_0_1(
		.clock(clock),
		.io_in_a_0(r_1_0),
		.io_in_b_0(b_8_0),
		.io_in_d_0(b_72_0),
		.io_in_control_0_dataflow(mesh_0_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_1_io_in_control_0_shift_b),
		.io_in_id_0(r_136_0),
		.io_in_last_0(r_200_0),
		.io_in_valid_0(r_72_0),
		.io_out_a_0(_mesh_0_1_io_out_a_0),
		.io_out_c_0(_mesh_0_1_io_out_c_0),
		.io_out_b_0(_mesh_0_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_1_io_out_id_0),
		.io_out_last_0(_mesh_0_1_io_out_last_0),
		.io_out_valid_0(_mesh_0_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((636 == GlobalFiModInstNr[0]) || (636 == GlobalFiModInstNr[1]) || (636 == GlobalFiModInstNr[2]) || (636 == GlobalFiModInstNr[3]))));
	Tile mesh_0_2(
		.clock(clock),
		.io_in_a_0(r_2_0),
		.io_in_b_0(b_16_0),
		.io_in_d_0(b_80_0),
		.io_in_control_0_dataflow(mesh_0_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_2_io_in_control_0_shift_b),
		.io_in_id_0(r_144_0),
		.io_in_last_0(r_208_0),
		.io_in_valid_0(r_80_0),
		.io_out_a_0(_mesh_0_2_io_out_a_0),
		.io_out_c_0(_mesh_0_2_io_out_c_0),
		.io_out_b_0(_mesh_0_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_2_io_out_id_0),
		.io_out_last_0(_mesh_0_2_io_out_last_0),
		.io_out_valid_0(_mesh_0_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((637 == GlobalFiModInstNr[0]) || (637 == GlobalFiModInstNr[1]) || (637 == GlobalFiModInstNr[2]) || (637 == GlobalFiModInstNr[3]))));
	Tile mesh_0_3(
		.clock(clock),
		.io_in_a_0(r_3_0),
		.io_in_b_0(b_24_0),
		.io_in_d_0(b_88_0),
		.io_in_control_0_dataflow(mesh_0_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_3_io_in_control_0_shift_b),
		.io_in_id_0(r_152_0),
		.io_in_last_0(r_216_0),
		.io_in_valid_0(r_88_0),
		.io_out_a_0(_mesh_0_3_io_out_a_0),
		.io_out_c_0(_mesh_0_3_io_out_c_0),
		.io_out_b_0(_mesh_0_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_3_io_out_id_0),
		.io_out_last_0(_mesh_0_3_io_out_last_0),
		.io_out_valid_0(_mesh_0_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((638 == GlobalFiModInstNr[0]) || (638 == GlobalFiModInstNr[1]) || (638 == GlobalFiModInstNr[2]) || (638 == GlobalFiModInstNr[3]))));
	Tile mesh_0_4(
		.clock(clock),
		.io_in_a_0(r_4_0),
		.io_in_b_0(b_32_0),
		.io_in_d_0(b_96_0),
		.io_in_control_0_dataflow(mesh_0_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_4_io_in_control_0_shift_b),
		.io_in_id_0(r_160_0),
		.io_in_last_0(r_224_0),
		.io_in_valid_0(r_96_0),
		.io_out_a_0(_mesh_0_4_io_out_a_0),
		.io_out_c_0(_mesh_0_4_io_out_c_0),
		.io_out_b_0(_mesh_0_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_4_io_out_id_0),
		.io_out_last_0(_mesh_0_4_io_out_last_0),
		.io_out_valid_0(_mesh_0_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((639 == GlobalFiModInstNr[0]) || (639 == GlobalFiModInstNr[1]) || (639 == GlobalFiModInstNr[2]) || (639 == GlobalFiModInstNr[3]))));
	Tile mesh_0_5(
		.clock(clock),
		.io_in_a_0(r_5_0),
		.io_in_b_0(b_40_0),
		.io_in_d_0(b_104_0),
		.io_in_control_0_dataflow(mesh_0_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_5_io_in_control_0_shift_b),
		.io_in_id_0(r_168_0),
		.io_in_last_0(r_232_0),
		.io_in_valid_0(r_104_0),
		.io_out_a_0(_mesh_0_5_io_out_a_0),
		.io_out_c_0(_mesh_0_5_io_out_c_0),
		.io_out_b_0(_mesh_0_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_5_io_out_id_0),
		.io_out_last_0(_mesh_0_5_io_out_last_0),
		.io_out_valid_0(_mesh_0_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((640 == GlobalFiModInstNr[0]) || (640 == GlobalFiModInstNr[1]) || (640 == GlobalFiModInstNr[2]) || (640 == GlobalFiModInstNr[3]))));
	Tile mesh_0_6(
		.clock(clock),
		.io_in_a_0(r_6_0),
		.io_in_b_0(b_48_0),
		.io_in_d_0(b_112_0),
		.io_in_control_0_dataflow(mesh_0_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_6_io_in_control_0_shift_b),
		.io_in_id_0(r_176_0),
		.io_in_last_0(r_240_0),
		.io_in_valid_0(r_112_0),
		.io_out_a_0(_mesh_0_6_io_out_a_0),
		.io_out_c_0(_mesh_0_6_io_out_c_0),
		.io_out_b_0(_mesh_0_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_6_io_out_id_0),
		.io_out_last_0(_mesh_0_6_io_out_last_0),
		.io_out_valid_0(_mesh_0_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((641 == GlobalFiModInstNr[0]) || (641 == GlobalFiModInstNr[1]) || (641 == GlobalFiModInstNr[2]) || (641 == GlobalFiModInstNr[3]))));
	Tile mesh_0_7(
		.clock(clock),
		.io_in_a_0(r_7_0),
		.io_in_b_0(b_56_0),
		.io_in_d_0(b_120_0),
		.io_in_control_0_dataflow(mesh_0_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_0_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_0_7_io_in_control_0_shift_b),
		.io_in_id_0(r_184_0),
		.io_in_last_0(r_248_0),
		.io_in_valid_0(r_120_0),
		.io_out_a_0(_mesh_0_7_io_out_a_0),
		.io_out_c_0(_mesh_0_7_io_out_c_0),
		.io_out_b_0(_mesh_0_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_0_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_0_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_0_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_0_7_io_out_id_0),
		.io_out_last_0(_mesh_0_7_io_out_last_0),
		.io_out_valid_0(_mesh_0_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((642 == GlobalFiModInstNr[0]) || (642 == GlobalFiModInstNr[1]) || (642 == GlobalFiModInstNr[2]) || (642 == GlobalFiModInstNr[3]))));
	Tile mesh_1_0(
		.clock(clock),
		.io_in_a_0(r_8_0),
		.io_in_b_0(b_1_0),
		.io_in_d_0(b_65_0),
		.io_in_control_0_dataflow(mesh_1_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_0_io_in_control_0_shift_b),
		.io_in_id_0(r_129_0),
		.io_in_last_0(r_193_0),
		.io_in_valid_0(r_65_0),
		.io_out_a_0(_mesh_1_0_io_out_a_0),
		.io_out_c_0(_mesh_1_0_io_out_c_0),
		.io_out_b_0(_mesh_1_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_0_io_out_id_0),
		.io_out_last_0(_mesh_1_0_io_out_last_0),
		.io_out_valid_0(_mesh_1_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((643 == GlobalFiModInstNr[0]) || (643 == GlobalFiModInstNr[1]) || (643 == GlobalFiModInstNr[2]) || (643 == GlobalFiModInstNr[3]))));
	Tile mesh_1_1(
		.clock(clock),
		.io_in_a_0(r_9_0),
		.io_in_b_0(b_9_0),
		.io_in_d_0(b_73_0),
		.io_in_control_0_dataflow(mesh_1_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_1_io_in_control_0_shift_b),
		.io_in_id_0(r_137_0),
		.io_in_last_0(r_201_0),
		.io_in_valid_0(r_73_0),
		.io_out_a_0(_mesh_1_1_io_out_a_0),
		.io_out_c_0(_mesh_1_1_io_out_c_0),
		.io_out_b_0(_mesh_1_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_1_io_out_id_0),
		.io_out_last_0(_mesh_1_1_io_out_last_0),
		.io_out_valid_0(_mesh_1_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((644 == GlobalFiModInstNr[0]) || (644 == GlobalFiModInstNr[1]) || (644 == GlobalFiModInstNr[2]) || (644 == GlobalFiModInstNr[3]))));
	Tile mesh_1_2(
		.clock(clock),
		.io_in_a_0(r_10_0),
		.io_in_b_0(b_17_0),
		.io_in_d_0(b_81_0),
		.io_in_control_0_dataflow(mesh_1_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_2_io_in_control_0_shift_b),
		.io_in_id_0(r_145_0),
		.io_in_last_0(r_209_0),
		.io_in_valid_0(r_81_0),
		.io_out_a_0(_mesh_1_2_io_out_a_0),
		.io_out_c_0(_mesh_1_2_io_out_c_0),
		.io_out_b_0(_mesh_1_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_2_io_out_id_0),
		.io_out_last_0(_mesh_1_2_io_out_last_0),
		.io_out_valid_0(_mesh_1_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((645 == GlobalFiModInstNr[0]) || (645 == GlobalFiModInstNr[1]) || (645 == GlobalFiModInstNr[2]) || (645 == GlobalFiModInstNr[3]))));
	Tile mesh_1_3(
		.clock(clock),
		.io_in_a_0(r_11_0),
		.io_in_b_0(b_25_0),
		.io_in_d_0(b_89_0),
		.io_in_control_0_dataflow(mesh_1_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_3_io_in_control_0_shift_b),
		.io_in_id_0(r_153_0),
		.io_in_last_0(r_217_0),
		.io_in_valid_0(r_89_0),
		.io_out_a_0(_mesh_1_3_io_out_a_0),
		.io_out_c_0(_mesh_1_3_io_out_c_0),
		.io_out_b_0(_mesh_1_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_3_io_out_id_0),
		.io_out_last_0(_mesh_1_3_io_out_last_0),
		.io_out_valid_0(_mesh_1_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((646 == GlobalFiModInstNr[0]) || (646 == GlobalFiModInstNr[1]) || (646 == GlobalFiModInstNr[2]) || (646 == GlobalFiModInstNr[3]))));
	Tile mesh_1_4(
		.clock(clock),
		.io_in_a_0(r_12_0),
		.io_in_b_0(b_33_0),
		.io_in_d_0(b_97_0),
		.io_in_control_0_dataflow(mesh_1_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_4_io_in_control_0_shift_b),
		.io_in_id_0(r_161_0),
		.io_in_last_0(r_225_0),
		.io_in_valid_0(r_97_0),
		.io_out_a_0(_mesh_1_4_io_out_a_0),
		.io_out_c_0(_mesh_1_4_io_out_c_0),
		.io_out_b_0(_mesh_1_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_4_io_out_id_0),
		.io_out_last_0(_mesh_1_4_io_out_last_0),
		.io_out_valid_0(_mesh_1_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((647 == GlobalFiModInstNr[0]) || (647 == GlobalFiModInstNr[1]) || (647 == GlobalFiModInstNr[2]) || (647 == GlobalFiModInstNr[3]))));
	Tile mesh_1_5(
		.clock(clock),
		.io_in_a_0(r_13_0),
		.io_in_b_0(b_41_0),
		.io_in_d_0(b_105_0),
		.io_in_control_0_dataflow(mesh_1_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_5_io_in_control_0_shift_b),
		.io_in_id_0(r_169_0),
		.io_in_last_0(r_233_0),
		.io_in_valid_0(r_105_0),
		.io_out_a_0(_mesh_1_5_io_out_a_0),
		.io_out_c_0(_mesh_1_5_io_out_c_0),
		.io_out_b_0(_mesh_1_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_5_io_out_id_0),
		.io_out_last_0(_mesh_1_5_io_out_last_0),
		.io_out_valid_0(_mesh_1_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((648 == GlobalFiModInstNr[0]) || (648 == GlobalFiModInstNr[1]) || (648 == GlobalFiModInstNr[2]) || (648 == GlobalFiModInstNr[3]))));
	Tile mesh_1_6(
		.clock(clock),
		.io_in_a_0(r_14_0),
		.io_in_b_0(b_49_0),
		.io_in_d_0(b_113_0),
		.io_in_control_0_dataflow(mesh_1_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_6_io_in_control_0_shift_b),
		.io_in_id_0(r_177_0),
		.io_in_last_0(r_241_0),
		.io_in_valid_0(r_113_0),
		.io_out_a_0(_mesh_1_6_io_out_a_0),
		.io_out_c_0(_mesh_1_6_io_out_c_0),
		.io_out_b_0(_mesh_1_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_6_io_out_id_0),
		.io_out_last_0(_mesh_1_6_io_out_last_0),
		.io_out_valid_0(_mesh_1_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((649 == GlobalFiModInstNr[0]) || (649 == GlobalFiModInstNr[1]) || (649 == GlobalFiModInstNr[2]) || (649 == GlobalFiModInstNr[3]))));
	Tile mesh_1_7(
		.clock(clock),
		.io_in_a_0(r_15_0),
		.io_in_b_0(b_57_0),
		.io_in_d_0(b_121_0),
		.io_in_control_0_dataflow(mesh_1_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_1_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_1_7_io_in_control_0_shift_b),
		.io_in_id_0(r_185_0),
		.io_in_last_0(r_249_0),
		.io_in_valid_0(r_121_0),
		.io_out_a_0(_mesh_1_7_io_out_a_0),
		.io_out_c_0(_mesh_1_7_io_out_c_0),
		.io_out_b_0(_mesh_1_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_1_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_1_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_1_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_1_7_io_out_id_0),
		.io_out_last_0(_mesh_1_7_io_out_last_0),
		.io_out_valid_0(_mesh_1_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((650 == GlobalFiModInstNr[0]) || (650 == GlobalFiModInstNr[1]) || (650 == GlobalFiModInstNr[2]) || (650 == GlobalFiModInstNr[3]))));
	Tile mesh_2_0(
		.clock(clock),
		.io_in_a_0(r_16_0),
		.io_in_b_0(b_2_0),
		.io_in_d_0(b_66_0),
		.io_in_control_0_dataflow(mesh_2_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_0_io_in_control_0_shift_b),
		.io_in_id_0(r_130_0),
		.io_in_last_0(r_194_0),
		.io_in_valid_0(r_66_0),
		.io_out_a_0(_mesh_2_0_io_out_a_0),
		.io_out_c_0(_mesh_2_0_io_out_c_0),
		.io_out_b_0(_mesh_2_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_0_io_out_id_0),
		.io_out_last_0(_mesh_2_0_io_out_last_0),
		.io_out_valid_0(_mesh_2_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((651 == GlobalFiModInstNr[0]) || (651 == GlobalFiModInstNr[1]) || (651 == GlobalFiModInstNr[2]) || (651 == GlobalFiModInstNr[3]))));
	Tile mesh_2_1(
		.clock(clock),
		.io_in_a_0(r_17_0),
		.io_in_b_0(b_10_0),
		.io_in_d_0(b_74_0),
		.io_in_control_0_dataflow(mesh_2_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_1_io_in_control_0_shift_b),
		.io_in_id_0(r_138_0),
		.io_in_last_0(r_202_0),
		.io_in_valid_0(r_74_0),
		.io_out_a_0(_mesh_2_1_io_out_a_0),
		.io_out_c_0(_mesh_2_1_io_out_c_0),
		.io_out_b_0(_mesh_2_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_1_io_out_id_0),
		.io_out_last_0(_mesh_2_1_io_out_last_0),
		.io_out_valid_0(_mesh_2_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((652 == GlobalFiModInstNr[0]) || (652 == GlobalFiModInstNr[1]) || (652 == GlobalFiModInstNr[2]) || (652 == GlobalFiModInstNr[3]))));
	Tile mesh_2_2(
		.clock(clock),
		.io_in_a_0(r_18_0),
		.io_in_b_0(b_18_0),
		.io_in_d_0(b_82_0),
		.io_in_control_0_dataflow(mesh_2_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_2_io_in_control_0_shift_b),
		.io_in_id_0(r_146_0),
		.io_in_last_0(r_210_0),
		.io_in_valid_0(r_82_0),
		.io_out_a_0(_mesh_2_2_io_out_a_0),
		.io_out_c_0(_mesh_2_2_io_out_c_0),
		.io_out_b_0(_mesh_2_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_2_io_out_id_0),
		.io_out_last_0(_mesh_2_2_io_out_last_0),
		.io_out_valid_0(_mesh_2_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((653 == GlobalFiModInstNr[0]) || (653 == GlobalFiModInstNr[1]) || (653 == GlobalFiModInstNr[2]) || (653 == GlobalFiModInstNr[3]))));
	Tile mesh_2_3(
		.clock(clock),
		.io_in_a_0(r_19_0),
		.io_in_b_0(b_26_0),
		.io_in_d_0(b_90_0),
		.io_in_control_0_dataflow(mesh_2_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_3_io_in_control_0_shift_b),
		.io_in_id_0(r_154_0),
		.io_in_last_0(r_218_0),
		.io_in_valid_0(r_90_0),
		.io_out_a_0(_mesh_2_3_io_out_a_0),
		.io_out_c_0(_mesh_2_3_io_out_c_0),
		.io_out_b_0(_mesh_2_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_3_io_out_id_0),
		.io_out_last_0(_mesh_2_3_io_out_last_0),
		.io_out_valid_0(_mesh_2_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((654 == GlobalFiModInstNr[0]) || (654 == GlobalFiModInstNr[1]) || (654 == GlobalFiModInstNr[2]) || (654 == GlobalFiModInstNr[3]))));
	Tile mesh_2_4(
		.clock(clock),
		.io_in_a_0(r_20_0),
		.io_in_b_0(b_34_0),
		.io_in_d_0(b_98_0),
		.io_in_control_0_dataflow(mesh_2_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_4_io_in_control_0_shift_b),
		.io_in_id_0(r_162_0),
		.io_in_last_0(r_226_0),
		.io_in_valid_0(r_98_0),
		.io_out_a_0(_mesh_2_4_io_out_a_0),
		.io_out_c_0(_mesh_2_4_io_out_c_0),
		.io_out_b_0(_mesh_2_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_4_io_out_id_0),
		.io_out_last_0(_mesh_2_4_io_out_last_0),
		.io_out_valid_0(_mesh_2_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((655 == GlobalFiModInstNr[0]) || (655 == GlobalFiModInstNr[1]) || (655 == GlobalFiModInstNr[2]) || (655 == GlobalFiModInstNr[3]))));
	Tile mesh_2_5(
		.clock(clock),
		.io_in_a_0(r_21_0),
		.io_in_b_0(b_42_0),
		.io_in_d_0(b_106_0),
		.io_in_control_0_dataflow(mesh_2_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_5_io_in_control_0_shift_b),
		.io_in_id_0(r_170_0),
		.io_in_last_0(r_234_0),
		.io_in_valid_0(r_106_0),
		.io_out_a_0(_mesh_2_5_io_out_a_0),
		.io_out_c_0(_mesh_2_5_io_out_c_0),
		.io_out_b_0(_mesh_2_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_5_io_out_id_0),
		.io_out_last_0(_mesh_2_5_io_out_last_0),
		.io_out_valid_0(_mesh_2_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((656 == GlobalFiModInstNr[0]) || (656 == GlobalFiModInstNr[1]) || (656 == GlobalFiModInstNr[2]) || (656 == GlobalFiModInstNr[3]))));
	Tile mesh_2_6(
		.clock(clock),
		.io_in_a_0(r_22_0),
		.io_in_b_0(b_50_0),
		.io_in_d_0(b_114_0),
		.io_in_control_0_dataflow(mesh_2_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_6_io_in_control_0_shift_b),
		.io_in_id_0(r_178_0),
		.io_in_last_0(r_242_0),
		.io_in_valid_0(r_114_0),
		.io_out_a_0(_mesh_2_6_io_out_a_0),
		.io_out_c_0(_mesh_2_6_io_out_c_0),
		.io_out_b_0(_mesh_2_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_6_io_out_id_0),
		.io_out_last_0(_mesh_2_6_io_out_last_0),
		.io_out_valid_0(_mesh_2_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((657 == GlobalFiModInstNr[0]) || (657 == GlobalFiModInstNr[1]) || (657 == GlobalFiModInstNr[2]) || (657 == GlobalFiModInstNr[3]))));
	Tile mesh_2_7(
		.clock(clock),
		.io_in_a_0(r_23_0),
		.io_in_b_0(b_58_0),
		.io_in_d_0(b_122_0),
		.io_in_control_0_dataflow(mesh_2_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_2_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_2_7_io_in_control_0_shift_b),
		.io_in_id_0(r_186_0),
		.io_in_last_0(r_250_0),
		.io_in_valid_0(r_122_0),
		.io_out_a_0(_mesh_2_7_io_out_a_0),
		.io_out_c_0(_mesh_2_7_io_out_c_0),
		.io_out_b_0(_mesh_2_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_2_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_2_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_2_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_2_7_io_out_id_0),
		.io_out_last_0(_mesh_2_7_io_out_last_0),
		.io_out_valid_0(_mesh_2_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((658 == GlobalFiModInstNr[0]) || (658 == GlobalFiModInstNr[1]) || (658 == GlobalFiModInstNr[2]) || (658 == GlobalFiModInstNr[3]))));
	Tile mesh_3_0(
		.clock(clock),
		.io_in_a_0(r_24_0),
		.io_in_b_0(b_3_0),
		.io_in_d_0(b_67_0),
		.io_in_control_0_dataflow(mesh_3_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_0_io_in_control_0_shift_b),
		.io_in_id_0(r_131_0),
		.io_in_last_0(r_195_0),
		.io_in_valid_0(r_67_0),
		.io_out_a_0(_mesh_3_0_io_out_a_0),
		.io_out_c_0(_mesh_3_0_io_out_c_0),
		.io_out_b_0(_mesh_3_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_0_io_out_id_0),
		.io_out_last_0(_mesh_3_0_io_out_last_0),
		.io_out_valid_0(_mesh_3_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((659 == GlobalFiModInstNr[0]) || (659 == GlobalFiModInstNr[1]) || (659 == GlobalFiModInstNr[2]) || (659 == GlobalFiModInstNr[3]))));
	Tile mesh_3_1(
		.clock(clock),
		.io_in_a_0(r_25_0),
		.io_in_b_0(b_11_0),
		.io_in_d_0(b_75_0),
		.io_in_control_0_dataflow(mesh_3_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_1_io_in_control_0_shift_b),
		.io_in_id_0(r_139_0),
		.io_in_last_0(r_203_0),
		.io_in_valid_0(r_75_0),
		.io_out_a_0(_mesh_3_1_io_out_a_0),
		.io_out_c_0(_mesh_3_1_io_out_c_0),
		.io_out_b_0(_mesh_3_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_1_io_out_id_0),
		.io_out_last_0(_mesh_3_1_io_out_last_0),
		.io_out_valid_0(_mesh_3_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((660 == GlobalFiModInstNr[0]) || (660 == GlobalFiModInstNr[1]) || (660 == GlobalFiModInstNr[2]) || (660 == GlobalFiModInstNr[3]))));
	Tile mesh_3_2(
		.clock(clock),
		.io_in_a_0(r_26_0),
		.io_in_b_0(b_19_0),
		.io_in_d_0(b_83_0),
		.io_in_control_0_dataflow(mesh_3_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_2_io_in_control_0_shift_b),
		.io_in_id_0(r_147_0),
		.io_in_last_0(r_211_0),
		.io_in_valid_0(r_83_0),
		.io_out_a_0(_mesh_3_2_io_out_a_0),
		.io_out_c_0(_mesh_3_2_io_out_c_0),
		.io_out_b_0(_mesh_3_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_2_io_out_id_0),
		.io_out_last_0(_mesh_3_2_io_out_last_0),
		.io_out_valid_0(_mesh_3_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((661 == GlobalFiModInstNr[0]) || (661 == GlobalFiModInstNr[1]) || (661 == GlobalFiModInstNr[2]) || (661 == GlobalFiModInstNr[3]))));
	Tile mesh_3_3(
		.clock(clock),
		.io_in_a_0(r_27_0),
		.io_in_b_0(b_27_0),
		.io_in_d_0(b_91_0),
		.io_in_control_0_dataflow(mesh_3_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_3_io_in_control_0_shift_b),
		.io_in_id_0(r_155_0),
		.io_in_last_0(r_219_0),
		.io_in_valid_0(r_91_0),
		.io_out_a_0(_mesh_3_3_io_out_a_0),
		.io_out_c_0(_mesh_3_3_io_out_c_0),
		.io_out_b_0(_mesh_3_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_3_io_out_id_0),
		.io_out_last_0(_mesh_3_3_io_out_last_0),
		.io_out_valid_0(_mesh_3_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((662 == GlobalFiModInstNr[0]) || (662 == GlobalFiModInstNr[1]) || (662 == GlobalFiModInstNr[2]) || (662 == GlobalFiModInstNr[3]))));
	Tile mesh_3_4(
		.clock(clock),
		.io_in_a_0(r_28_0),
		.io_in_b_0(b_35_0),
		.io_in_d_0(b_99_0),
		.io_in_control_0_dataflow(mesh_3_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_4_io_in_control_0_shift_b),
		.io_in_id_0(r_163_0),
		.io_in_last_0(r_227_0),
		.io_in_valid_0(r_99_0),
		.io_out_a_0(_mesh_3_4_io_out_a_0),
		.io_out_c_0(_mesh_3_4_io_out_c_0),
		.io_out_b_0(_mesh_3_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_4_io_out_id_0),
		.io_out_last_0(_mesh_3_4_io_out_last_0),
		.io_out_valid_0(_mesh_3_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((663 == GlobalFiModInstNr[0]) || (663 == GlobalFiModInstNr[1]) || (663 == GlobalFiModInstNr[2]) || (663 == GlobalFiModInstNr[3]))));
	Tile mesh_3_5(
		.clock(clock),
		.io_in_a_0(r_29_0),
		.io_in_b_0(b_43_0),
		.io_in_d_0(b_107_0),
		.io_in_control_0_dataflow(mesh_3_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_5_io_in_control_0_shift_b),
		.io_in_id_0(r_171_0),
		.io_in_last_0(r_235_0),
		.io_in_valid_0(r_107_0),
		.io_out_a_0(_mesh_3_5_io_out_a_0),
		.io_out_c_0(_mesh_3_5_io_out_c_0),
		.io_out_b_0(_mesh_3_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_5_io_out_id_0),
		.io_out_last_0(_mesh_3_5_io_out_last_0),
		.io_out_valid_0(_mesh_3_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((664 == GlobalFiModInstNr[0]) || (664 == GlobalFiModInstNr[1]) || (664 == GlobalFiModInstNr[2]) || (664 == GlobalFiModInstNr[3]))));
	Tile mesh_3_6(
		.clock(clock),
		.io_in_a_0(r_30_0),
		.io_in_b_0(b_51_0),
		.io_in_d_0(b_115_0),
		.io_in_control_0_dataflow(mesh_3_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_6_io_in_control_0_shift_b),
		.io_in_id_0(r_179_0),
		.io_in_last_0(r_243_0),
		.io_in_valid_0(r_115_0),
		.io_out_a_0(_mesh_3_6_io_out_a_0),
		.io_out_c_0(_mesh_3_6_io_out_c_0),
		.io_out_b_0(_mesh_3_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_6_io_out_id_0),
		.io_out_last_0(_mesh_3_6_io_out_last_0),
		.io_out_valid_0(_mesh_3_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((665 == GlobalFiModInstNr[0]) || (665 == GlobalFiModInstNr[1]) || (665 == GlobalFiModInstNr[2]) || (665 == GlobalFiModInstNr[3]))));
	Tile mesh_3_7(
		.clock(clock),
		.io_in_a_0(r_31_0),
		.io_in_b_0(b_59_0),
		.io_in_d_0(b_123_0),
		.io_in_control_0_dataflow(mesh_3_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_3_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_3_7_io_in_control_0_shift_b),
		.io_in_id_0(r_187_0),
		.io_in_last_0(r_251_0),
		.io_in_valid_0(r_123_0),
		.io_out_a_0(_mesh_3_7_io_out_a_0),
		.io_out_c_0(_mesh_3_7_io_out_c_0),
		.io_out_b_0(_mesh_3_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_3_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_3_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_3_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_3_7_io_out_id_0),
		.io_out_last_0(_mesh_3_7_io_out_last_0),
		.io_out_valid_0(_mesh_3_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((666 == GlobalFiModInstNr[0]) || (666 == GlobalFiModInstNr[1]) || (666 == GlobalFiModInstNr[2]) || (666 == GlobalFiModInstNr[3]))));
	Tile mesh_4_0(
		.clock(clock),
		.io_in_a_0(r_32_0),
		.io_in_b_0(b_4_0),
		.io_in_d_0(b_68_0),
		.io_in_control_0_dataflow(mesh_4_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_0_io_in_control_0_shift_b),
		.io_in_id_0(r_132_0),
		.io_in_last_0(r_196_0),
		.io_in_valid_0(r_68_0),
		.io_out_a_0(_mesh_4_0_io_out_a_0),
		.io_out_c_0(_mesh_4_0_io_out_c_0),
		.io_out_b_0(_mesh_4_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_0_io_out_id_0),
		.io_out_last_0(_mesh_4_0_io_out_last_0),
		.io_out_valid_0(_mesh_4_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((667 == GlobalFiModInstNr[0]) || (667 == GlobalFiModInstNr[1]) || (667 == GlobalFiModInstNr[2]) || (667 == GlobalFiModInstNr[3]))));
	Tile mesh_4_1(
		.clock(clock),
		.io_in_a_0(r_33_0),
		.io_in_b_0(b_12_0),
		.io_in_d_0(b_76_0),
		.io_in_control_0_dataflow(mesh_4_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_1_io_in_control_0_shift_b),
		.io_in_id_0(r_140_0),
		.io_in_last_0(r_204_0),
		.io_in_valid_0(r_76_0),
		.io_out_a_0(_mesh_4_1_io_out_a_0),
		.io_out_c_0(_mesh_4_1_io_out_c_0),
		.io_out_b_0(_mesh_4_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_1_io_out_id_0),
		.io_out_last_0(_mesh_4_1_io_out_last_0),
		.io_out_valid_0(_mesh_4_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((668 == GlobalFiModInstNr[0]) || (668 == GlobalFiModInstNr[1]) || (668 == GlobalFiModInstNr[2]) || (668 == GlobalFiModInstNr[3]))));
	Tile mesh_4_2(
		.clock(clock),
		.io_in_a_0(r_34_0),
		.io_in_b_0(b_20_0),
		.io_in_d_0(b_84_0),
		.io_in_control_0_dataflow(mesh_4_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_2_io_in_control_0_shift_b),
		.io_in_id_0(r_148_0),
		.io_in_last_0(r_212_0),
		.io_in_valid_0(r_84_0),
		.io_out_a_0(_mesh_4_2_io_out_a_0),
		.io_out_c_0(_mesh_4_2_io_out_c_0),
		.io_out_b_0(_mesh_4_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_2_io_out_id_0),
		.io_out_last_0(_mesh_4_2_io_out_last_0),
		.io_out_valid_0(_mesh_4_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((669 == GlobalFiModInstNr[0]) || (669 == GlobalFiModInstNr[1]) || (669 == GlobalFiModInstNr[2]) || (669 == GlobalFiModInstNr[3]))));
	Tile mesh_4_3(
		.clock(clock),
		.io_in_a_0(r_35_0),
		.io_in_b_0(b_28_0),
		.io_in_d_0(b_92_0),
		.io_in_control_0_dataflow(mesh_4_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_3_io_in_control_0_shift_b),
		.io_in_id_0(r_156_0),
		.io_in_last_0(r_220_0),
		.io_in_valid_0(r_92_0),
		.io_out_a_0(_mesh_4_3_io_out_a_0),
		.io_out_c_0(_mesh_4_3_io_out_c_0),
		.io_out_b_0(_mesh_4_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_3_io_out_id_0),
		.io_out_last_0(_mesh_4_3_io_out_last_0),
		.io_out_valid_0(_mesh_4_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((670 == GlobalFiModInstNr[0]) || (670 == GlobalFiModInstNr[1]) || (670 == GlobalFiModInstNr[2]) || (670 == GlobalFiModInstNr[3]))));
	Tile mesh_4_4(
		.clock(clock),
		.io_in_a_0(r_36_0),
		.io_in_b_0(b_36_0),
		.io_in_d_0(b_100_0),
		.io_in_control_0_dataflow(mesh_4_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_4_io_in_control_0_shift_b),
		.io_in_id_0(r_164_0),
		.io_in_last_0(r_228_0),
		.io_in_valid_0(r_100_0),
		.io_out_a_0(_mesh_4_4_io_out_a_0),
		.io_out_c_0(_mesh_4_4_io_out_c_0),
		.io_out_b_0(_mesh_4_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_4_io_out_id_0),
		.io_out_last_0(_mesh_4_4_io_out_last_0),
		.io_out_valid_0(_mesh_4_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((671 == GlobalFiModInstNr[0]) || (671 == GlobalFiModInstNr[1]) || (671 == GlobalFiModInstNr[2]) || (671 == GlobalFiModInstNr[3]))));
	Tile mesh_4_5(
		.clock(clock),
		.io_in_a_0(r_37_0),
		.io_in_b_0(b_44_0),
		.io_in_d_0(b_108_0),
		.io_in_control_0_dataflow(mesh_4_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_5_io_in_control_0_shift_b),
		.io_in_id_0(r_172_0),
		.io_in_last_0(r_236_0),
		.io_in_valid_0(r_108_0),
		.io_out_a_0(_mesh_4_5_io_out_a_0),
		.io_out_c_0(_mesh_4_5_io_out_c_0),
		.io_out_b_0(_mesh_4_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_5_io_out_id_0),
		.io_out_last_0(_mesh_4_5_io_out_last_0),
		.io_out_valid_0(_mesh_4_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((672 == GlobalFiModInstNr[0]) || (672 == GlobalFiModInstNr[1]) || (672 == GlobalFiModInstNr[2]) || (672 == GlobalFiModInstNr[3]))));
	Tile mesh_4_6(
		.clock(clock),
		.io_in_a_0(r_38_0),
		.io_in_b_0(b_52_0),
		.io_in_d_0(b_116_0),
		.io_in_control_0_dataflow(mesh_4_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_6_io_in_control_0_shift_b),
		.io_in_id_0(r_180_0),
		.io_in_last_0(r_244_0),
		.io_in_valid_0(r_116_0),
		.io_out_a_0(_mesh_4_6_io_out_a_0),
		.io_out_c_0(_mesh_4_6_io_out_c_0),
		.io_out_b_0(_mesh_4_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_6_io_out_id_0),
		.io_out_last_0(_mesh_4_6_io_out_last_0),
		.io_out_valid_0(_mesh_4_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((673 == GlobalFiModInstNr[0]) || (673 == GlobalFiModInstNr[1]) || (673 == GlobalFiModInstNr[2]) || (673 == GlobalFiModInstNr[3]))));
	Tile mesh_4_7(
		.clock(clock),
		.io_in_a_0(r_39_0),
		.io_in_b_0(b_60_0),
		.io_in_d_0(b_124_0),
		.io_in_control_0_dataflow(mesh_4_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_4_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_4_7_io_in_control_0_shift_b),
		.io_in_id_0(r_188_0),
		.io_in_last_0(r_252_0),
		.io_in_valid_0(r_124_0),
		.io_out_a_0(_mesh_4_7_io_out_a_0),
		.io_out_c_0(_mesh_4_7_io_out_c_0),
		.io_out_b_0(_mesh_4_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_4_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_4_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_4_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_4_7_io_out_id_0),
		.io_out_last_0(_mesh_4_7_io_out_last_0),
		.io_out_valid_0(_mesh_4_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((674 == GlobalFiModInstNr[0]) || (674 == GlobalFiModInstNr[1]) || (674 == GlobalFiModInstNr[2]) || (674 == GlobalFiModInstNr[3]))));
	Tile mesh_5_0(
		.clock(clock),
		.io_in_a_0(r_40_0),
		.io_in_b_0(b_5_0),
		.io_in_d_0(b_69_0),
		.io_in_control_0_dataflow(mesh_5_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_0_io_in_control_0_shift_b),
		.io_in_id_0(r_133_0),
		.io_in_last_0(r_197_0),
		.io_in_valid_0(r_69_0),
		.io_out_a_0(_mesh_5_0_io_out_a_0),
		.io_out_c_0(_mesh_5_0_io_out_c_0),
		.io_out_b_0(_mesh_5_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_0_io_out_id_0),
		.io_out_last_0(_mesh_5_0_io_out_last_0),
		.io_out_valid_0(_mesh_5_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((675 == GlobalFiModInstNr[0]) || (675 == GlobalFiModInstNr[1]) || (675 == GlobalFiModInstNr[2]) || (675 == GlobalFiModInstNr[3]))));
	Tile mesh_5_1(
		.clock(clock),
		.io_in_a_0(r_41_0),
		.io_in_b_0(b_13_0),
		.io_in_d_0(b_77_0),
		.io_in_control_0_dataflow(mesh_5_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_1_io_in_control_0_shift_b),
		.io_in_id_0(r_141_0),
		.io_in_last_0(r_205_0),
		.io_in_valid_0(r_77_0),
		.io_out_a_0(_mesh_5_1_io_out_a_0),
		.io_out_c_0(_mesh_5_1_io_out_c_0),
		.io_out_b_0(_mesh_5_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_1_io_out_id_0),
		.io_out_last_0(_mesh_5_1_io_out_last_0),
		.io_out_valid_0(_mesh_5_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((676 == GlobalFiModInstNr[0]) || (676 == GlobalFiModInstNr[1]) || (676 == GlobalFiModInstNr[2]) || (676 == GlobalFiModInstNr[3]))));
	Tile mesh_5_2(
		.clock(clock),
		.io_in_a_0(r_42_0),
		.io_in_b_0(b_21_0),
		.io_in_d_0(b_85_0),
		.io_in_control_0_dataflow(mesh_5_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_2_io_in_control_0_shift_b),
		.io_in_id_0(r_149_0),
		.io_in_last_0(r_213_0),
		.io_in_valid_0(r_85_0),
		.io_out_a_0(_mesh_5_2_io_out_a_0),
		.io_out_c_0(_mesh_5_2_io_out_c_0),
		.io_out_b_0(_mesh_5_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_2_io_out_id_0),
		.io_out_last_0(_mesh_5_2_io_out_last_0),
		.io_out_valid_0(_mesh_5_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((677 == GlobalFiModInstNr[0]) || (677 == GlobalFiModInstNr[1]) || (677 == GlobalFiModInstNr[2]) || (677 == GlobalFiModInstNr[3]))));
	Tile mesh_5_3(
		.clock(clock),
		.io_in_a_0(r_43_0),
		.io_in_b_0(b_29_0),
		.io_in_d_0(b_93_0),
		.io_in_control_0_dataflow(mesh_5_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_3_io_in_control_0_shift_b),
		.io_in_id_0(r_157_0),
		.io_in_last_0(r_221_0),
		.io_in_valid_0(r_93_0),
		.io_out_a_0(_mesh_5_3_io_out_a_0),
		.io_out_c_0(_mesh_5_3_io_out_c_0),
		.io_out_b_0(_mesh_5_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_3_io_out_id_0),
		.io_out_last_0(_mesh_5_3_io_out_last_0),
		.io_out_valid_0(_mesh_5_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((678 == GlobalFiModInstNr[0]) || (678 == GlobalFiModInstNr[1]) || (678 == GlobalFiModInstNr[2]) || (678 == GlobalFiModInstNr[3]))));
	Tile mesh_5_4(
		.clock(clock),
		.io_in_a_0(r_44_0),
		.io_in_b_0(b_37_0),
		.io_in_d_0(b_101_0),
		.io_in_control_0_dataflow(mesh_5_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_4_io_in_control_0_shift_b),
		.io_in_id_0(r_165_0),
		.io_in_last_0(r_229_0),
		.io_in_valid_0(r_101_0),
		.io_out_a_0(_mesh_5_4_io_out_a_0),
		.io_out_c_0(_mesh_5_4_io_out_c_0),
		.io_out_b_0(_mesh_5_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_4_io_out_id_0),
		.io_out_last_0(_mesh_5_4_io_out_last_0),
		.io_out_valid_0(_mesh_5_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((679 == GlobalFiModInstNr[0]) || (679 == GlobalFiModInstNr[1]) || (679 == GlobalFiModInstNr[2]) || (679 == GlobalFiModInstNr[3]))));
	Tile mesh_5_5(
		.clock(clock),
		.io_in_a_0(r_45_0),
		.io_in_b_0(b_45_0),
		.io_in_d_0(b_109_0),
		.io_in_control_0_dataflow(mesh_5_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_5_io_in_control_0_shift_b),
		.io_in_id_0(r_173_0),
		.io_in_last_0(r_237_0),
		.io_in_valid_0(r_109_0),
		.io_out_a_0(_mesh_5_5_io_out_a_0),
		.io_out_c_0(_mesh_5_5_io_out_c_0),
		.io_out_b_0(_mesh_5_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_5_io_out_id_0),
		.io_out_last_0(_mesh_5_5_io_out_last_0),
		.io_out_valid_0(_mesh_5_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((680 == GlobalFiModInstNr[0]) || (680 == GlobalFiModInstNr[1]) || (680 == GlobalFiModInstNr[2]) || (680 == GlobalFiModInstNr[3]))));
	Tile mesh_5_6(
		.clock(clock),
		.io_in_a_0(r_46_0),
		.io_in_b_0(b_53_0),
		.io_in_d_0(b_117_0),
		.io_in_control_0_dataflow(mesh_5_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_6_io_in_control_0_shift_b),
		.io_in_id_0(r_181_0),
		.io_in_last_0(r_245_0),
		.io_in_valid_0(r_117_0),
		.io_out_a_0(_mesh_5_6_io_out_a_0),
		.io_out_c_0(_mesh_5_6_io_out_c_0),
		.io_out_b_0(_mesh_5_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_6_io_out_id_0),
		.io_out_last_0(_mesh_5_6_io_out_last_0),
		.io_out_valid_0(_mesh_5_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((681 == GlobalFiModInstNr[0]) || (681 == GlobalFiModInstNr[1]) || (681 == GlobalFiModInstNr[2]) || (681 == GlobalFiModInstNr[3]))));
	Tile mesh_5_7(
		.clock(clock),
		.io_in_a_0(r_47_0),
		.io_in_b_0(b_61_0),
		.io_in_d_0(b_125_0),
		.io_in_control_0_dataflow(mesh_5_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_5_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_5_7_io_in_control_0_shift_b),
		.io_in_id_0(r_189_0),
		.io_in_last_0(r_253_0),
		.io_in_valid_0(r_125_0),
		.io_out_a_0(_mesh_5_7_io_out_a_0),
		.io_out_c_0(_mesh_5_7_io_out_c_0),
		.io_out_b_0(_mesh_5_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_5_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_5_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_5_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_5_7_io_out_id_0),
		.io_out_last_0(_mesh_5_7_io_out_last_0),
		.io_out_valid_0(_mesh_5_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((682 == GlobalFiModInstNr[0]) || (682 == GlobalFiModInstNr[1]) || (682 == GlobalFiModInstNr[2]) || (682 == GlobalFiModInstNr[3]))));
	Tile mesh_6_0(
		.clock(clock),
		.io_in_a_0(r_48_0),
		.io_in_b_0(b_6_0),
		.io_in_d_0(b_70_0),
		.io_in_control_0_dataflow(mesh_6_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_0_io_in_control_0_shift_b),
		.io_in_id_0(r_134_0),
		.io_in_last_0(r_198_0),
		.io_in_valid_0(r_70_0),
		.io_out_a_0(_mesh_6_0_io_out_a_0),
		.io_out_c_0(_mesh_6_0_io_out_c_0),
		.io_out_b_0(_mesh_6_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_0_io_out_id_0),
		.io_out_last_0(_mesh_6_0_io_out_last_0),
		.io_out_valid_0(_mesh_6_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((683 == GlobalFiModInstNr[0]) || (683 == GlobalFiModInstNr[1]) || (683 == GlobalFiModInstNr[2]) || (683 == GlobalFiModInstNr[3]))));
	Tile mesh_6_1(
		.clock(clock),
		.io_in_a_0(r_49_0),
		.io_in_b_0(b_14_0),
		.io_in_d_0(b_78_0),
		.io_in_control_0_dataflow(mesh_6_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_1_io_in_control_0_shift_b),
		.io_in_id_0(r_142_0),
		.io_in_last_0(r_206_0),
		.io_in_valid_0(r_78_0),
		.io_out_a_0(_mesh_6_1_io_out_a_0),
		.io_out_c_0(_mesh_6_1_io_out_c_0),
		.io_out_b_0(_mesh_6_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_1_io_out_id_0),
		.io_out_last_0(_mesh_6_1_io_out_last_0),
		.io_out_valid_0(_mesh_6_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((684 == GlobalFiModInstNr[0]) || (684 == GlobalFiModInstNr[1]) || (684 == GlobalFiModInstNr[2]) || (684 == GlobalFiModInstNr[3]))));
	Tile mesh_6_2(
		.clock(clock),
		.io_in_a_0(r_50_0),
		.io_in_b_0(b_22_0),
		.io_in_d_0(b_86_0),
		.io_in_control_0_dataflow(mesh_6_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_2_io_in_control_0_shift_b),
		.io_in_id_0(r_150_0),
		.io_in_last_0(r_214_0),
		.io_in_valid_0(r_86_0),
		.io_out_a_0(_mesh_6_2_io_out_a_0),
		.io_out_c_0(_mesh_6_2_io_out_c_0),
		.io_out_b_0(_mesh_6_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_2_io_out_id_0),
		.io_out_last_0(_mesh_6_2_io_out_last_0),
		.io_out_valid_0(_mesh_6_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((685 == GlobalFiModInstNr[0]) || (685 == GlobalFiModInstNr[1]) || (685 == GlobalFiModInstNr[2]) || (685 == GlobalFiModInstNr[3]))));
	Tile mesh_6_3(
		.clock(clock),
		.io_in_a_0(r_51_0),
		.io_in_b_0(b_30_0),
		.io_in_d_0(b_94_0),
		.io_in_control_0_dataflow(mesh_6_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_3_io_in_control_0_shift_b),
		.io_in_id_0(r_158_0),
		.io_in_last_0(r_222_0),
		.io_in_valid_0(r_94_0),
		.io_out_a_0(_mesh_6_3_io_out_a_0),
		.io_out_c_0(_mesh_6_3_io_out_c_0),
		.io_out_b_0(_mesh_6_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_3_io_out_id_0),
		.io_out_last_0(_mesh_6_3_io_out_last_0),
		.io_out_valid_0(_mesh_6_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((686 == GlobalFiModInstNr[0]) || (686 == GlobalFiModInstNr[1]) || (686 == GlobalFiModInstNr[2]) || (686 == GlobalFiModInstNr[3]))));
	Tile mesh_6_4(
		.clock(clock),
		.io_in_a_0(r_52_0),
		.io_in_b_0(b_38_0),
		.io_in_d_0(b_102_0),
		.io_in_control_0_dataflow(mesh_6_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_4_io_in_control_0_shift_b),
		.io_in_id_0(r_166_0),
		.io_in_last_0(r_230_0),
		.io_in_valid_0(r_102_0),
		.io_out_a_0(_mesh_6_4_io_out_a_0),
		.io_out_c_0(_mesh_6_4_io_out_c_0),
		.io_out_b_0(_mesh_6_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_4_io_out_id_0),
		.io_out_last_0(_mesh_6_4_io_out_last_0),
		.io_out_valid_0(_mesh_6_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((687 == GlobalFiModInstNr[0]) || (687 == GlobalFiModInstNr[1]) || (687 == GlobalFiModInstNr[2]) || (687 == GlobalFiModInstNr[3]))));
	Tile mesh_6_5(
		.clock(clock),
		.io_in_a_0(r_53_0),
		.io_in_b_0(b_46_0),
		.io_in_d_0(b_110_0),
		.io_in_control_0_dataflow(mesh_6_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_5_io_in_control_0_shift_b),
		.io_in_id_0(r_174_0),
		.io_in_last_0(r_238_0),
		.io_in_valid_0(r_110_0),
		.io_out_a_0(_mesh_6_5_io_out_a_0),
		.io_out_c_0(_mesh_6_5_io_out_c_0),
		.io_out_b_0(_mesh_6_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_5_io_out_id_0),
		.io_out_last_0(_mesh_6_5_io_out_last_0),
		.io_out_valid_0(_mesh_6_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((688 == GlobalFiModInstNr[0]) || (688 == GlobalFiModInstNr[1]) || (688 == GlobalFiModInstNr[2]) || (688 == GlobalFiModInstNr[3]))));
	Tile mesh_6_6(
		.clock(clock),
		.io_in_a_0(r_54_0),
		.io_in_b_0(b_54_0),
		.io_in_d_0(b_118_0),
		.io_in_control_0_dataflow(mesh_6_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_6_io_in_control_0_shift_b),
		.io_in_id_0(r_182_0),
		.io_in_last_0(r_246_0),
		.io_in_valid_0(r_118_0),
		.io_out_a_0(_mesh_6_6_io_out_a_0),
		.io_out_c_0(_mesh_6_6_io_out_c_0),
		.io_out_b_0(_mesh_6_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_6_io_out_id_0),
		.io_out_last_0(_mesh_6_6_io_out_last_0),
		.io_out_valid_0(_mesh_6_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((689 == GlobalFiModInstNr[0]) || (689 == GlobalFiModInstNr[1]) || (689 == GlobalFiModInstNr[2]) || (689 == GlobalFiModInstNr[3]))));
	Tile mesh_6_7(
		.clock(clock),
		.io_in_a_0(r_55_0),
		.io_in_b_0(b_62_0),
		.io_in_d_0(b_126_0),
		.io_in_control_0_dataflow(mesh_6_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_6_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_6_7_io_in_control_0_shift_b),
		.io_in_id_0(r_190_0),
		.io_in_last_0(r_254_0),
		.io_in_valid_0(r_126_0),
		.io_out_a_0(_mesh_6_7_io_out_a_0),
		.io_out_c_0(_mesh_6_7_io_out_c_0),
		.io_out_b_0(_mesh_6_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_6_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_6_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_6_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_6_7_io_out_id_0),
		.io_out_last_0(_mesh_6_7_io_out_last_0),
		.io_out_valid_0(_mesh_6_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((690 == GlobalFiModInstNr[0]) || (690 == GlobalFiModInstNr[1]) || (690 == GlobalFiModInstNr[2]) || (690 == GlobalFiModInstNr[3]))));
	Tile mesh_7_0(
		.clock(clock),
		.io_in_a_0(r_56_0),
		.io_in_b_0(b_7_0),
		.io_in_d_0(b_71_0),
		.io_in_control_0_dataflow(mesh_7_0_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_0_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_0_io_in_control_0_shift_b),
		.io_in_id_0(r_135_0),
		.io_in_last_0(r_199_0),
		.io_in_valid_0(r_71_0),
		.io_out_a_0(_mesh_7_0_io_out_a_0),
		.io_out_c_0(_mesh_7_0_io_out_c_0),
		.io_out_b_0(_mesh_7_0_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_0_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_0_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_0_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_0_io_out_id_0),
		.io_out_last_0(_mesh_7_0_io_out_last_0),
		.io_out_valid_0(_mesh_7_0_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((691 == GlobalFiModInstNr[0]) || (691 == GlobalFiModInstNr[1]) || (691 == GlobalFiModInstNr[2]) || (691 == GlobalFiModInstNr[3]))));
	Tile mesh_7_1(
		.clock(clock),
		.io_in_a_0(r_57_0),
		.io_in_b_0(b_15_0),
		.io_in_d_0(b_79_0),
		.io_in_control_0_dataflow(mesh_7_1_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_1_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_1_io_in_control_0_shift_b),
		.io_in_id_0(r_143_0),
		.io_in_last_0(r_207_0),
		.io_in_valid_0(r_79_0),
		.io_out_a_0(_mesh_7_1_io_out_a_0),
		.io_out_c_0(_mesh_7_1_io_out_c_0),
		.io_out_b_0(_mesh_7_1_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_1_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_1_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_1_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_1_io_out_id_0),
		.io_out_last_0(_mesh_7_1_io_out_last_0),
		.io_out_valid_0(_mesh_7_1_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((692 == GlobalFiModInstNr[0]) || (692 == GlobalFiModInstNr[1]) || (692 == GlobalFiModInstNr[2]) || (692 == GlobalFiModInstNr[3]))));
	Tile mesh_7_2(
		.clock(clock),
		.io_in_a_0(r_58_0),
		.io_in_b_0(b_23_0),
		.io_in_d_0(b_87_0),
		.io_in_control_0_dataflow(mesh_7_2_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_2_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_2_io_in_control_0_shift_b),
		.io_in_id_0(r_151_0),
		.io_in_last_0(r_215_0),
		.io_in_valid_0(r_87_0),
		.io_out_a_0(_mesh_7_2_io_out_a_0),
		.io_out_c_0(_mesh_7_2_io_out_c_0),
		.io_out_b_0(_mesh_7_2_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_2_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_2_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_2_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_2_io_out_id_0),
		.io_out_last_0(_mesh_7_2_io_out_last_0),
		.io_out_valid_0(_mesh_7_2_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((693 == GlobalFiModInstNr[0]) || (693 == GlobalFiModInstNr[1]) || (693 == GlobalFiModInstNr[2]) || (693 == GlobalFiModInstNr[3]))));
	Tile mesh_7_3(
		.clock(clock),
		.io_in_a_0(r_59_0),
		.io_in_b_0(b_31_0),
		.io_in_d_0(b_95_0),
		.io_in_control_0_dataflow(mesh_7_3_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_3_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_3_io_in_control_0_shift_b),
		.io_in_id_0(r_159_0),
		.io_in_last_0(r_223_0),
		.io_in_valid_0(r_95_0),
		.io_out_a_0(_mesh_7_3_io_out_a_0),
		.io_out_c_0(_mesh_7_3_io_out_c_0),
		.io_out_b_0(_mesh_7_3_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_3_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_3_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_3_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_3_io_out_id_0),
		.io_out_last_0(_mesh_7_3_io_out_last_0),
		.io_out_valid_0(_mesh_7_3_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((694 == GlobalFiModInstNr[0]) || (694 == GlobalFiModInstNr[1]) || (694 == GlobalFiModInstNr[2]) || (694 == GlobalFiModInstNr[3]))));
	Tile mesh_7_4(
		.clock(clock),
		.io_in_a_0(r_60_0),
		.io_in_b_0(b_39_0),
		.io_in_d_0(b_103_0),
		.io_in_control_0_dataflow(mesh_7_4_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_4_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_4_io_in_control_0_shift_b),
		.io_in_id_0(r_167_0),
		.io_in_last_0(r_231_0),
		.io_in_valid_0(r_103_0),
		.io_out_a_0(_mesh_7_4_io_out_a_0),
		.io_out_c_0(_mesh_7_4_io_out_c_0),
		.io_out_b_0(_mesh_7_4_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_4_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_4_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_4_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_4_io_out_id_0),
		.io_out_last_0(_mesh_7_4_io_out_last_0),
		.io_out_valid_0(_mesh_7_4_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((695 == GlobalFiModInstNr[0]) || (695 == GlobalFiModInstNr[1]) || (695 == GlobalFiModInstNr[2]) || (695 == GlobalFiModInstNr[3]))));
	Tile mesh_7_5(
		.clock(clock),
		.io_in_a_0(r_61_0),
		.io_in_b_0(b_47_0),
		.io_in_d_0(b_111_0),
		.io_in_control_0_dataflow(mesh_7_5_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_5_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_5_io_in_control_0_shift_b),
		.io_in_id_0(r_175_0),
		.io_in_last_0(r_239_0),
		.io_in_valid_0(r_111_0),
		.io_out_a_0(_mesh_7_5_io_out_a_0),
		.io_out_c_0(_mesh_7_5_io_out_c_0),
		.io_out_b_0(_mesh_7_5_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_5_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_5_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_5_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_5_io_out_id_0),
		.io_out_last_0(_mesh_7_5_io_out_last_0),
		.io_out_valid_0(_mesh_7_5_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((696 == GlobalFiModInstNr[0]) || (696 == GlobalFiModInstNr[1]) || (696 == GlobalFiModInstNr[2]) || (696 == GlobalFiModInstNr[3]))));
	Tile mesh_7_6(
		.clock(clock),
		.io_in_a_0(r_62_0),
		.io_in_b_0(b_55_0),
		.io_in_d_0(b_119_0),
		.io_in_control_0_dataflow(mesh_7_6_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_6_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_6_io_in_control_0_shift_b),
		.io_in_id_0(r_183_0),
		.io_in_last_0(r_247_0),
		.io_in_valid_0(r_119_0),
		.io_out_a_0(_mesh_7_6_io_out_a_0),
		.io_out_c_0(_mesh_7_6_io_out_c_0),
		.io_out_b_0(_mesh_7_6_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_6_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_6_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_6_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_6_io_out_id_0),
		.io_out_last_0(_mesh_7_6_io_out_last_0),
		.io_out_valid_0(_mesh_7_6_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((697 == GlobalFiModInstNr[0]) || (697 == GlobalFiModInstNr[1]) || (697 == GlobalFiModInstNr[2]) || (697 == GlobalFiModInstNr[3]))));
	Tile mesh_7_7(
		.clock(clock),
		.io_in_a_0(r_63_0),
		.io_in_b_0(b_63_0),
		.io_in_d_0(b_127_0),
		.io_in_control_0_dataflow(mesh_7_7_io_in_control_0_dataflow_b),
		.io_in_control_0_propagate(mesh_7_7_io_in_control_0_propagate_b),
		.io_in_control_0_shift(mesh_7_7_io_in_control_0_shift_b),
		.io_in_id_0(r_191_0),
		.io_in_last_0(r_255_0),
		.io_in_valid_0(r_127_0),
		.io_out_a_0(_mesh_7_7_io_out_a_0),
		.io_out_c_0(_mesh_7_7_io_out_c_0),
		.io_out_b_0(_mesh_7_7_io_out_b_0),
		.io_out_control_0_dataflow(_mesh_7_7_io_out_control_0_dataflow),
		.io_out_control_0_propagate(_mesh_7_7_io_out_control_0_propagate),
		.io_out_control_0_shift(_mesh_7_7_io_out_control_0_shift),
		.io_out_id_0(_mesh_7_7_io_out_id_0),
		.io_out_last_0(_mesh_7_7_io_out_last_0),
		.io_out_valid_0(_mesh_7_7_io_out_valid_0)
	,
    .fiEnable(fiEnable && ((698 == GlobalFiModInstNr[0]) || (698 == GlobalFiModInstNr[1]) || (698 == GlobalFiModInstNr[2]) || (698 == GlobalFiModInstNr[3]))));
	assign io_out_b_0_0 =( r_256_0) ^ ((fiEnable && (613 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_1_0 =( r_262_0) ^ ((fiEnable && (614 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_2_0 =( r_268_0) ^ ((fiEnable && (615 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_3_0 =( r_274_0) ^ ((fiEnable && (616 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_4_0 =( r_280_0) ^ ((fiEnable && (617 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_5_0 =( r_286_0) ^ ((fiEnable && (618 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_6_0 =( r_292_0) ^ ((fiEnable && (619 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_b_7_0 =( r_298_0) ^ ((fiEnable && (620 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_0_0 =( r_257_0) ^ ((fiEnable && (621 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_1_0 =( r_263_0) ^ ((fiEnable && (622 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_2_0 =( r_269_0) ^ ((fiEnable && (623 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_3_0 =( r_275_0) ^ ((fiEnable && (624 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_4_0 =( r_281_0) ^ ((fiEnable && (625 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_5_0 =( r_287_0) ^ ((fiEnable && (626 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_6_0 =( r_293_0) ^ ((fiEnable && (627 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_c_7_0 =( r_299_0) ^ ((fiEnable && (628 == GlobalFiNumber)) ? GlobalFiSignal[31:0] : {32{1'b0}});
	assign io_out_valid_0_0 =( r_258_0) ^ ((fiEnable && (629 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_control_0_0_dataflow =( r_259_0_dataflow) ^ ((fiEnable && (630 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
	assign io_out_id_0_0 =( r_260_0) ^ ((fiEnable && (631 == GlobalFiNumber)) ? GlobalFiSignal[2:0] : {3{1'b0}});
	assign io_out_last_0_0 =( r_261_0) ^ ((fiEnable && (632 == GlobalFiNumber)) ? GlobalFiSignal[0] : {1{1'b0}});
endmodule